magic
tech sky130A
magscale 1 2
timestamp 1668282613
<< pwell >>
rect 945 14715 4089 17471
<< psubdiff >>
rect 971 17421 4063 17445
rect 971 17406 1168 17421
rect 971 17372 995 17406
rect 1029 17372 1067 17406
rect 1101 17387 1168 17406
rect 1202 17387 1240 17421
rect 1274 17387 1312 17421
rect 1346 17387 1384 17421
rect 1418 17387 1456 17421
rect 1490 17387 1528 17421
rect 1562 17387 1600 17421
rect 1634 17387 1672 17421
rect 1706 17387 1744 17421
rect 1778 17387 1816 17421
rect 1850 17387 1888 17421
rect 1922 17387 1960 17421
rect 1994 17387 2032 17421
rect 2066 17387 2104 17421
rect 2138 17387 2176 17421
rect 2210 17387 2248 17421
rect 2282 17387 2320 17421
rect 2354 17387 2392 17421
rect 2426 17387 2464 17421
rect 2498 17387 2536 17421
rect 2570 17387 2608 17421
rect 2642 17387 2680 17421
rect 2714 17387 2752 17421
rect 2786 17387 2824 17421
rect 2858 17387 2896 17421
rect 2930 17387 2968 17421
rect 3002 17387 3040 17421
rect 3074 17387 3112 17421
rect 3146 17387 3184 17421
rect 3218 17387 3256 17421
rect 3290 17387 3328 17421
rect 3362 17387 3400 17421
rect 3434 17387 3472 17421
rect 3506 17387 3544 17421
rect 3578 17387 3616 17421
rect 3650 17387 3688 17421
rect 3722 17387 3760 17421
rect 3794 17387 3832 17421
rect 3866 17406 4063 17421
rect 3866 17387 3933 17406
rect 1101 17372 3933 17387
rect 3967 17372 4005 17406
rect 4039 17372 4063 17406
rect 971 17349 4063 17372
rect 971 17334 1168 17349
rect 971 17300 995 17334
rect 1029 17300 1067 17334
rect 1101 17315 1168 17334
rect 1202 17315 1240 17349
rect 1274 17315 1312 17349
rect 1346 17315 1384 17349
rect 1418 17315 1456 17349
rect 1490 17315 1528 17349
rect 1562 17315 1600 17349
rect 1634 17315 1672 17349
rect 1706 17315 1744 17349
rect 1778 17315 1816 17349
rect 1850 17315 1888 17349
rect 1922 17315 1960 17349
rect 1994 17315 2032 17349
rect 2066 17315 2104 17349
rect 2138 17315 2176 17349
rect 2210 17315 2248 17349
rect 2282 17315 2320 17349
rect 2354 17315 2392 17349
rect 2426 17315 2464 17349
rect 2498 17315 2536 17349
rect 2570 17315 2608 17349
rect 2642 17315 2680 17349
rect 2714 17315 2752 17349
rect 2786 17315 2824 17349
rect 2858 17315 2896 17349
rect 2930 17315 2968 17349
rect 3002 17315 3040 17349
rect 3074 17315 3112 17349
rect 3146 17315 3184 17349
rect 3218 17315 3256 17349
rect 3290 17315 3328 17349
rect 3362 17315 3400 17349
rect 3434 17315 3472 17349
rect 3506 17315 3544 17349
rect 3578 17315 3616 17349
rect 3650 17315 3688 17349
rect 3722 17315 3760 17349
rect 3794 17315 3832 17349
rect 3866 17334 4063 17349
rect 3866 17315 3933 17334
rect 1101 17300 3933 17315
rect 3967 17300 4005 17334
rect 4039 17300 4063 17334
rect 971 17291 4063 17300
rect 971 17262 1125 17291
rect 971 17228 995 17262
rect 1029 17228 1067 17262
rect 1101 17228 1125 17262
rect 971 17190 1125 17228
rect 971 17156 995 17190
rect 1029 17156 1067 17190
rect 1101 17156 1125 17190
rect 971 17118 1125 17156
rect 971 17084 995 17118
rect 1029 17084 1067 17118
rect 1101 17084 1125 17118
rect 971 17046 1125 17084
rect 971 17012 995 17046
rect 1029 17012 1067 17046
rect 1101 17012 1125 17046
rect 971 16974 1125 17012
rect 971 16940 995 16974
rect 1029 16940 1067 16974
rect 1101 16940 1125 16974
rect 971 16902 1125 16940
rect 971 16868 995 16902
rect 1029 16868 1067 16902
rect 1101 16868 1125 16902
rect 971 16830 1125 16868
rect 971 16796 995 16830
rect 1029 16796 1067 16830
rect 1101 16796 1125 16830
rect 971 16758 1125 16796
rect 971 16724 995 16758
rect 1029 16724 1067 16758
rect 1101 16724 1125 16758
rect 971 16686 1125 16724
rect 971 16652 995 16686
rect 1029 16652 1067 16686
rect 1101 16652 1125 16686
rect 971 16614 1125 16652
rect 971 16580 995 16614
rect 1029 16580 1067 16614
rect 1101 16580 1125 16614
rect 971 16542 1125 16580
rect 971 16508 995 16542
rect 1029 16508 1067 16542
rect 1101 16508 1125 16542
rect 971 16470 1125 16508
rect 971 16436 995 16470
rect 1029 16436 1067 16470
rect 1101 16436 1125 16470
rect 971 16398 1125 16436
rect 971 16364 995 16398
rect 1029 16364 1067 16398
rect 1101 16364 1125 16398
rect 971 16326 1125 16364
rect 971 16292 995 16326
rect 1029 16292 1067 16326
rect 1101 16292 1125 16326
rect 971 16254 1125 16292
rect 971 16220 995 16254
rect 1029 16220 1067 16254
rect 1101 16220 1125 16254
rect 971 16182 1125 16220
rect 971 16148 995 16182
rect 1029 16148 1067 16182
rect 1101 16148 1125 16182
rect 971 16110 1125 16148
rect 971 16076 995 16110
rect 1029 16076 1067 16110
rect 1101 16076 1125 16110
rect 971 16038 1125 16076
rect 971 16004 995 16038
rect 1029 16004 1067 16038
rect 1101 16004 1125 16038
rect 971 15966 1125 16004
rect 971 15932 995 15966
rect 1029 15932 1067 15966
rect 1101 15932 1125 15966
rect 971 15894 1125 15932
rect 971 15860 995 15894
rect 1029 15860 1067 15894
rect 1101 15860 1125 15894
rect 971 15822 1125 15860
rect 971 15788 995 15822
rect 1029 15788 1067 15822
rect 1101 15788 1125 15822
rect 971 15750 1125 15788
rect 971 15716 995 15750
rect 1029 15716 1067 15750
rect 1101 15716 1125 15750
rect 971 15678 1125 15716
rect 971 15644 995 15678
rect 1029 15644 1067 15678
rect 1101 15644 1125 15678
rect 971 15606 1125 15644
rect 971 15572 995 15606
rect 1029 15572 1067 15606
rect 1101 15572 1125 15606
rect 971 15534 1125 15572
rect 971 15500 995 15534
rect 1029 15500 1067 15534
rect 1101 15500 1125 15534
rect 971 15462 1125 15500
rect 971 15428 995 15462
rect 1029 15428 1067 15462
rect 1101 15428 1125 15462
rect 971 15390 1125 15428
rect 971 15356 995 15390
rect 1029 15356 1067 15390
rect 1101 15356 1125 15390
rect 971 15318 1125 15356
rect 971 15284 995 15318
rect 1029 15284 1067 15318
rect 1101 15284 1125 15318
rect 971 15246 1125 15284
rect 971 15212 995 15246
rect 1029 15212 1067 15246
rect 1101 15212 1125 15246
rect 971 15174 1125 15212
rect 971 15140 995 15174
rect 1029 15140 1067 15174
rect 1101 15140 1125 15174
rect 971 15102 1125 15140
rect 971 15068 995 15102
rect 1029 15068 1067 15102
rect 1101 15068 1125 15102
rect 971 15030 1125 15068
rect 971 14996 995 15030
rect 1029 14996 1067 15030
rect 1101 14996 1125 15030
rect 971 14958 1125 14996
rect 971 14924 995 14958
rect 1029 14924 1067 14958
rect 1101 14924 1125 14958
rect 971 14895 1125 14924
rect 3909 17262 4063 17291
rect 3909 17228 3933 17262
rect 3967 17228 4005 17262
rect 4039 17228 4063 17262
rect 3909 17190 4063 17228
rect 3909 17156 3933 17190
rect 3967 17156 4005 17190
rect 4039 17156 4063 17190
rect 3909 17118 4063 17156
rect 3909 17084 3933 17118
rect 3967 17084 4005 17118
rect 4039 17084 4063 17118
rect 3909 17046 4063 17084
rect 3909 17012 3933 17046
rect 3967 17012 4005 17046
rect 4039 17012 4063 17046
rect 3909 16974 4063 17012
rect 3909 16940 3933 16974
rect 3967 16940 4005 16974
rect 4039 16940 4063 16974
rect 3909 16902 4063 16940
rect 3909 16868 3933 16902
rect 3967 16868 4005 16902
rect 4039 16868 4063 16902
rect 3909 16830 4063 16868
rect 3909 16796 3933 16830
rect 3967 16796 4005 16830
rect 4039 16796 4063 16830
rect 3909 16758 4063 16796
rect 3909 16724 3933 16758
rect 3967 16724 4005 16758
rect 4039 16724 4063 16758
rect 3909 16686 4063 16724
rect 3909 16652 3933 16686
rect 3967 16652 4005 16686
rect 4039 16652 4063 16686
rect 3909 16614 4063 16652
rect 3909 16580 3933 16614
rect 3967 16580 4005 16614
rect 4039 16580 4063 16614
rect 3909 16542 4063 16580
rect 3909 16508 3933 16542
rect 3967 16508 4005 16542
rect 4039 16508 4063 16542
rect 3909 16470 4063 16508
rect 3909 16436 3933 16470
rect 3967 16436 4005 16470
rect 4039 16436 4063 16470
rect 3909 16398 4063 16436
rect 3909 16364 3933 16398
rect 3967 16364 4005 16398
rect 4039 16364 4063 16398
rect 3909 16326 4063 16364
rect 3909 16292 3933 16326
rect 3967 16292 4005 16326
rect 4039 16292 4063 16326
rect 3909 16254 4063 16292
rect 3909 16220 3933 16254
rect 3967 16220 4005 16254
rect 4039 16220 4063 16254
rect 3909 16182 4063 16220
rect 3909 16148 3933 16182
rect 3967 16148 4005 16182
rect 4039 16148 4063 16182
rect 3909 16110 4063 16148
rect 3909 16076 3933 16110
rect 3967 16076 4005 16110
rect 4039 16076 4063 16110
rect 3909 16038 4063 16076
rect 3909 16004 3933 16038
rect 3967 16004 4005 16038
rect 4039 16004 4063 16038
rect 3909 15966 4063 16004
rect 3909 15932 3933 15966
rect 3967 15932 4005 15966
rect 4039 15932 4063 15966
rect 3909 15894 4063 15932
rect 3909 15860 3933 15894
rect 3967 15860 4005 15894
rect 4039 15860 4063 15894
rect 3909 15822 4063 15860
rect 3909 15788 3933 15822
rect 3967 15788 4005 15822
rect 4039 15788 4063 15822
rect 3909 15750 4063 15788
rect 3909 15716 3933 15750
rect 3967 15716 4005 15750
rect 4039 15716 4063 15750
rect 3909 15678 4063 15716
rect 3909 15644 3933 15678
rect 3967 15644 4005 15678
rect 4039 15644 4063 15678
rect 3909 15606 4063 15644
rect 3909 15572 3933 15606
rect 3967 15572 4005 15606
rect 4039 15572 4063 15606
rect 3909 15534 4063 15572
rect 3909 15500 3933 15534
rect 3967 15500 4005 15534
rect 4039 15500 4063 15534
rect 3909 15462 4063 15500
rect 3909 15428 3933 15462
rect 3967 15428 4005 15462
rect 4039 15428 4063 15462
rect 3909 15390 4063 15428
rect 3909 15356 3933 15390
rect 3967 15356 4005 15390
rect 4039 15356 4063 15390
rect 3909 15318 4063 15356
rect 3909 15284 3933 15318
rect 3967 15284 4005 15318
rect 4039 15284 4063 15318
rect 3909 15246 4063 15284
rect 3909 15212 3933 15246
rect 3967 15212 4005 15246
rect 4039 15212 4063 15246
rect 3909 15174 4063 15212
rect 3909 15140 3933 15174
rect 3967 15140 4005 15174
rect 4039 15140 4063 15174
rect 3909 15102 4063 15140
rect 3909 15068 3933 15102
rect 3967 15068 4005 15102
rect 4039 15068 4063 15102
rect 3909 15030 4063 15068
rect 3909 14996 3933 15030
rect 3967 14996 4005 15030
rect 4039 14996 4063 15030
rect 3909 14958 4063 14996
rect 3909 14924 3933 14958
rect 3967 14924 4005 14958
rect 4039 14924 4063 14958
rect 3909 14895 4063 14924
rect 971 14886 4063 14895
rect 971 14852 995 14886
rect 1029 14852 1067 14886
rect 1101 14871 3933 14886
rect 1101 14852 1168 14871
rect 971 14837 1168 14852
rect 1202 14837 1240 14871
rect 1274 14837 1312 14871
rect 1346 14837 1384 14871
rect 1418 14837 1456 14871
rect 1490 14837 1528 14871
rect 1562 14837 1600 14871
rect 1634 14837 1672 14871
rect 1706 14837 1744 14871
rect 1778 14837 1816 14871
rect 1850 14837 1888 14871
rect 1922 14837 1960 14871
rect 1994 14837 2032 14871
rect 2066 14837 2104 14871
rect 2138 14837 2176 14871
rect 2210 14837 2248 14871
rect 2282 14837 2320 14871
rect 2354 14837 2392 14871
rect 2426 14837 2464 14871
rect 2498 14837 2536 14871
rect 2570 14837 2608 14871
rect 2642 14837 2680 14871
rect 2714 14837 2752 14871
rect 2786 14837 2824 14871
rect 2858 14837 2896 14871
rect 2930 14837 2968 14871
rect 3002 14837 3040 14871
rect 3074 14837 3112 14871
rect 3146 14837 3184 14871
rect 3218 14837 3256 14871
rect 3290 14837 3328 14871
rect 3362 14837 3400 14871
rect 3434 14837 3472 14871
rect 3506 14837 3544 14871
rect 3578 14837 3616 14871
rect 3650 14837 3688 14871
rect 3722 14837 3760 14871
rect 3794 14837 3832 14871
rect 3866 14852 3933 14871
rect 3967 14852 4005 14886
rect 4039 14852 4063 14886
rect 3866 14837 4063 14852
rect 971 14814 4063 14837
rect 971 14780 995 14814
rect 1029 14780 1067 14814
rect 1101 14799 3933 14814
rect 1101 14780 1168 14799
rect 971 14765 1168 14780
rect 1202 14765 1240 14799
rect 1274 14765 1312 14799
rect 1346 14765 1384 14799
rect 1418 14765 1456 14799
rect 1490 14765 1528 14799
rect 1562 14765 1600 14799
rect 1634 14765 1672 14799
rect 1706 14765 1744 14799
rect 1778 14765 1816 14799
rect 1850 14765 1888 14799
rect 1922 14765 1960 14799
rect 1994 14765 2032 14799
rect 2066 14765 2104 14799
rect 2138 14765 2176 14799
rect 2210 14765 2248 14799
rect 2282 14765 2320 14799
rect 2354 14765 2392 14799
rect 2426 14765 2464 14799
rect 2498 14765 2536 14799
rect 2570 14765 2608 14799
rect 2642 14765 2680 14799
rect 2714 14765 2752 14799
rect 2786 14765 2824 14799
rect 2858 14765 2896 14799
rect 2930 14765 2968 14799
rect 3002 14765 3040 14799
rect 3074 14765 3112 14799
rect 3146 14765 3184 14799
rect 3218 14765 3256 14799
rect 3290 14765 3328 14799
rect 3362 14765 3400 14799
rect 3434 14765 3472 14799
rect 3506 14765 3544 14799
rect 3578 14765 3616 14799
rect 3650 14765 3688 14799
rect 3722 14765 3760 14799
rect 3794 14765 3832 14799
rect 3866 14780 3933 14799
rect 3967 14780 4005 14814
rect 4039 14780 4063 14814
rect 3866 14765 4063 14780
rect 971 14741 4063 14765
<< psubdiffcont >>
rect 995 17372 1029 17406
rect 1067 17372 1101 17406
rect 1168 17387 1202 17421
rect 1240 17387 1274 17421
rect 1312 17387 1346 17421
rect 1384 17387 1418 17421
rect 1456 17387 1490 17421
rect 1528 17387 1562 17421
rect 1600 17387 1634 17421
rect 1672 17387 1706 17421
rect 1744 17387 1778 17421
rect 1816 17387 1850 17421
rect 1888 17387 1922 17421
rect 1960 17387 1994 17421
rect 2032 17387 2066 17421
rect 2104 17387 2138 17421
rect 2176 17387 2210 17421
rect 2248 17387 2282 17421
rect 2320 17387 2354 17421
rect 2392 17387 2426 17421
rect 2464 17387 2498 17421
rect 2536 17387 2570 17421
rect 2608 17387 2642 17421
rect 2680 17387 2714 17421
rect 2752 17387 2786 17421
rect 2824 17387 2858 17421
rect 2896 17387 2930 17421
rect 2968 17387 3002 17421
rect 3040 17387 3074 17421
rect 3112 17387 3146 17421
rect 3184 17387 3218 17421
rect 3256 17387 3290 17421
rect 3328 17387 3362 17421
rect 3400 17387 3434 17421
rect 3472 17387 3506 17421
rect 3544 17387 3578 17421
rect 3616 17387 3650 17421
rect 3688 17387 3722 17421
rect 3760 17387 3794 17421
rect 3832 17387 3866 17421
rect 3933 17372 3967 17406
rect 4005 17372 4039 17406
rect 995 17300 1029 17334
rect 1067 17300 1101 17334
rect 1168 17315 1202 17349
rect 1240 17315 1274 17349
rect 1312 17315 1346 17349
rect 1384 17315 1418 17349
rect 1456 17315 1490 17349
rect 1528 17315 1562 17349
rect 1600 17315 1634 17349
rect 1672 17315 1706 17349
rect 1744 17315 1778 17349
rect 1816 17315 1850 17349
rect 1888 17315 1922 17349
rect 1960 17315 1994 17349
rect 2032 17315 2066 17349
rect 2104 17315 2138 17349
rect 2176 17315 2210 17349
rect 2248 17315 2282 17349
rect 2320 17315 2354 17349
rect 2392 17315 2426 17349
rect 2464 17315 2498 17349
rect 2536 17315 2570 17349
rect 2608 17315 2642 17349
rect 2680 17315 2714 17349
rect 2752 17315 2786 17349
rect 2824 17315 2858 17349
rect 2896 17315 2930 17349
rect 2968 17315 3002 17349
rect 3040 17315 3074 17349
rect 3112 17315 3146 17349
rect 3184 17315 3218 17349
rect 3256 17315 3290 17349
rect 3328 17315 3362 17349
rect 3400 17315 3434 17349
rect 3472 17315 3506 17349
rect 3544 17315 3578 17349
rect 3616 17315 3650 17349
rect 3688 17315 3722 17349
rect 3760 17315 3794 17349
rect 3832 17315 3866 17349
rect 3933 17300 3967 17334
rect 4005 17300 4039 17334
rect 995 17228 1029 17262
rect 1067 17228 1101 17262
rect 995 17156 1029 17190
rect 1067 17156 1101 17190
rect 995 17084 1029 17118
rect 1067 17084 1101 17118
rect 995 17012 1029 17046
rect 1067 17012 1101 17046
rect 995 16940 1029 16974
rect 1067 16940 1101 16974
rect 995 16868 1029 16902
rect 1067 16868 1101 16902
rect 995 16796 1029 16830
rect 1067 16796 1101 16830
rect 995 16724 1029 16758
rect 1067 16724 1101 16758
rect 995 16652 1029 16686
rect 1067 16652 1101 16686
rect 995 16580 1029 16614
rect 1067 16580 1101 16614
rect 995 16508 1029 16542
rect 1067 16508 1101 16542
rect 995 16436 1029 16470
rect 1067 16436 1101 16470
rect 995 16364 1029 16398
rect 1067 16364 1101 16398
rect 995 16292 1029 16326
rect 1067 16292 1101 16326
rect 995 16220 1029 16254
rect 1067 16220 1101 16254
rect 995 16148 1029 16182
rect 1067 16148 1101 16182
rect 995 16076 1029 16110
rect 1067 16076 1101 16110
rect 995 16004 1029 16038
rect 1067 16004 1101 16038
rect 995 15932 1029 15966
rect 1067 15932 1101 15966
rect 995 15860 1029 15894
rect 1067 15860 1101 15894
rect 995 15788 1029 15822
rect 1067 15788 1101 15822
rect 995 15716 1029 15750
rect 1067 15716 1101 15750
rect 995 15644 1029 15678
rect 1067 15644 1101 15678
rect 995 15572 1029 15606
rect 1067 15572 1101 15606
rect 995 15500 1029 15534
rect 1067 15500 1101 15534
rect 995 15428 1029 15462
rect 1067 15428 1101 15462
rect 995 15356 1029 15390
rect 1067 15356 1101 15390
rect 995 15284 1029 15318
rect 1067 15284 1101 15318
rect 995 15212 1029 15246
rect 1067 15212 1101 15246
rect 995 15140 1029 15174
rect 1067 15140 1101 15174
rect 995 15068 1029 15102
rect 1067 15068 1101 15102
rect 995 14996 1029 15030
rect 1067 14996 1101 15030
rect 995 14924 1029 14958
rect 1067 14924 1101 14958
rect 3933 17228 3967 17262
rect 4005 17228 4039 17262
rect 3933 17156 3967 17190
rect 4005 17156 4039 17190
rect 3933 17084 3967 17118
rect 4005 17084 4039 17118
rect 3933 17012 3967 17046
rect 4005 17012 4039 17046
rect 3933 16940 3967 16974
rect 4005 16940 4039 16974
rect 3933 16868 3967 16902
rect 4005 16868 4039 16902
rect 3933 16796 3967 16830
rect 4005 16796 4039 16830
rect 3933 16724 3967 16758
rect 4005 16724 4039 16758
rect 3933 16652 3967 16686
rect 4005 16652 4039 16686
rect 3933 16580 3967 16614
rect 4005 16580 4039 16614
rect 3933 16508 3967 16542
rect 4005 16508 4039 16542
rect 3933 16436 3967 16470
rect 4005 16436 4039 16470
rect 3933 16364 3967 16398
rect 4005 16364 4039 16398
rect 3933 16292 3967 16326
rect 4005 16292 4039 16326
rect 3933 16220 3967 16254
rect 4005 16220 4039 16254
rect 3933 16148 3967 16182
rect 4005 16148 4039 16182
rect 3933 16076 3967 16110
rect 4005 16076 4039 16110
rect 3933 16004 3967 16038
rect 4005 16004 4039 16038
rect 3933 15932 3967 15966
rect 4005 15932 4039 15966
rect 3933 15860 3967 15894
rect 4005 15860 4039 15894
rect 3933 15788 3967 15822
rect 4005 15788 4039 15822
rect 3933 15716 3967 15750
rect 4005 15716 4039 15750
rect 3933 15644 3967 15678
rect 4005 15644 4039 15678
rect 3933 15572 3967 15606
rect 4005 15572 4039 15606
rect 3933 15500 3967 15534
rect 4005 15500 4039 15534
rect 3933 15428 3967 15462
rect 4005 15428 4039 15462
rect 3933 15356 3967 15390
rect 4005 15356 4039 15390
rect 3933 15284 3967 15318
rect 4005 15284 4039 15318
rect 3933 15212 3967 15246
rect 4005 15212 4039 15246
rect 3933 15140 3967 15174
rect 4005 15140 4039 15174
rect 3933 15068 3967 15102
rect 4005 15068 4039 15102
rect 3933 14996 3967 15030
rect 4005 14996 4039 15030
rect 3933 14924 3967 14958
rect 4005 14924 4039 14958
rect 995 14852 1029 14886
rect 1067 14852 1101 14886
rect 1168 14837 1202 14871
rect 1240 14837 1274 14871
rect 1312 14837 1346 14871
rect 1384 14837 1418 14871
rect 1456 14837 1490 14871
rect 1528 14837 1562 14871
rect 1600 14837 1634 14871
rect 1672 14837 1706 14871
rect 1744 14837 1778 14871
rect 1816 14837 1850 14871
rect 1888 14837 1922 14871
rect 1960 14837 1994 14871
rect 2032 14837 2066 14871
rect 2104 14837 2138 14871
rect 2176 14837 2210 14871
rect 2248 14837 2282 14871
rect 2320 14837 2354 14871
rect 2392 14837 2426 14871
rect 2464 14837 2498 14871
rect 2536 14837 2570 14871
rect 2608 14837 2642 14871
rect 2680 14837 2714 14871
rect 2752 14837 2786 14871
rect 2824 14837 2858 14871
rect 2896 14837 2930 14871
rect 2968 14837 3002 14871
rect 3040 14837 3074 14871
rect 3112 14837 3146 14871
rect 3184 14837 3218 14871
rect 3256 14837 3290 14871
rect 3328 14837 3362 14871
rect 3400 14837 3434 14871
rect 3472 14837 3506 14871
rect 3544 14837 3578 14871
rect 3616 14837 3650 14871
rect 3688 14837 3722 14871
rect 3760 14837 3794 14871
rect 3832 14837 3866 14871
rect 3933 14852 3967 14886
rect 4005 14852 4039 14886
rect 995 14780 1029 14814
rect 1067 14780 1101 14814
rect 1168 14765 1202 14799
rect 1240 14765 1274 14799
rect 1312 14765 1346 14799
rect 1384 14765 1418 14799
rect 1456 14765 1490 14799
rect 1528 14765 1562 14799
rect 1600 14765 1634 14799
rect 1672 14765 1706 14799
rect 1744 14765 1778 14799
rect 1816 14765 1850 14799
rect 1888 14765 1922 14799
rect 1960 14765 1994 14799
rect 2032 14765 2066 14799
rect 2104 14765 2138 14799
rect 2176 14765 2210 14799
rect 2248 14765 2282 14799
rect 2320 14765 2354 14799
rect 2392 14765 2426 14799
rect 2464 14765 2498 14799
rect 2536 14765 2570 14799
rect 2608 14765 2642 14799
rect 2680 14765 2714 14799
rect 2752 14765 2786 14799
rect 2824 14765 2858 14799
rect 2896 14765 2930 14799
rect 2968 14765 3002 14799
rect 3040 14765 3074 14799
rect 3112 14765 3146 14799
rect 3184 14765 3218 14799
rect 3256 14765 3290 14799
rect 3328 14765 3362 14799
rect 3400 14765 3434 14799
rect 3472 14765 3506 14799
rect 3544 14765 3578 14799
rect 3616 14765 3650 14799
rect 3688 14765 3722 14799
rect 3760 14765 3794 14799
rect 3832 14765 3866 14799
rect 3933 14780 3967 14814
rect 4005 14780 4039 14814
<< locali >>
rect 979 17421 4055 17437
rect 979 17406 1168 17421
rect 979 14780 995 17406
rect 1101 17315 1168 17406
rect 3866 17406 4055 17421
rect 3866 17315 3933 17406
rect 1101 17299 3933 17315
rect 1101 14887 1117 17299
rect 3917 14887 3933 17299
rect 1101 14871 3933 14887
rect 1101 14780 1168 14871
rect 979 14765 1168 14780
rect 3866 14780 3933 14871
rect 4039 14780 4055 17406
rect 3866 14765 4055 14780
rect 979 14749 4055 14765
<< viali >>
rect 995 17372 1029 17406
rect 1029 17372 1067 17406
rect 1067 17372 1101 17406
rect 995 17334 1101 17372
rect 995 17300 1029 17334
rect 1029 17300 1067 17334
rect 1067 17300 1101 17334
rect 1168 17387 1202 17421
rect 1202 17387 1240 17421
rect 1240 17387 1274 17421
rect 1274 17387 1312 17421
rect 1312 17387 1346 17421
rect 1346 17387 1384 17421
rect 1384 17387 1418 17421
rect 1418 17387 1456 17421
rect 1456 17387 1490 17421
rect 1490 17387 1528 17421
rect 1528 17387 1562 17421
rect 1562 17387 1600 17421
rect 1600 17387 1634 17421
rect 1634 17387 1672 17421
rect 1672 17387 1706 17421
rect 1706 17387 1744 17421
rect 1744 17387 1778 17421
rect 1778 17387 1816 17421
rect 1816 17387 1850 17421
rect 1850 17387 1888 17421
rect 1888 17387 1922 17421
rect 1922 17387 1960 17421
rect 1960 17387 1994 17421
rect 1994 17387 2032 17421
rect 2032 17387 2066 17421
rect 2066 17387 2104 17421
rect 2104 17387 2138 17421
rect 2138 17387 2176 17421
rect 2176 17387 2210 17421
rect 2210 17387 2248 17421
rect 2248 17387 2282 17421
rect 2282 17387 2320 17421
rect 2320 17387 2354 17421
rect 2354 17387 2392 17421
rect 2392 17387 2426 17421
rect 2426 17387 2464 17421
rect 2464 17387 2498 17421
rect 2498 17387 2536 17421
rect 2536 17387 2570 17421
rect 2570 17387 2608 17421
rect 2608 17387 2642 17421
rect 2642 17387 2680 17421
rect 2680 17387 2714 17421
rect 2714 17387 2752 17421
rect 2752 17387 2786 17421
rect 2786 17387 2824 17421
rect 2824 17387 2858 17421
rect 2858 17387 2896 17421
rect 2896 17387 2930 17421
rect 2930 17387 2968 17421
rect 2968 17387 3002 17421
rect 3002 17387 3040 17421
rect 3040 17387 3074 17421
rect 3074 17387 3112 17421
rect 3112 17387 3146 17421
rect 3146 17387 3184 17421
rect 3184 17387 3218 17421
rect 3218 17387 3256 17421
rect 3256 17387 3290 17421
rect 3290 17387 3328 17421
rect 3328 17387 3362 17421
rect 3362 17387 3400 17421
rect 3400 17387 3434 17421
rect 3434 17387 3472 17421
rect 3472 17387 3506 17421
rect 3506 17387 3544 17421
rect 3544 17387 3578 17421
rect 3578 17387 3616 17421
rect 3616 17387 3650 17421
rect 3650 17387 3688 17421
rect 3688 17387 3722 17421
rect 3722 17387 3760 17421
rect 3760 17387 3794 17421
rect 3794 17387 3832 17421
rect 3832 17387 3866 17421
rect 1168 17349 3866 17387
rect 1168 17315 1202 17349
rect 1202 17315 1240 17349
rect 1240 17315 1274 17349
rect 1274 17315 1312 17349
rect 1312 17315 1346 17349
rect 1346 17315 1384 17349
rect 1384 17315 1418 17349
rect 1418 17315 1456 17349
rect 1456 17315 1490 17349
rect 1490 17315 1528 17349
rect 1528 17315 1562 17349
rect 1562 17315 1600 17349
rect 1600 17315 1634 17349
rect 1634 17315 1672 17349
rect 1672 17315 1706 17349
rect 1706 17315 1744 17349
rect 1744 17315 1778 17349
rect 1778 17315 1816 17349
rect 1816 17315 1850 17349
rect 1850 17315 1888 17349
rect 1888 17315 1922 17349
rect 1922 17315 1960 17349
rect 1960 17315 1994 17349
rect 1994 17315 2032 17349
rect 2032 17315 2066 17349
rect 2066 17315 2104 17349
rect 2104 17315 2138 17349
rect 2138 17315 2176 17349
rect 2176 17315 2210 17349
rect 2210 17315 2248 17349
rect 2248 17315 2282 17349
rect 2282 17315 2320 17349
rect 2320 17315 2354 17349
rect 2354 17315 2392 17349
rect 2392 17315 2426 17349
rect 2426 17315 2464 17349
rect 2464 17315 2498 17349
rect 2498 17315 2536 17349
rect 2536 17315 2570 17349
rect 2570 17315 2608 17349
rect 2608 17315 2642 17349
rect 2642 17315 2680 17349
rect 2680 17315 2714 17349
rect 2714 17315 2752 17349
rect 2752 17315 2786 17349
rect 2786 17315 2824 17349
rect 2824 17315 2858 17349
rect 2858 17315 2896 17349
rect 2896 17315 2930 17349
rect 2930 17315 2968 17349
rect 2968 17315 3002 17349
rect 3002 17315 3040 17349
rect 3040 17315 3074 17349
rect 3074 17315 3112 17349
rect 3112 17315 3146 17349
rect 3146 17315 3184 17349
rect 3184 17315 3218 17349
rect 3218 17315 3256 17349
rect 3256 17315 3290 17349
rect 3290 17315 3328 17349
rect 3328 17315 3362 17349
rect 3362 17315 3400 17349
rect 3400 17315 3434 17349
rect 3434 17315 3472 17349
rect 3472 17315 3506 17349
rect 3506 17315 3544 17349
rect 3544 17315 3578 17349
rect 3578 17315 3616 17349
rect 3616 17315 3650 17349
rect 3650 17315 3688 17349
rect 3688 17315 3722 17349
rect 3722 17315 3760 17349
rect 3760 17315 3794 17349
rect 3794 17315 3832 17349
rect 3832 17315 3866 17349
rect 3933 17372 3967 17406
rect 3967 17372 4005 17406
rect 4005 17372 4039 17406
rect 3933 17334 4039 17372
rect 995 17262 1101 17300
rect 3933 17300 3967 17334
rect 3967 17300 4005 17334
rect 4005 17300 4039 17334
rect 995 17228 1029 17262
rect 1029 17228 1067 17262
rect 1067 17228 1101 17262
rect 995 17190 1101 17228
rect 995 17156 1029 17190
rect 1029 17156 1067 17190
rect 1067 17156 1101 17190
rect 995 17118 1101 17156
rect 995 17084 1029 17118
rect 1029 17084 1067 17118
rect 1067 17084 1101 17118
rect 995 17046 1101 17084
rect 995 17012 1029 17046
rect 1029 17012 1067 17046
rect 1067 17012 1101 17046
rect 995 16974 1101 17012
rect 995 16940 1029 16974
rect 1029 16940 1067 16974
rect 1067 16940 1101 16974
rect 995 16902 1101 16940
rect 995 16868 1029 16902
rect 1029 16868 1067 16902
rect 1067 16868 1101 16902
rect 995 16830 1101 16868
rect 995 16796 1029 16830
rect 1029 16796 1067 16830
rect 1067 16796 1101 16830
rect 995 16758 1101 16796
rect 995 16724 1029 16758
rect 1029 16724 1067 16758
rect 1067 16724 1101 16758
rect 995 16686 1101 16724
rect 995 16652 1029 16686
rect 1029 16652 1067 16686
rect 1067 16652 1101 16686
rect 995 16614 1101 16652
rect 995 16580 1029 16614
rect 1029 16580 1067 16614
rect 1067 16580 1101 16614
rect 995 16542 1101 16580
rect 995 16508 1029 16542
rect 1029 16508 1067 16542
rect 1067 16508 1101 16542
rect 995 16470 1101 16508
rect 995 16436 1029 16470
rect 1029 16436 1067 16470
rect 1067 16436 1101 16470
rect 995 16398 1101 16436
rect 995 16364 1029 16398
rect 1029 16364 1067 16398
rect 1067 16364 1101 16398
rect 995 16326 1101 16364
rect 995 16292 1029 16326
rect 1029 16292 1067 16326
rect 1067 16292 1101 16326
rect 995 16254 1101 16292
rect 995 16220 1029 16254
rect 1029 16220 1067 16254
rect 1067 16220 1101 16254
rect 995 16182 1101 16220
rect 995 16148 1029 16182
rect 1029 16148 1067 16182
rect 1067 16148 1101 16182
rect 995 16110 1101 16148
rect 995 16076 1029 16110
rect 1029 16076 1067 16110
rect 1067 16076 1101 16110
rect 995 16038 1101 16076
rect 995 16004 1029 16038
rect 1029 16004 1067 16038
rect 1067 16004 1101 16038
rect 995 15966 1101 16004
rect 995 15932 1029 15966
rect 1029 15932 1067 15966
rect 1067 15932 1101 15966
rect 995 15894 1101 15932
rect 995 15860 1029 15894
rect 1029 15860 1067 15894
rect 1067 15860 1101 15894
rect 995 15822 1101 15860
rect 995 15788 1029 15822
rect 1029 15788 1067 15822
rect 1067 15788 1101 15822
rect 995 15750 1101 15788
rect 995 15716 1029 15750
rect 1029 15716 1067 15750
rect 1067 15716 1101 15750
rect 995 15678 1101 15716
rect 995 15644 1029 15678
rect 1029 15644 1067 15678
rect 1067 15644 1101 15678
rect 995 15606 1101 15644
rect 995 15572 1029 15606
rect 1029 15572 1067 15606
rect 1067 15572 1101 15606
rect 995 15534 1101 15572
rect 995 15500 1029 15534
rect 1029 15500 1067 15534
rect 1067 15500 1101 15534
rect 995 15462 1101 15500
rect 995 15428 1029 15462
rect 1029 15428 1067 15462
rect 1067 15428 1101 15462
rect 995 15390 1101 15428
rect 995 15356 1029 15390
rect 1029 15356 1067 15390
rect 1067 15356 1101 15390
rect 995 15318 1101 15356
rect 995 15284 1029 15318
rect 1029 15284 1067 15318
rect 1067 15284 1101 15318
rect 995 15246 1101 15284
rect 995 15212 1029 15246
rect 1029 15212 1067 15246
rect 1067 15212 1101 15246
rect 995 15174 1101 15212
rect 995 15140 1029 15174
rect 1029 15140 1067 15174
rect 1067 15140 1101 15174
rect 995 15102 1101 15140
rect 995 15068 1029 15102
rect 1029 15068 1067 15102
rect 1067 15068 1101 15102
rect 995 15030 1101 15068
rect 995 14996 1029 15030
rect 1029 14996 1067 15030
rect 1067 14996 1101 15030
rect 995 14958 1101 14996
rect 995 14924 1029 14958
rect 1029 14924 1067 14958
rect 1067 14924 1101 14958
rect 995 14886 1101 14924
rect 3933 17262 4039 17300
rect 3933 17228 3967 17262
rect 3967 17228 4005 17262
rect 4005 17228 4039 17262
rect 3933 17190 4039 17228
rect 3933 17156 3967 17190
rect 3967 17156 4005 17190
rect 4005 17156 4039 17190
rect 3933 17118 4039 17156
rect 3933 17084 3967 17118
rect 3967 17084 4005 17118
rect 4005 17084 4039 17118
rect 3933 17046 4039 17084
rect 3933 17012 3967 17046
rect 3967 17012 4005 17046
rect 4005 17012 4039 17046
rect 3933 16974 4039 17012
rect 3933 16940 3967 16974
rect 3967 16940 4005 16974
rect 4005 16940 4039 16974
rect 3933 16902 4039 16940
rect 3933 16868 3967 16902
rect 3967 16868 4005 16902
rect 4005 16868 4039 16902
rect 3933 16830 4039 16868
rect 3933 16796 3967 16830
rect 3967 16796 4005 16830
rect 4005 16796 4039 16830
rect 3933 16758 4039 16796
rect 3933 16724 3967 16758
rect 3967 16724 4005 16758
rect 4005 16724 4039 16758
rect 3933 16686 4039 16724
rect 3933 16652 3967 16686
rect 3967 16652 4005 16686
rect 4005 16652 4039 16686
rect 3933 16614 4039 16652
rect 3933 16580 3967 16614
rect 3967 16580 4005 16614
rect 4005 16580 4039 16614
rect 3933 16542 4039 16580
rect 3933 16508 3967 16542
rect 3967 16508 4005 16542
rect 4005 16508 4039 16542
rect 3933 16470 4039 16508
rect 3933 16436 3967 16470
rect 3967 16436 4005 16470
rect 4005 16436 4039 16470
rect 3933 16398 4039 16436
rect 3933 16364 3967 16398
rect 3967 16364 4005 16398
rect 4005 16364 4039 16398
rect 3933 16326 4039 16364
rect 3933 16292 3967 16326
rect 3967 16292 4005 16326
rect 4005 16292 4039 16326
rect 3933 16254 4039 16292
rect 3933 16220 3967 16254
rect 3967 16220 4005 16254
rect 4005 16220 4039 16254
rect 3933 16182 4039 16220
rect 3933 16148 3967 16182
rect 3967 16148 4005 16182
rect 4005 16148 4039 16182
rect 3933 16110 4039 16148
rect 3933 16076 3967 16110
rect 3967 16076 4005 16110
rect 4005 16076 4039 16110
rect 3933 16038 4039 16076
rect 3933 16004 3967 16038
rect 3967 16004 4005 16038
rect 4005 16004 4039 16038
rect 3933 15966 4039 16004
rect 3933 15932 3967 15966
rect 3967 15932 4005 15966
rect 4005 15932 4039 15966
rect 3933 15894 4039 15932
rect 3933 15860 3967 15894
rect 3967 15860 4005 15894
rect 4005 15860 4039 15894
rect 3933 15822 4039 15860
rect 3933 15788 3967 15822
rect 3967 15788 4005 15822
rect 4005 15788 4039 15822
rect 3933 15750 4039 15788
rect 3933 15716 3967 15750
rect 3967 15716 4005 15750
rect 4005 15716 4039 15750
rect 3933 15678 4039 15716
rect 3933 15644 3967 15678
rect 3967 15644 4005 15678
rect 4005 15644 4039 15678
rect 3933 15606 4039 15644
rect 3933 15572 3967 15606
rect 3967 15572 4005 15606
rect 4005 15572 4039 15606
rect 3933 15534 4039 15572
rect 3933 15500 3967 15534
rect 3967 15500 4005 15534
rect 4005 15500 4039 15534
rect 3933 15462 4039 15500
rect 3933 15428 3967 15462
rect 3967 15428 4005 15462
rect 4005 15428 4039 15462
rect 3933 15390 4039 15428
rect 3933 15356 3967 15390
rect 3967 15356 4005 15390
rect 4005 15356 4039 15390
rect 3933 15318 4039 15356
rect 3933 15284 3967 15318
rect 3967 15284 4005 15318
rect 4005 15284 4039 15318
rect 3933 15246 4039 15284
rect 3933 15212 3967 15246
rect 3967 15212 4005 15246
rect 4005 15212 4039 15246
rect 3933 15174 4039 15212
rect 3933 15140 3967 15174
rect 3967 15140 4005 15174
rect 4005 15140 4039 15174
rect 3933 15102 4039 15140
rect 3933 15068 3967 15102
rect 3967 15068 4005 15102
rect 4005 15068 4039 15102
rect 3933 15030 4039 15068
rect 3933 14996 3967 15030
rect 3967 14996 4005 15030
rect 4005 14996 4039 15030
rect 3933 14958 4039 14996
rect 3933 14924 3967 14958
rect 3967 14924 4005 14958
rect 4005 14924 4039 14958
rect 995 14852 1029 14886
rect 1029 14852 1067 14886
rect 1067 14852 1101 14886
rect 3933 14886 4039 14924
rect 995 14814 1101 14852
rect 995 14780 1029 14814
rect 1029 14780 1067 14814
rect 1067 14780 1101 14814
rect 1168 14837 1202 14871
rect 1202 14837 1240 14871
rect 1240 14837 1274 14871
rect 1274 14837 1312 14871
rect 1312 14837 1346 14871
rect 1346 14837 1384 14871
rect 1384 14837 1418 14871
rect 1418 14837 1456 14871
rect 1456 14837 1490 14871
rect 1490 14837 1528 14871
rect 1528 14837 1562 14871
rect 1562 14837 1600 14871
rect 1600 14837 1634 14871
rect 1634 14837 1672 14871
rect 1672 14837 1706 14871
rect 1706 14837 1744 14871
rect 1744 14837 1778 14871
rect 1778 14837 1816 14871
rect 1816 14837 1850 14871
rect 1850 14837 1888 14871
rect 1888 14837 1922 14871
rect 1922 14837 1960 14871
rect 1960 14837 1994 14871
rect 1994 14837 2032 14871
rect 2032 14837 2066 14871
rect 2066 14837 2104 14871
rect 2104 14837 2138 14871
rect 2138 14837 2176 14871
rect 2176 14837 2210 14871
rect 2210 14837 2248 14871
rect 2248 14837 2282 14871
rect 2282 14837 2320 14871
rect 2320 14837 2354 14871
rect 2354 14837 2392 14871
rect 2392 14837 2426 14871
rect 2426 14837 2464 14871
rect 2464 14837 2498 14871
rect 2498 14837 2536 14871
rect 2536 14837 2570 14871
rect 2570 14837 2608 14871
rect 2608 14837 2642 14871
rect 2642 14837 2680 14871
rect 2680 14837 2714 14871
rect 2714 14837 2752 14871
rect 2752 14837 2786 14871
rect 2786 14837 2824 14871
rect 2824 14837 2858 14871
rect 2858 14837 2896 14871
rect 2896 14837 2930 14871
rect 2930 14837 2968 14871
rect 2968 14837 3002 14871
rect 3002 14837 3040 14871
rect 3040 14837 3074 14871
rect 3074 14837 3112 14871
rect 3112 14837 3146 14871
rect 3146 14837 3184 14871
rect 3184 14837 3218 14871
rect 3218 14837 3256 14871
rect 3256 14837 3290 14871
rect 3290 14837 3328 14871
rect 3328 14837 3362 14871
rect 3362 14837 3400 14871
rect 3400 14837 3434 14871
rect 3434 14837 3472 14871
rect 3472 14837 3506 14871
rect 3506 14837 3544 14871
rect 3544 14837 3578 14871
rect 3578 14837 3616 14871
rect 3616 14837 3650 14871
rect 3650 14837 3688 14871
rect 3688 14837 3722 14871
rect 3722 14837 3760 14871
rect 3760 14837 3794 14871
rect 3794 14837 3832 14871
rect 3832 14837 3866 14871
rect 1168 14799 3866 14837
rect 1168 14765 1202 14799
rect 1202 14765 1240 14799
rect 1240 14765 1274 14799
rect 1274 14765 1312 14799
rect 1312 14765 1346 14799
rect 1346 14765 1384 14799
rect 1384 14765 1418 14799
rect 1418 14765 1456 14799
rect 1456 14765 1490 14799
rect 1490 14765 1528 14799
rect 1528 14765 1562 14799
rect 1562 14765 1600 14799
rect 1600 14765 1634 14799
rect 1634 14765 1672 14799
rect 1672 14765 1706 14799
rect 1706 14765 1744 14799
rect 1744 14765 1778 14799
rect 1778 14765 1816 14799
rect 1816 14765 1850 14799
rect 1850 14765 1888 14799
rect 1888 14765 1922 14799
rect 1922 14765 1960 14799
rect 1960 14765 1994 14799
rect 1994 14765 2032 14799
rect 2032 14765 2066 14799
rect 2066 14765 2104 14799
rect 2104 14765 2138 14799
rect 2138 14765 2176 14799
rect 2176 14765 2210 14799
rect 2210 14765 2248 14799
rect 2248 14765 2282 14799
rect 2282 14765 2320 14799
rect 2320 14765 2354 14799
rect 2354 14765 2392 14799
rect 2392 14765 2426 14799
rect 2426 14765 2464 14799
rect 2464 14765 2498 14799
rect 2498 14765 2536 14799
rect 2536 14765 2570 14799
rect 2570 14765 2608 14799
rect 2608 14765 2642 14799
rect 2642 14765 2680 14799
rect 2680 14765 2714 14799
rect 2714 14765 2752 14799
rect 2752 14765 2786 14799
rect 2786 14765 2824 14799
rect 2824 14765 2858 14799
rect 2858 14765 2896 14799
rect 2896 14765 2930 14799
rect 2930 14765 2968 14799
rect 2968 14765 3002 14799
rect 3002 14765 3040 14799
rect 3040 14765 3074 14799
rect 3074 14765 3112 14799
rect 3112 14765 3146 14799
rect 3146 14765 3184 14799
rect 3184 14765 3218 14799
rect 3218 14765 3256 14799
rect 3256 14765 3290 14799
rect 3290 14765 3328 14799
rect 3328 14765 3362 14799
rect 3362 14765 3400 14799
rect 3400 14765 3434 14799
rect 3434 14765 3472 14799
rect 3472 14765 3506 14799
rect 3506 14765 3544 14799
rect 3544 14765 3578 14799
rect 3578 14765 3616 14799
rect 3616 14765 3650 14799
rect 3650 14765 3688 14799
rect 3688 14765 3722 14799
rect 3722 14765 3760 14799
rect 3760 14765 3794 14799
rect 3794 14765 3832 14799
rect 3832 14765 3866 14799
rect 3933 14852 3967 14886
rect 3967 14852 4005 14886
rect 4005 14852 4039 14886
rect 3933 14814 4039 14852
rect 3933 14780 3967 14814
rect 3967 14780 4005 14814
rect 4005 14780 4039 14814
<< metal1 >>
rect 983 17421 4051 17433
rect 983 17406 1168 17421
rect 983 14780 995 17406
rect 1101 17315 1168 17406
rect 3866 17406 4051 17421
rect 3866 17315 3933 17406
rect 1101 17303 3933 17315
rect 1101 14883 1113 17303
rect 3921 14883 3933 17303
rect 1101 14871 3933 14883
rect 1101 14780 1168 14871
rect 983 14765 1168 14780
rect 3866 14780 3933 14871
rect 4039 14780 4051 17406
rect 3866 14765 4051 14780
rect 983 14753 4051 14765
<< metal3 >>
rect 1525 16885 1681 16891
rect 1525 15301 1531 16885
rect 1675 16587 1681 16885
rect 3353 16885 3509 16891
rect 3353 16739 3359 16885
rect 1757 16733 3359 16739
rect 1757 16669 1877 16733
rect 1941 16669 2181 16733
rect 2245 16669 2485 16733
rect 2549 16669 2789 16733
rect 2853 16669 3093 16733
rect 3157 16669 3359 16733
rect 1757 16663 3359 16669
rect 1675 16581 3277 16587
rect 1675 16517 2029 16581
rect 2093 16517 2333 16581
rect 2397 16517 2637 16581
rect 2701 16517 2941 16581
rect 3005 16517 3277 16581
rect 1675 16511 3277 16517
rect 1675 16283 1681 16511
rect 3353 16435 3359 16663
rect 1757 16429 3359 16435
rect 1757 16365 1877 16429
rect 1941 16365 2181 16429
rect 2245 16365 2485 16429
rect 2549 16365 2789 16429
rect 2853 16365 3093 16429
rect 3157 16365 3359 16429
rect 1757 16359 3359 16365
rect 1675 16277 3277 16283
rect 1675 16213 2029 16277
rect 2093 16213 2333 16277
rect 2397 16213 2637 16277
rect 2701 16213 2941 16277
rect 3005 16213 3277 16277
rect 1675 16207 3277 16213
rect 1675 15979 1681 16207
rect 3353 16131 3359 16359
rect 1757 16125 3359 16131
rect 1757 16061 1877 16125
rect 1941 16061 2181 16125
rect 2245 16061 2485 16125
rect 2549 16061 2789 16125
rect 2853 16061 3093 16125
rect 3157 16061 3359 16125
rect 1757 16055 3359 16061
rect 1675 15973 3277 15979
rect 1675 15909 2029 15973
rect 2093 15909 2333 15973
rect 2397 15909 2637 15973
rect 2701 15909 2941 15973
rect 3005 15909 3277 15973
rect 1675 15903 3277 15909
rect 1675 15675 1681 15903
rect 3353 15827 3359 16055
rect 1757 15821 3359 15827
rect 1757 15757 1877 15821
rect 1941 15757 2181 15821
rect 2245 15757 2485 15821
rect 2549 15757 2789 15821
rect 2853 15757 3093 15821
rect 3157 15757 3359 15821
rect 1757 15751 3359 15757
rect 1675 15669 3277 15675
rect 1675 15605 2029 15669
rect 2093 15605 2333 15669
rect 2397 15605 2637 15669
rect 2701 15605 2941 15669
rect 3005 15605 3277 15669
rect 1675 15599 3277 15605
rect 1675 15301 1681 15599
rect 3353 15523 3359 15751
rect 1757 15517 3359 15523
rect 1757 15453 1877 15517
rect 1941 15453 2181 15517
rect 2245 15453 2485 15517
rect 2549 15453 2789 15517
rect 2853 15453 3093 15517
rect 3157 15453 3359 15517
rect 1757 15447 3359 15453
rect 1525 15295 1681 15301
rect 3353 15301 3359 15447
rect 3503 15301 3509 16885
rect 3353 15295 3509 15301
<< via3 >>
rect 1531 15301 1675 16885
rect 1877 16669 1941 16733
rect 2181 16669 2245 16733
rect 2485 16669 2549 16733
rect 2789 16669 2853 16733
rect 3093 16669 3157 16733
rect 2029 16517 2093 16581
rect 2333 16517 2397 16581
rect 2637 16517 2701 16581
rect 2941 16517 3005 16581
rect 1877 16365 1941 16429
rect 2181 16365 2245 16429
rect 2485 16365 2549 16429
rect 2789 16365 2853 16429
rect 3093 16365 3157 16429
rect 2029 16213 2093 16277
rect 2333 16213 2397 16277
rect 2637 16213 2701 16277
rect 2941 16213 3005 16277
rect 1877 16061 1941 16125
rect 2181 16061 2245 16125
rect 2485 16061 2549 16125
rect 2789 16061 2853 16125
rect 3093 16061 3157 16125
rect 2029 15909 2093 15973
rect 2333 15909 2397 15973
rect 2637 15909 2701 15973
rect 2941 15909 3005 15973
rect 1877 15757 1941 15821
rect 2181 15757 2245 15821
rect 2485 15757 2549 15821
rect 2789 15757 2853 15821
rect 3093 15757 3157 15821
rect 2029 15605 2093 15669
rect 2333 15605 2397 15669
rect 2637 15605 2701 15669
rect 2941 15605 3005 15669
rect 1877 15453 1941 15517
rect 2181 15453 2245 15517
rect 2485 15453 2549 15517
rect 2789 15453 2853 15517
rect 3093 15453 3157 15517
rect 3359 15301 3503 16885
<< metal4 >>
rect 1525 16885 1681 16891
rect 1525 16851 1531 16885
rect 1675 16851 1681 16885
rect 3353 16885 3509 16891
rect 3353 16851 3359 16885
rect 3503 16851 3509 16885
rect 1445 16531 1531 16615
rect 1675 16531 1681 16615
rect 1445 16211 1531 16295
rect 1675 16211 1681 16295
rect 1445 15891 1531 15975
rect 1675 15891 1681 15975
rect 1445 15571 1531 15655
rect 1675 15571 1681 15655
rect 1871 16733 1947 16777
rect 1871 16669 1877 16733
rect 1941 16669 1947 16733
rect 1871 16429 1947 16669
rect 1871 16365 1877 16429
rect 1941 16365 1947 16429
rect 1871 16125 1947 16365
rect 1871 16061 1877 16125
rect 1941 16061 1947 16125
rect 1871 15821 1947 16061
rect 1871 15757 1877 15821
rect 1941 15757 1947 15821
rect 1871 15517 1947 15757
rect 1871 15453 1877 15517
rect 1941 15453 1947 15517
rect 1871 15409 1947 15453
rect 2023 16581 2099 16777
rect 2023 16517 2029 16581
rect 2093 16517 2099 16581
rect 2023 16277 2099 16517
rect 2023 16213 2029 16277
rect 2093 16213 2099 16277
rect 2023 15973 2099 16213
rect 2023 15909 2029 15973
rect 2093 15909 2099 15973
rect 2023 15669 2099 15909
rect 2023 15605 2029 15669
rect 2093 15605 2099 15669
rect 2023 15409 2099 15605
rect 2175 16733 2251 16777
rect 2175 16669 2181 16733
rect 2245 16669 2251 16733
rect 2175 16429 2251 16669
rect 2175 16365 2181 16429
rect 2245 16365 2251 16429
rect 2175 16125 2251 16365
rect 2175 16061 2181 16125
rect 2245 16061 2251 16125
rect 2175 15821 2251 16061
rect 2175 15757 2181 15821
rect 2245 15757 2251 15821
rect 2175 15517 2251 15757
rect 2175 15453 2181 15517
rect 2245 15453 2251 15517
rect 2175 15409 2251 15453
rect 2327 16581 2403 16777
rect 2327 16517 2333 16581
rect 2397 16517 2403 16581
rect 2327 16277 2403 16517
rect 2327 16213 2333 16277
rect 2397 16213 2403 16277
rect 2327 15973 2403 16213
rect 2327 15909 2333 15973
rect 2397 15909 2403 15973
rect 2327 15669 2403 15909
rect 2327 15605 2333 15669
rect 2397 15605 2403 15669
rect 2327 15409 2403 15605
rect 2479 16733 2555 16777
rect 2479 16669 2485 16733
rect 2549 16669 2555 16733
rect 2479 16429 2555 16669
rect 2479 16365 2485 16429
rect 2549 16365 2555 16429
rect 2479 16125 2555 16365
rect 2479 16061 2485 16125
rect 2549 16061 2555 16125
rect 2479 15821 2555 16061
rect 2479 15757 2485 15821
rect 2549 15757 2555 15821
rect 2479 15517 2555 15757
rect 2479 15453 2485 15517
rect 2549 15453 2555 15517
rect 2479 15409 2555 15453
rect 2631 16581 2707 16777
rect 2631 16517 2637 16581
rect 2701 16517 2707 16581
rect 2631 16277 2707 16517
rect 2631 16213 2637 16277
rect 2701 16213 2707 16277
rect 2631 15973 2707 16213
rect 2631 15909 2637 15973
rect 2701 15909 2707 15973
rect 2631 15669 2707 15909
rect 2631 15605 2637 15669
rect 2701 15605 2707 15669
rect 2631 15409 2707 15605
rect 2783 16733 2859 16777
rect 2783 16669 2789 16733
rect 2853 16669 2859 16733
rect 2783 16429 2859 16669
rect 2783 16365 2789 16429
rect 2853 16365 2859 16429
rect 2783 16125 2859 16365
rect 2783 16061 2789 16125
rect 2853 16061 2859 16125
rect 2783 15821 2859 16061
rect 2783 15757 2789 15821
rect 2853 15757 2859 15821
rect 2783 15517 2859 15757
rect 2783 15453 2789 15517
rect 2853 15453 2859 15517
rect 2783 15409 2859 15453
rect 2935 16581 3011 16777
rect 2935 16517 2941 16581
rect 3005 16517 3011 16581
rect 2935 16277 3011 16517
rect 2935 16213 2941 16277
rect 3005 16213 3011 16277
rect 2935 15973 3011 16213
rect 2935 15909 2941 15973
rect 3005 15909 3011 15973
rect 2935 15669 3011 15909
rect 2935 15605 2941 15669
rect 3005 15605 3011 15669
rect 2935 15409 3011 15605
rect 3087 16733 3163 16777
rect 3087 16669 3093 16733
rect 3157 16669 3163 16733
rect 3087 16429 3163 16669
rect 3087 16365 3093 16429
rect 3157 16365 3163 16429
rect 3087 16125 3163 16365
rect 3087 16061 3093 16125
rect 3157 16061 3163 16125
rect 3087 15821 3163 16061
rect 3087 15757 3093 15821
rect 3157 15757 3163 15821
rect 3087 15517 3163 15757
rect 3087 15453 3093 15517
rect 3157 15453 3163 15517
rect 3087 15409 3163 15453
rect 3353 16531 3359 16615
rect 3503 16531 3589 16615
rect 3353 16211 3359 16295
rect 3503 16211 3589 16295
rect 3353 15891 3359 15975
rect 3503 15891 3589 15975
rect 3353 15571 3359 15655
rect 3503 15571 3589 15655
rect 1525 15301 1531 15335
rect 1675 15301 1681 15335
rect 1525 15295 1681 15301
rect 3353 15301 3359 15335
rect 3503 15301 3509 15335
rect 3353 15295 3509 15301
<< via4 >>
rect 1445 16615 1531 16851
rect 1531 16615 1675 16851
rect 1675 16615 1681 16851
rect 1445 16295 1531 16531
rect 1531 16295 1675 16531
rect 1675 16295 1681 16531
rect 1445 15975 1531 16211
rect 1531 15975 1675 16211
rect 1675 15975 1681 16211
rect 1445 15655 1531 15891
rect 1531 15655 1675 15891
rect 1675 15655 1681 15891
rect 1445 15335 1531 15571
rect 1531 15335 1675 15571
rect 1675 15335 1681 15571
rect 3353 16615 3359 16851
rect 3359 16615 3503 16851
rect 3503 16615 3589 16851
rect 3353 16295 3359 16531
rect 3359 16295 3503 16531
rect 3503 16295 3589 16531
rect 3353 15975 3359 16211
rect 3359 15975 3503 16211
rect 3503 15975 3589 16211
rect 3353 15655 3359 15891
rect 3359 15655 3503 15891
rect 3503 15655 3589 15891
rect 3353 15335 3359 15571
rect 3359 15335 3503 15571
rect 3503 15335 3589 15571
<< metal5 >>
rect 1152 16851 1723 16875
rect 1152 16615 1445 16851
rect 1681 16615 1723 16851
rect 1152 16531 1723 16615
rect 1152 16295 1445 16531
rect 1681 16295 1723 16531
rect 1152 16211 1723 16295
rect 1152 15975 1445 16211
rect 1681 15975 1723 16211
rect 1152 15891 1723 15975
rect 1152 15655 1445 15891
rect 1681 15655 1723 15891
rect 1152 15571 1723 15655
rect 1152 15335 1445 15571
rect 1681 15335 1723 15571
rect 1152 15311 1723 15335
rect 3311 16851 3886 16875
rect 3311 16615 3353 16851
rect 3589 16615 3886 16851
rect 3311 16531 3886 16615
rect 3311 16295 3353 16531
rect 3589 16295 3886 16531
rect 3311 16211 3886 16295
rect 3311 15975 3353 16211
rect 3589 15975 3886 16211
rect 3311 15891 3886 15975
rect 3311 15655 3353 15891
rect 3589 15655 3886 15891
rect 3311 15571 3886 15655
rect 3311 15335 3353 15571
rect 3589 15335 3886 15571
rect 3311 15311 3886 15335
<< labels >>
flabel metal5 s 1152 15311 1192 16875 2 FreeSans 2000 0 0 0 in
port 1 nsew
flabel metal5 s 3846 15311 3886 16875 2 FreeSans 2000 0 0 0 out
port 2 nsew
flabel metal1 s 2389 14771 2480 14858 2 FreeSans 2000 0 0 0 gnd
port 3 nsew
<< properties >>
string device primitive
<< end >>
