* NGSPICE file created from LNA_final.ext - technology: sky130A

.subckt LNA_final Vgg_1v2 Vdd_1v8 Gnd
XMOM_capacitor_0 Vdd_1v8 MOM_capacitor_0/out Gnd MOM_capacitor
X0 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X21 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X24 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X28 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X31 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X34 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X38 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X41 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X42 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X45 a_n27544_n39610# a_n12387_n39359# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=1e+07u
X46 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X48 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X49 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X50 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X53 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X56 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X57 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X60 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X69 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X70 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 Vgg_1v2 a_n27544_n39610# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X71 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X72 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X73 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X74 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X79 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X83 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 Gnd MOM_capacitor_0/out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X85 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X86 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X88 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X93 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X94 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X98 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X100 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 Gnd MOM_capacitor_0/out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X104 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X105 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X106 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X107 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X109 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X110 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X120 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X123 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X124 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X126 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 a_n12387_n39359# m4_38188_n46509# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X129 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X130 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X133 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X135 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X136 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X143 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X144 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X145 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X146 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X147 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X149 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X150 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X151 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X153 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X163 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X164 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X165 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X167 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X169 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X171 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X172 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X173 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X175 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X176 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X177 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X178 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X179 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X180 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X181 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X183 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X185 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X186 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X188 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X189 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X190 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X191 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X193 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X195 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X196 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X197 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X198 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X201 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X202 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X203 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X207 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X208 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X209 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X213 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X214 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X215 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X216 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X217 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X218 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X219 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X222 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X223 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X224 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X225 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D0 Gnd Vdd_1v8 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X226 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X228 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X229 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X230 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X231 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X232 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X234 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X235 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X236 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X237 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X239 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X241 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X245 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X246 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X247 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

