* NGSPICE file created from VGA_gainCellv3.ext - technology: sky130A

X0 a_n2543_2314# Vctrl.t0 Vdd.t29 gnd.t69 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n2543_2314# gate.t0 out.t29 gnd.t105 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 Vdd.t28 Vctrl.t1 a_n2543_2314# gnd.t68 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_n2543_2314# Vctrl.t2 Vdd.t27 gnd.t67 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 out.t28 gate.t1 a_n2543_2314# gnd.t28 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_n2543_2314# gate.t2 out.t27 gnd.t106 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 out.t26 gate.t3 a_n2543_2314# gnd.t109 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_n2543_2314# Vctrl.t3 Vdd.t26 gnd.t66 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 Vdd.t25 Vctrl.t4 a_n2543_2314# gnd.t65 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 Vdd.t24 Vctrl.t5 a_n2543_2314# gnd.t64 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 out.t25 gate.t4 a_n2543_2314# gnd.t108 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 out.t24 gate.t5 a_n2543_2314# gnd.t103 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_n2543_2314# gate.t6 out.t23 gnd.t104 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_n2543_2314# gate.t7 out.t22 gnd.t29 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 a_n2543_2314# Vctrl.t6 Vdd.t23 gnd.t63 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_n2543_2314# Vctrl.t7 Vdd.t22 gnd.t62 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_n2543_2314# gate.t8 out.t21 gnd.t0 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 a_n2543_2314# Vctrl.t8 Vdd.t21 gnd.t61 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 Vdd.t20 Vctrl.t9 a_n2543_2314# gnd.t60 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 gnd.t101 in.t0 a_n2543_2314# gnd.t100 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 Vdd.t19 Vctrl.t10 a_n2543_2314# gnd.t59 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 gnd.t111 in.t1 a_n2543_2314# gnd.t110 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 a_n2543_2314# in.t2 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_n2543_2314# in.t3 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 gnd.t88 in.t4 a_n2543_2314# gnd.t87 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 a_n2543_2314# in.t5 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_n2543_2314# Vctrl.t11 Vdd.t18 gnd.t58 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 a_n2543_2314# gate.t9 out.t20 gnd.t23 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 gnd.t6 in.t6 a_n2543_2314# gnd.t5 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 a_n2543_2314# in.t7 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 a_n2543_2314# gate.t10 out.t19 gnd.t107 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 a_n2543_2314# Vctrl.t12 Vdd.t17 gnd.t57 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X32 gnd.t27 in.t8 a_n2543_2314# gnd.t26 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 gnd.t77 in.t9 a_n2543_2314# gnd.t76 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X34 a_n2543_2314# in.t10 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 a_n2543_2314# in.t11 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 gnd.t34 in.t12 a_n2543_2314# gnd.t33 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 Vdd.t16 Vctrl.t13 a_n2543_2314# gnd.t56 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 Vdd.t15 Vctrl.t14 a_n2543_2314# gnd.t55 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 gnd.t10 in.t13 a_n2543_2314# gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 Vdd.t14 Vctrl.t15 a_n2543_2314# gnd.t54 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 Vdd.t13 Vctrl.t16 a_n2543_2314# gnd.t53 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 a_n2543_2314# gate.t11 out.t18 gnd.t30 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X43 a_n2543_2314# in.t14 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X44 gnd.t90 in.t15 a_n2543_2314# gnd.t89 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X45 out.t17 gate.t12 a_n2543_2314# gnd.t39 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X46 a_n2543_2314# gate.t13 out.t16 gnd.t38 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X47 gnd.t86 in.t16 a_n2543_2314# gnd.t85 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X48 a_n2543_2314# in.t17 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X49 gnd.t75 in.t18 a_n2543_2314# gnd.t74 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X50 a_n2543_2314# in.t19 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X51 a_n2543_2314# in.t20 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X52 a_n2543_2314# in.t21 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X53 gnd.t36 in.t22 a_n2543_2314# gnd.t35 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X54 gnd.t119 in.t23 a_n2543_2314# gnd.t118 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X55 a_n2543_2314# in.t24 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X56 a_n2543_2314# in.t25 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X57 gnd.t114 in.t26 a_n2543_2314# gnd.t113 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X58 gnd.t14 in.t27 a_n2543_2314# gnd.t13 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X59 a_n2543_2314# gate.t14 out.t15 gnd.t37 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X60 out.t14 gate.t15 a_n2543_2314# gnd.t1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X61 Vdd.t12 Vctrl.t17 a_n2543_2314# gnd.t52 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X62 out.t13 gate.t16 a_n2543_2314# gnd.t71 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X63 out.t12 gate.t17 a_n2543_2314# gnd.t112 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X64 a_n2543_2314# in.t28 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X65 a_n2543_2314# gate.t18 out.t11 gnd.t102 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X66 Vdd.t11 Vctrl.t18 a_n2543_2314# gnd.t51 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X67 out.t10 gate.t19 a_n2543_2314# gnd.t15 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X68 Vdd.t10 Vctrl.t19 a_n2543_2314# gnd.t50 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X69 a_n2543_2314# Vctrl.t20 Vdd.t9 gnd.t49 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X70 a_n2543_2314# gate.t20 out.t9 gnd.t82 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X71 a_n2543_2314# Vctrl.t21 Vdd.t8 gnd.t48 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X72 out.t8 gate.t21 a_n2543_2314# gnd.t70 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X73 a_n2543_2314# Vctrl.t22 Vdd.t7 gnd.t47 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X74 out.t7 gate.t22 a_n2543_2314# gnd.t4 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X75 Vdd.t6 Vctrl.t23 a_n2543_2314# gnd.t46 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X76 a_n2543_2314# gate.t23 out.t6 gnd.t2 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X77 a_n2543_2314# Vctrl.t24 Vdd.t5 gnd.t45 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X78 Vdd.t4 Vctrl.t25 a_n2543_2314# gnd.t44 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X79 Vdd.t3 Vctrl.t26 a_n2543_2314# gnd.t43 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X80 a_n2543_2314# Vctrl.t27 Vdd.t2 gnd.t42 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X81 out.t5 gate.t24 a_n2543_2314# gnd.t73 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X82 a_n2543_2314# gate.t25 out.t4 gnd.t72 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X83 a_n2543_2314# in.t29 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X84 a_n2543_2314# Vctrl.t28 Vdd.t1 gnd.t41 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X85 a_n2543_2314# Vctrl.t29 Vdd.t0 gnd.t40 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X86 out.t3 gate.t26 a_n2543_2314# gnd.t115 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X87 a_n2543_2314# gate.t27 out.t2 gnd.t99 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X88 out.t1 gate.t28 a_n2543_2314# gnd.t3 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X89 out.t0 gate.t29 a_n2543_2314# gnd.t16 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 Vctrl.n28 Vctrl.t15 179.593
R1 Vctrl.n28 Vctrl.t29 179.476
R2 Vctrl.n29 Vctrl.t25 170.306
R3 Vctrl.n26 Vctrl.t20 170.306
R4 Vctrl.n33 Vctrl.t13 170.306
R5 Vctrl.n24 Vctrl.t27 170.306
R6 Vctrl.n37 Vctrl.t23 170.306
R7 Vctrl.n22 Vctrl.t0 170.306
R8 Vctrl.n41 Vctrl.t4 170.306
R9 Vctrl.n20 Vctrl.t11 170.306
R10 Vctrl.n45 Vctrl.t10 170.306
R11 Vctrl.n18 Vctrl.t22 170.306
R12 Vctrl.n49 Vctrl.t18 170.306
R13 Vctrl.n16 Vctrl.t21 170.306
R14 Vctrl.n53 Vctrl.t17 170.306
R15 Vctrl.n14 Vctrl.t3 170.306
R16 Vctrl.n57 Vctrl.t14 170.306
R17 Vctrl.n12 Vctrl.t6 170.306
R18 Vctrl.n61 Vctrl.t1 170.306
R19 Vctrl.n10 Vctrl.t24 170.306
R20 Vctrl.n65 Vctrl.t26 170.306
R21 Vctrl.n8 Vctrl.t12 170.306
R22 Vctrl.n69 Vctrl.t16 170.306
R23 Vctrl.n6 Vctrl.t8 170.306
R24 Vctrl.n73 Vctrl.t19 170.306
R25 Vctrl.n4 Vctrl.t7 170.306
R26 Vctrl.n77 Vctrl.t9 170.306
R27 Vctrl.n2 Vctrl.t2 170.306
R28 Vctrl.n81 Vctrl.t5 170.306
R29 Vctrl.n0 Vctrl.t28 170.306
R30 Vctrl.n27 Vctrl.n26 8.764
R31 Vctrl.n25 Vctrl.n24 8.764
R32 Vctrl.n23 Vctrl.n22 8.764
R33 Vctrl.n21 Vctrl.n20 8.764
R34 Vctrl.n19 Vctrl.n18 8.764
R35 Vctrl.n17 Vctrl.n16 8.764
R36 Vctrl.n15 Vctrl.n14 8.764
R37 Vctrl.n13 Vctrl.n12 8.764
R38 Vctrl.n11 Vctrl.n10 8.764
R39 Vctrl.n9 Vctrl.n8 8.764
R40 Vctrl.n7 Vctrl.n6 8.764
R41 Vctrl.n5 Vctrl.n4 8.764
R42 Vctrl.n3 Vctrl.n2 8.764
R43 Vctrl.n1 Vctrl.n0 8.764
R44 Vctrl.n82 Vctrl.n81 8.764
R45 Vctrl.n78 Vctrl.n77 8.764
R46 Vctrl.n74 Vctrl.n73 8.764
R47 Vctrl.n70 Vctrl.n69 8.764
R48 Vctrl.n66 Vctrl.n65 8.764
R49 Vctrl.n62 Vctrl.n61 8.764
R50 Vctrl.n58 Vctrl.n57 8.764
R51 Vctrl.n54 Vctrl.n53 8.764
R52 Vctrl.n50 Vctrl.n49 8.764
R53 Vctrl.n46 Vctrl.n45 8.764
R54 Vctrl.n42 Vctrl.n41 8.764
R55 Vctrl.n38 Vctrl.n37 8.764
R56 Vctrl.n34 Vctrl.n33 8.764
R57 Vctrl.n30 Vctrl.n29 8.764
R58 Vctrl.n84 Vctrl.n1 4.65
R59 Vctrl.n83 Vctrl.n82 4.65
R60 Vctrl.n80 Vctrl.n3 4.65
R61 Vctrl.n79 Vctrl.n78 4.65
R62 Vctrl.n76 Vctrl.n5 4.65
R63 Vctrl.n75 Vctrl.n74 4.65
R64 Vctrl.n72 Vctrl.n7 4.65
R65 Vctrl.n71 Vctrl.n70 4.65
R66 Vctrl.n68 Vctrl.n9 4.65
R67 Vctrl.n67 Vctrl.n66 4.65
R68 Vctrl.n64 Vctrl.n11 4.65
R69 Vctrl.n63 Vctrl.n62 4.65
R70 Vctrl.n60 Vctrl.n13 4.65
R71 Vctrl.n59 Vctrl.n58 4.65
R72 Vctrl.n56 Vctrl.n15 4.65
R73 Vctrl.n55 Vctrl.n54 4.65
R74 Vctrl.n52 Vctrl.n17 4.65
R75 Vctrl.n51 Vctrl.n50 4.65
R76 Vctrl.n48 Vctrl.n19 4.65
R77 Vctrl.n47 Vctrl.n46 4.65
R78 Vctrl.n44 Vctrl.n21 4.65
R79 Vctrl.n43 Vctrl.n42 4.65
R80 Vctrl.n40 Vctrl.n23 4.65
R81 Vctrl.n39 Vctrl.n38 4.65
R82 Vctrl.n36 Vctrl.n25 4.65
R83 Vctrl.n35 Vctrl.n34 4.65
R84 Vctrl.n32 Vctrl.n27 4.65
R85 Vctrl.n31 Vctrl.n30 4.65
R86 Vctrl.n31 Vctrl.n28 2.744
R87 Vctrl Vctrl.n84 2.669
R88 Vctrl.n83 Vctrl.n80 0.6
R89 Vctrl.n79 Vctrl.n76 0.6
R90 Vctrl.n75 Vctrl.n72 0.6
R91 Vctrl.n71 Vctrl.n68 0.6
R92 Vctrl.n67 Vctrl.n64 0.6
R93 Vctrl.n63 Vctrl.n60 0.6
R94 Vctrl.n59 Vctrl.n56 0.6
R95 Vctrl.n55 Vctrl.n52 0.6
R96 Vctrl.n51 Vctrl.n48 0.6
R97 Vctrl.n47 Vctrl.n44 0.6
R98 Vctrl.n43 Vctrl.n40 0.6
R99 Vctrl.n39 Vctrl.n36 0.6
R100 Vctrl.n35 Vctrl.n32 0.6
R101 Vctrl.n84 Vctrl.n83 0.2
R102 Vctrl.n80 Vctrl.n79 0.2
R103 Vctrl.n76 Vctrl.n75 0.2
R104 Vctrl.n72 Vctrl.n71 0.2
R105 Vctrl.n68 Vctrl.n67 0.2
R106 Vctrl.n64 Vctrl.n63 0.2
R107 Vctrl.n60 Vctrl.n59 0.2
R108 Vctrl.n56 Vctrl.n55 0.2
R109 Vctrl.n52 Vctrl.n51 0.2
R110 Vctrl.n48 Vctrl.n47 0.2
R111 Vctrl.n44 Vctrl.n43 0.2
R112 Vctrl.n40 Vctrl.n39 0.2
R113 Vctrl.n36 Vctrl.n35 0.2
R114 Vctrl.n32 Vctrl.n31 0.2
R115 Vdd.n0 Vdd.t0 23.571
R116 Vdd.n0 Vdd.t14 23.571
R117 Vdd.n9 Vdd.t9 23.571
R118 Vdd.n9 Vdd.t4 23.571
R119 Vdd.n18 Vdd.t2 23.571
R120 Vdd.n18 Vdd.t16 23.571
R121 Vdd.n27 Vdd.t29 23.571
R122 Vdd.n27 Vdd.t6 23.571
R123 Vdd.n36 Vdd.t18 23.571
R124 Vdd.n36 Vdd.t25 23.571
R125 Vdd.n45 Vdd.t7 23.571
R126 Vdd.n45 Vdd.t19 23.571
R127 Vdd.n54 Vdd.t8 23.571
R128 Vdd.n54 Vdd.t11 23.571
R129 Vdd.n63 Vdd.t26 23.571
R130 Vdd.n63 Vdd.t12 23.571
R131 Vdd.n72 Vdd.t23 23.571
R132 Vdd.n72 Vdd.t15 23.571
R133 Vdd.n81 Vdd.t5 23.571
R134 Vdd.n81 Vdd.t28 23.571
R135 Vdd.n90 Vdd.t17 23.571
R136 Vdd.n90 Vdd.t3 23.571
R137 Vdd.n99 Vdd.t21 23.571
R138 Vdd.n99 Vdd.t13 23.571
R139 Vdd.n108 Vdd.t22 23.571
R140 Vdd.n108 Vdd.t10 23.571
R141 Vdd.n117 Vdd.t27 23.571
R142 Vdd.n117 Vdd.t20 23.571
R143 Vdd.n126 Vdd.t1 23.571
R144 Vdd.n126 Vdd.t24 23.571
R145 Vdd.n15 Vdd.n10 8.032
R146 Vdd.n24 Vdd.n19 8.032
R147 Vdd.n33 Vdd.n28 8.032
R148 Vdd.n42 Vdd.n37 8.032
R149 Vdd.n51 Vdd.n46 8.032
R150 Vdd.n60 Vdd.n55 8.032
R151 Vdd.n69 Vdd.n64 8.032
R152 Vdd.n78 Vdd.n73 8.032
R153 Vdd.n87 Vdd.n82 8.032
R154 Vdd.n96 Vdd.n91 8.032
R155 Vdd.n105 Vdd.n100 8.032
R156 Vdd.n114 Vdd.n109 8.032
R157 Vdd.n123 Vdd.n118 8.032
R158 Vdd.n132 Vdd.n127 8.032
R159 Vdd.n6 Vdd.n1 8.031
R160 Vdd.n3 Vdd.n2 3.85
R161 Vdd.n12 Vdd.n11 3.85
R162 Vdd.n21 Vdd.n20 3.85
R163 Vdd.n30 Vdd.n29 3.85
R164 Vdd.n39 Vdd.n38 3.85
R165 Vdd.n48 Vdd.n47 3.85
R166 Vdd.n57 Vdd.n56 3.85
R167 Vdd.n66 Vdd.n65 3.85
R168 Vdd.n75 Vdd.n74 3.85
R169 Vdd.n84 Vdd.n83 3.85
R170 Vdd.n93 Vdd.n92 3.85
R171 Vdd.n102 Vdd.n101 3.85
R172 Vdd.n111 Vdd.n110 3.85
R173 Vdd.n120 Vdd.n119 3.85
R174 Vdd.n129 Vdd.n128 3.85
R175 Vdd.n1 Vdd.n0 1.601
R176 Vdd.n10 Vdd.n9 1.601
R177 Vdd.n19 Vdd.n18 1.601
R178 Vdd.n28 Vdd.n27 1.601
R179 Vdd.n37 Vdd.n36 1.601
R180 Vdd.n46 Vdd.n45 1.601
R181 Vdd.n55 Vdd.n54 1.601
R182 Vdd.n64 Vdd.n63 1.601
R183 Vdd.n73 Vdd.n72 1.601
R184 Vdd.n82 Vdd.n81 1.601
R185 Vdd.n91 Vdd.n90 1.601
R186 Vdd.n100 Vdd.n99 1.601
R187 Vdd.n109 Vdd.n108 1.601
R188 Vdd.n118 Vdd.n117 1.601
R189 Vdd.n127 Vdd.n126 1.601
R190 Vdd.n7 Vdd.n6 0.619
R191 Vdd.n16 Vdd.n15 0.618
R192 Vdd.n25 Vdd.n24 0.618
R193 Vdd.n34 Vdd.n33 0.618
R194 Vdd.n43 Vdd.n42 0.618
R195 Vdd.n52 Vdd.n51 0.618
R196 Vdd.n61 Vdd.n60 0.618
R197 Vdd.n70 Vdd.n69 0.618
R198 Vdd.n79 Vdd.n78 0.618
R199 Vdd.n88 Vdd.n87 0.618
R200 Vdd.n97 Vdd.n96 0.618
R201 Vdd.n106 Vdd.n105 0.618
R202 Vdd.n115 Vdd.n114 0.618
R203 Vdd.n124 Vdd.n123 0.618
R204 Vdd.n133 Vdd.n132 0.618
R205 Vdd.n135 Vdd.n134 0.616
R206 Vdd.n148 Vdd.n8 0.539
R207 Vdd.n147 Vdd.n17 0.539
R208 Vdd.n146 Vdd.n26 0.539
R209 Vdd.n145 Vdd.n35 0.539
R210 Vdd.n144 Vdd.n44 0.539
R211 Vdd.n143 Vdd.n53 0.539
R212 Vdd.n142 Vdd.n62 0.539
R213 Vdd.n141 Vdd.n71 0.539
R214 Vdd.n140 Vdd.n80 0.539
R215 Vdd.n139 Vdd.n89 0.539
R216 Vdd.n138 Vdd.n98 0.539
R217 Vdd.n137 Vdd.n107 0.539
R218 Vdd.n136 Vdd.n116 0.539
R219 Vdd.n135 Vdd.n125 0.539
R220 Vdd Vdd.n148 0.291
R221 Vdd.n6 Vdd.n5 0.098
R222 Vdd.n15 Vdd.n14 0.098
R223 Vdd.n24 Vdd.n23 0.098
R224 Vdd.n33 Vdd.n32 0.098
R225 Vdd.n42 Vdd.n41 0.098
R226 Vdd.n51 Vdd.n50 0.098
R227 Vdd.n60 Vdd.n59 0.098
R228 Vdd.n69 Vdd.n68 0.098
R229 Vdd.n78 Vdd.n77 0.098
R230 Vdd.n87 Vdd.n86 0.098
R231 Vdd.n96 Vdd.n95 0.098
R232 Vdd.n105 Vdd.n104 0.098
R233 Vdd.n114 Vdd.n113 0.098
R234 Vdd.n123 Vdd.n122 0.098
R235 Vdd.n132 Vdd.n131 0.098
R236 Vdd.n136 Vdd.n135 0.077
R237 Vdd.n137 Vdd.n136 0.077
R238 Vdd.n138 Vdd.n137 0.077
R239 Vdd.n139 Vdd.n138 0.077
R240 Vdd.n140 Vdd.n139 0.077
R241 Vdd.n141 Vdd.n140 0.077
R242 Vdd.n142 Vdd.n141 0.077
R243 Vdd.n143 Vdd.n142 0.077
R244 Vdd.n144 Vdd.n143 0.077
R245 Vdd.n145 Vdd.n144 0.077
R246 Vdd.n146 Vdd.n145 0.077
R247 Vdd.n147 Vdd.n146 0.077
R248 Vdd.n148 Vdd.n147 0.077
R249 Vdd.n8 Vdd.n7 0.037
R250 Vdd.n17 Vdd.n16 0.037
R251 Vdd.n26 Vdd.n25 0.037
R252 Vdd.n35 Vdd.n34 0.037
R253 Vdd.n44 Vdd.n43 0.037
R254 Vdd.n53 Vdd.n52 0.037
R255 Vdd.n62 Vdd.n61 0.037
R256 Vdd.n71 Vdd.n70 0.037
R257 Vdd.n80 Vdd.n79 0.037
R258 Vdd.n89 Vdd.n88 0.037
R259 Vdd.n98 Vdd.n97 0.037
R260 Vdd.n107 Vdd.n106 0.037
R261 Vdd.n116 Vdd.n115 0.037
R262 Vdd.n125 Vdd.n124 0.037
R263 Vdd.n134 Vdd.n133 0.037
R264 Vdd.n4 Vdd.n3 0.008
R265 Vdd.n13 Vdd.n12 0.008
R266 Vdd.n22 Vdd.n21 0.008
R267 Vdd.n31 Vdd.n30 0.008
R268 Vdd.n40 Vdd.n39 0.008
R269 Vdd.n49 Vdd.n48 0.008
R270 Vdd.n58 Vdd.n57 0.008
R271 Vdd.n67 Vdd.n66 0.008
R272 Vdd.n76 Vdd.n75 0.008
R273 Vdd.n85 Vdd.n84 0.008
R274 Vdd.n94 Vdd.n93 0.008
R275 Vdd.n103 Vdd.n102 0.008
R276 Vdd.n112 Vdd.n111 0.008
R277 Vdd.n121 Vdd.n120 0.008
R278 Vdd.n130 Vdd.n129 0.008
R279 Vdd.n5 Vdd.n4 0.001
R280 Vdd.n14 Vdd.n13 0.001
R281 Vdd.n23 Vdd.n22 0.001
R282 Vdd.n32 Vdd.n31 0.001
R283 Vdd.n41 Vdd.n40 0.001
R284 Vdd.n50 Vdd.n49 0.001
R285 Vdd.n59 Vdd.n58 0.001
R286 Vdd.n68 Vdd.n67 0.001
R287 Vdd.n77 Vdd.n76 0.001
R288 Vdd.n86 Vdd.n85 0.001
R289 Vdd.n95 Vdd.n94 0.001
R290 Vdd.n104 Vdd.n103 0.001
R291 Vdd.n113 Vdd.n112 0.001
R292 Vdd.n122 Vdd.n121 0.001
R293 Vdd.n131 Vdd.n130 0.001
R294 gnd.n285 gnd.n284 380.388
R295 gnd.n6 gnd.n5 380.388
R296 gnd.n565 gnd.n564 378.245
R297 gnd.n626 gnd.n625 378.245
R298 gnd.n630 gnd.n626 378.245
R299 gnd.n567 gnd.n566 295.014
R300 gnd.n287 gnd.n286 294.881
R301 gnd.n8 gnd.n7 294.881
R302 gnd.n291 gnd.n290 292.5
R303 gnd.n298 gnd.n297 292.5
R304 gnd.n309 gnd.n308 292.5
R305 gnd.n305 gnd.n304 292.5
R306 gnd.n316 gnd.n315 292.5
R307 gnd.n323 gnd.n322 292.5
R308 gnd.n330 gnd.n329 292.5
R309 gnd.n331 gnd.n330 292.5
R310 gnd.n338 gnd.n337 292.5
R311 gnd.n339 gnd.n338 292.5
R312 gnd.n346 gnd.n345 292.5
R313 gnd.t24 gnd.n346 292.5
R314 gnd.n353 gnd.n352 292.5
R315 gnd.n354 gnd.n353 292.5
R316 gnd.n361 gnd.n360 292.5
R317 gnd.n362 gnd.n361 292.5
R318 gnd.n369 gnd.n368 292.5
R319 gnd.n370 gnd.n369 292.5
R320 gnd.n376 gnd.n375 292.5
R321 gnd.n377 gnd.n376 292.5
R322 gnd.n384 gnd.n383 292.5
R323 gnd.n385 gnd.n384 292.5
R324 gnd.n392 gnd.n391 292.5
R325 gnd.n393 gnd.n392 292.5
R326 gnd.n400 gnd.n399 292.5
R327 gnd.n401 gnd.n400 292.5
R328 gnd.n408 gnd.n407 292.5
R329 gnd.n409 gnd.n408 292.5
R330 gnd.n416 gnd.n415 292.5
R331 gnd.n417 gnd.n416 292.5
R332 gnd.n424 gnd.n423 292.5
R333 gnd.n425 gnd.n424 292.5
R334 gnd.n432 gnd.n431 292.5
R335 gnd.n433 gnd.n432 292.5
R336 gnd.n158 gnd.n157 292.5
R337 gnd.n159 gnd.n158 292.5
R338 gnd.n153 gnd.n152 292.5
R339 gnd.n154 gnd.n153 292.5
R340 gnd.n145 gnd.n144 292.5
R341 gnd.n146 gnd.n145 292.5
R342 gnd.n137 gnd.n136 292.5
R343 gnd.n138 gnd.n137 292.5
R344 gnd.n129 gnd.n128 292.5
R345 gnd.n130 gnd.n129 292.5
R346 gnd.n121 gnd.n120 292.5
R347 gnd.n122 gnd.n121 292.5
R348 gnd.n113 gnd.n112 292.5
R349 gnd.n114 gnd.n113 292.5
R350 gnd.n105 gnd.n104 292.5
R351 gnd.n106 gnd.n105 292.5
R352 gnd.n97 gnd.n96 292.5
R353 gnd.n98 gnd.n97 292.5
R354 gnd.n90 gnd.n89 292.5
R355 gnd.n91 gnd.n90 292.5
R356 gnd.n82 gnd.n81 292.5
R357 gnd.n83 gnd.n82 292.5
R358 gnd.n74 gnd.n73 292.5
R359 gnd.n75 gnd.n74 292.5
R360 gnd.n67 gnd.n66 292.5
R361 gnd.t26 gnd.n67 292.5
R362 gnd.n59 gnd.n58 292.5
R363 gnd.n60 gnd.n59 292.5
R364 gnd.n51 gnd.n50 292.5
R365 gnd.n52 gnd.n51 292.5
R366 gnd.n44 gnd.n43 292.5
R367 gnd.n37 gnd.n36 292.5
R368 gnd.n30 gnd.n29 292.5
R369 gnd.n26 gnd.n25 292.5
R370 gnd.n19 gnd.n18 292.5
R371 gnd.n12 gnd.n11 292.5
R372 gnd.n68 gnd.t26 292.5
R373 gnd.n347 gnd.t24 292.5
R374 gnd.n14 gnd.n13 292.5
R375 gnd.n13 gnd.n12 292.5
R376 gnd.n21 gnd.n20 292.5
R377 gnd.n20 gnd.n19 292.5
R378 gnd.n28 gnd.n27 292.5
R379 gnd.n27 gnd.n26 292.5
R380 gnd.n32 gnd.n31 292.5
R381 gnd.n31 gnd.n30 292.5
R382 gnd.n39 gnd.n38 292.5
R383 gnd.n38 gnd.n37 292.5
R384 gnd.n46 gnd.n45 292.5
R385 gnd.n45 gnd.n44 292.5
R386 gnd.n54 gnd.n53 292.5
R387 gnd.n53 gnd.n52 292.5
R388 gnd.n62 gnd.n61 292.5
R389 gnd.n61 gnd.n60 292.5
R390 gnd.n69 gnd.n68 292.5
R391 gnd.n77 gnd.n76 292.5
R392 gnd.n76 gnd.n75 292.5
R393 gnd.n85 gnd.n84 292.5
R394 gnd.n84 gnd.n83 292.5
R395 gnd.n93 gnd.n92 292.5
R396 gnd.n92 gnd.n91 292.5
R397 gnd.n100 gnd.n99 292.5
R398 gnd.n99 gnd.n98 292.5
R399 gnd.n108 gnd.n107 292.5
R400 gnd.n107 gnd.n106 292.5
R401 gnd.n116 gnd.n115 292.5
R402 gnd.n115 gnd.n114 292.5
R403 gnd.n124 gnd.n123 292.5
R404 gnd.n123 gnd.n122 292.5
R405 gnd.n132 gnd.n131 292.5
R406 gnd.n131 gnd.n130 292.5
R407 gnd.n140 gnd.n139 292.5
R408 gnd.n139 gnd.n138 292.5
R409 gnd.n148 gnd.n147 292.5
R410 gnd.n147 gnd.n146 292.5
R411 gnd.n156 gnd.n155 292.5
R412 gnd.n155 gnd.n154 292.5
R413 gnd.n161 gnd.n160 292.5
R414 gnd.n160 gnd.n159 292.5
R415 gnd.n435 gnd.n434 292.5
R416 gnd.n434 gnd.n433 292.5
R417 gnd.n427 gnd.n426 292.5
R418 gnd.n426 gnd.n425 292.5
R419 gnd.n419 gnd.n418 292.5
R420 gnd.n418 gnd.n417 292.5
R421 gnd.n411 gnd.n410 292.5
R422 gnd.n410 gnd.n409 292.5
R423 gnd.n403 gnd.n402 292.5
R424 gnd.n402 gnd.n401 292.5
R425 gnd.n395 gnd.n394 292.5
R426 gnd.n394 gnd.n393 292.5
R427 gnd.n387 gnd.n386 292.5
R428 gnd.n386 gnd.n385 292.5
R429 gnd.n379 gnd.n378 292.5
R430 gnd.n378 gnd.n377 292.5
R431 gnd.n372 gnd.n371 292.5
R432 gnd.n371 gnd.n370 292.5
R433 gnd.n364 gnd.n363 292.5
R434 gnd.n363 gnd.n362 292.5
R435 gnd.n356 gnd.n355 292.5
R436 gnd.n355 gnd.n354 292.5
R437 gnd.n348 gnd.n347 292.5
R438 gnd.n341 gnd.n340 292.5
R439 gnd.n340 gnd.n339 292.5
R440 gnd.n333 gnd.n332 292.5
R441 gnd.n332 gnd.n331 292.5
R442 gnd.n325 gnd.n324 292.5
R443 gnd.n324 gnd.n323 292.5
R444 gnd.n318 gnd.n317 292.5
R445 gnd.n317 gnd.n316 292.5
R446 gnd.n307 gnd.n306 292.5
R447 gnd.n306 gnd.n305 292.5
R448 gnd.n311 gnd.n310 292.5
R449 gnd.n310 gnd.n309 292.5
R450 gnd.n300 gnd.n299 292.5
R451 gnd.n299 gnd.n298 292.5
R452 gnd.n293 gnd.n292 292.5
R453 gnd.n292 gnd.n291 292.5
R454 gnd.n628 gnd.n627 292.5
R455 gnd.n632 gnd.n631 292.5
R456 gnd.n636 gnd.n635 292.5
R457 gnd.n640 gnd.n639 292.5
R458 gnd.n644 gnd.n643 292.5
R459 gnd.n648 gnd.n647 292.5
R460 gnd.n649 gnd.n648 292.5
R461 gnd.n653 gnd.n652 292.5
R462 gnd.n657 gnd.n656 292.5
R463 gnd.n663 gnd.n662 292.5
R464 gnd.n664 gnd.n663 292.5
R465 gnd.n668 gnd.n667 292.5
R466 gnd.n669 gnd.n668 292.5
R467 gnd.n673 gnd.n672 292.5
R468 gnd.n678 gnd.n677 292.5
R469 gnd.n679 gnd.n678 292.5
R470 gnd.n683 gnd.n682 292.5
R471 gnd.n688 gnd.n687 292.5
R472 gnd.n689 gnd.n688 292.5
R473 gnd.n693 gnd.n692 292.5
R474 gnd.n694 gnd.n693 292.5
R475 gnd.n698 gnd.n697 292.5
R476 gnd.n699 gnd.n698 292.5
R477 gnd.n703 gnd.n702 292.5
R478 gnd.n704 gnd.n703 292.5
R479 gnd.n708 gnd.n707 292.5
R480 gnd.n709 gnd.n708 292.5
R481 gnd.n713 gnd.n712 292.5
R482 gnd.n714 gnd.n713 292.5
R483 gnd.n718 gnd.n717 292.5
R484 gnd.n719 gnd.n718 292.5
R485 gnd.n723 gnd.n722 292.5
R486 gnd.n724 gnd.n723 292.5
R487 gnd.n728 gnd.n727 292.5
R488 gnd.n729 gnd.n728 292.5
R489 gnd.n733 gnd.n732 292.5
R490 gnd.n737 gnd.n736 292.5
R491 gnd.n741 gnd.n740 292.5
R492 gnd.n748 gnd.n747 292.5
R493 gnd.n749 gnd.n748 292.5
R494 gnd.n753 gnd.n752 292.5
R495 gnd.n754 gnd.n753 292.5
R496 gnd.n758 gnd.n757 292.5
R497 gnd.n763 gnd.n762 292.5
R498 gnd.n764 gnd.n763 292.5
R499 gnd.n768 gnd.n767 292.5
R500 gnd.n769 gnd.n768 292.5
R501 gnd.n773 gnd.n772 292.5
R502 gnd.n774 gnd.n773 292.5
R503 gnd.n778 gnd.n777 292.5
R504 gnd.n779 gnd.n778 292.5
R505 gnd.n783 gnd.n782 292.5
R506 gnd.n788 gnd.n787 292.5
R507 gnd.n789 gnd.n788 292.5
R508 gnd.n793 gnd.n792 292.5
R509 gnd.n797 gnd.n796 292.5
R510 gnd.n803 gnd.n802 292.5
R511 gnd.n804 gnd.n803 292.5
R512 gnd.n808 gnd.n807 292.5
R513 gnd.n813 gnd.n812 292.5
R514 gnd.n814 gnd.n813 292.5
R515 gnd.n818 gnd.n817 292.5
R516 gnd.n819 gnd.n818 292.5
R517 gnd.n823 gnd.n822 292.5
R518 gnd.n824 gnd.n823 292.5
R519 gnd.n828 gnd.n827 292.5
R520 gnd.n829 gnd.n828 292.5
R521 gnd.n833 gnd.n832 292.5
R522 gnd.n834 gnd.n833 292.5
R523 gnd.n838 gnd.n837 292.5
R524 gnd.n839 gnd.n838 292.5
R525 gnd.n843 gnd.n842 292.5
R526 gnd.n844 gnd.n843 292.5
R527 gnd.n848 gnd.n847 292.5
R528 gnd.n849 gnd.n848 292.5
R529 gnd.n853 gnd.n852 292.5
R530 gnd.n858 gnd.n857 292.5
R531 gnd.n859 gnd.n858 292.5
R532 gnd.n863 gnd.n862 292.5
R533 gnd.n864 gnd.n863 292.5
R534 gnd.n868 gnd.n867 292.5
R535 gnd.n869 gnd.n868 292.5
R536 gnd.n873 gnd.n872 292.5
R537 gnd.n874 gnd.n873 292.5
R538 gnd.n878 gnd.n877 292.5
R539 gnd.n879 gnd.n878 292.5
R540 gnd.n883 gnd.n882 292.5
R541 gnd.n884 gnd.n883 292.5
R542 gnd.n888 gnd.n887 292.5
R543 gnd.n889 gnd.n888 292.5
R544 gnd.n893 gnd.n892 292.5
R545 gnd.n894 gnd.n893 292.5
R546 gnd.n898 gnd.n897 292.5
R547 gnd.n899 gnd.n898 292.5
R548 gnd.n903 gnd.n902 292.5
R549 gnd.n904 gnd.n903 292.5
R550 gnd.n908 gnd.n907 292.5
R551 gnd.n909 gnd.n908 292.5
R552 gnd.n913 gnd.n912 292.5
R553 gnd.n914 gnd.n913 292.5
R554 gnd.n918 gnd.n917 292.5
R555 gnd.n919 gnd.n918 292.5
R556 gnd.n923 gnd.n922 292.5
R557 gnd.n928 gnd.n927 292.5
R558 gnd.n929 gnd.n928 292.5
R559 gnd.n933 gnd.n932 292.5
R560 gnd.n938 gnd.n937 292.5
R561 gnd.n939 gnd.n938 292.5
R562 gnd.n618 gnd.n617 292.5
R563 gnd.n619 gnd.n618 292.5
R564 gnd.n944 gnd.n943 292.5
R565 gnd.n945 gnd.n944 292.5
R566 gnd.n950 gnd.n949 292.5
R567 gnd.n951 gnd.n950 292.5
R568 gnd.n957 gnd.n956 292.5
R569 gnd.n958 gnd.n957 292.5
R570 gnd.n964 gnd.n963 292.5
R571 gnd.n965 gnd.n964 292.5
R572 gnd.n971 gnd.n970 292.5
R573 gnd.n972 gnd.n971 292.5
R574 gnd.n978 gnd.n977 292.5
R575 gnd.n979 gnd.n978 292.5
R576 gnd.n985 gnd.n984 292.5
R577 gnd.n986 gnd.n985 292.5
R578 gnd.n992 gnd.n991 292.5
R579 gnd.n993 gnd.n992 292.5
R580 gnd.n1004 gnd.n1003 292.5
R581 gnd.n1005 gnd.n1004 292.5
R582 gnd.n999 gnd.n998 292.5
R583 gnd.n1000 gnd.n999 292.5
R584 gnd.n611 gnd.n610 292.5
R585 gnd.n612 gnd.n611 292.5
R586 gnd.n604 gnd.n603 292.5
R587 gnd.n605 gnd.n604 292.5
R588 gnd.n598 gnd.n597 292.5
R589 gnd.n592 gnd.n591 292.5
R590 gnd.n586 gnd.n585 292.5
R591 gnd.n580 gnd.n579 292.5
R592 gnd.n574 gnd.n573 292.5
R593 gnd.n569 gnd.n568 292.5
R594 gnd.n555 gnd.n554 292.5
R595 gnd.n942 gnd.n620 292.5
R596 gnd.n620 gnd.n619 292.5
R597 gnd.n941 gnd.n940 292.5
R598 gnd.n940 gnd.n939 292.5
R599 gnd.n935 gnd.n934 292.5
R600 gnd.n934 gnd.n933 292.5
R601 gnd.n931 gnd.n930 292.5
R602 gnd.n930 gnd.n929 292.5
R603 gnd.n925 gnd.n924 292.5
R604 gnd.n924 gnd.n923 292.5
R605 gnd.n921 gnd.n920 292.5
R606 gnd.n920 gnd.n919 292.5
R607 gnd.n916 gnd.n915 292.5
R608 gnd.n915 gnd.n914 292.5
R609 gnd.n911 gnd.n910 292.5
R610 gnd.n910 gnd.n909 292.5
R611 gnd.n906 gnd.n905 292.5
R612 gnd.n905 gnd.n904 292.5
R613 gnd.n901 gnd.n900 292.5
R614 gnd.n900 gnd.n899 292.5
R615 gnd.n896 gnd.n895 292.5
R616 gnd.n895 gnd.n894 292.5
R617 gnd.n891 gnd.n890 292.5
R618 gnd.n890 gnd.n889 292.5
R619 gnd.n886 gnd.n885 292.5
R620 gnd.n885 gnd.n884 292.5
R621 gnd.n881 gnd.n880 292.5
R622 gnd.n880 gnd.n879 292.5
R623 gnd.n876 gnd.n875 292.5
R624 gnd.n875 gnd.n874 292.5
R625 gnd.n871 gnd.n870 292.5
R626 gnd.n870 gnd.n869 292.5
R627 gnd.n866 gnd.n865 292.5
R628 gnd.n865 gnd.n864 292.5
R629 gnd.n861 gnd.n860 292.5
R630 gnd.n860 gnd.n859 292.5
R631 gnd.n855 gnd.n854 292.5
R632 gnd.n854 gnd.n853 292.5
R633 gnd.n851 gnd.n850 292.5
R634 gnd.n850 gnd.n849 292.5
R635 gnd.n846 gnd.n845 292.5
R636 gnd.n845 gnd.n844 292.5
R637 gnd.n841 gnd.n840 292.5
R638 gnd.n840 gnd.n839 292.5
R639 gnd.n836 gnd.n835 292.5
R640 gnd.n835 gnd.n834 292.5
R641 gnd.n831 gnd.n830 292.5
R642 gnd.n830 gnd.n829 292.5
R643 gnd.n826 gnd.n825 292.5
R644 gnd.n825 gnd.n824 292.5
R645 gnd.n821 gnd.n820 292.5
R646 gnd.n820 gnd.n819 292.5
R647 gnd.n816 gnd.n815 292.5
R648 gnd.n815 gnd.n814 292.5
R649 gnd.n810 gnd.n809 292.5
R650 gnd.n809 gnd.n808 292.5
R651 gnd.n806 gnd.n805 292.5
R652 gnd.n805 gnd.n804 292.5
R653 gnd.n799 gnd.n798 292.5
R654 gnd.n798 gnd.n797 292.5
R655 gnd.n795 gnd.n794 292.5
R656 gnd.n794 gnd.n793 292.5
R657 gnd.n791 gnd.n790 292.5
R658 gnd.n790 gnd.n789 292.5
R659 gnd.n785 gnd.n784 292.5
R660 gnd.n784 gnd.n783 292.5
R661 gnd.n781 gnd.n780 292.5
R662 gnd.n780 gnd.n779 292.5
R663 gnd.n776 gnd.n775 292.5
R664 gnd.n775 gnd.n774 292.5
R665 gnd.n771 gnd.n770 292.5
R666 gnd.n770 gnd.n769 292.5
R667 gnd.n766 gnd.n765 292.5
R668 gnd.n765 gnd.n764 292.5
R669 gnd.n760 gnd.n759 292.5
R670 gnd.n759 gnd.n758 292.5
R671 gnd.n756 gnd.n755 292.5
R672 gnd.n755 gnd.n754 292.5
R673 gnd.n751 gnd.n750 292.5
R674 gnd.n750 gnd.n749 292.5
R675 gnd.n743 gnd.n742 292.5
R676 gnd.n742 gnd.n741 292.5
R677 gnd.n739 gnd.n738 292.5
R678 gnd.n738 gnd.n737 292.5
R679 gnd.n735 gnd.n734 292.5
R680 gnd.n734 gnd.n733 292.5
R681 gnd.n731 gnd.n730 292.5
R682 gnd.n730 gnd.n729 292.5
R683 gnd.n726 gnd.n725 292.5
R684 gnd.n725 gnd.n724 292.5
R685 gnd.n721 gnd.n720 292.5
R686 gnd.n720 gnd.n719 292.5
R687 gnd.n716 gnd.n715 292.5
R688 gnd.n715 gnd.n714 292.5
R689 gnd.n711 gnd.n710 292.5
R690 gnd.n710 gnd.n709 292.5
R691 gnd.n706 gnd.n705 292.5
R692 gnd.n705 gnd.n704 292.5
R693 gnd.n701 gnd.n700 292.5
R694 gnd.n700 gnd.n699 292.5
R695 gnd.n696 gnd.n695 292.5
R696 gnd.n695 gnd.n694 292.5
R697 gnd.n691 gnd.n690 292.5
R698 gnd.n690 gnd.n689 292.5
R699 gnd.n685 gnd.n684 292.5
R700 gnd.n684 gnd.n683 292.5
R701 gnd.n681 gnd.n680 292.5
R702 gnd.n680 gnd.n679 292.5
R703 gnd.n675 gnd.n674 292.5
R704 gnd.n674 gnd.n673 292.5
R705 gnd.n671 gnd.n670 292.5
R706 gnd.n670 gnd.n669 292.5
R707 gnd.n666 gnd.n665 292.5
R708 gnd.n665 gnd.n664 292.5
R709 gnd.n659 gnd.n658 292.5
R710 gnd.n658 gnd.n657 292.5
R711 gnd.n655 gnd.n654 292.5
R712 gnd.n654 gnd.n653 292.5
R713 gnd.n651 gnd.n650 292.5
R714 gnd.n650 gnd.n649 292.5
R715 gnd.n646 gnd.n645 292.5
R716 gnd.n645 gnd.n644 292.5
R717 gnd.n642 gnd.n641 292.5
R718 gnd.n641 gnd.n640 292.5
R719 gnd.n638 gnd.n637 292.5
R720 gnd.n637 gnd.n636 292.5
R721 gnd.n634 gnd.n633 292.5
R722 gnd.n633 gnd.n632 292.5
R723 gnd.n629 gnd.n628 292.5
R724 gnd.n557 gnd.n556 292.5
R725 gnd.n556 gnd.n555 292.5
R726 gnd.n571 gnd.n570 292.5
R727 gnd.n570 gnd.n569 292.5
R728 gnd.n576 gnd.n575 292.5
R729 gnd.n575 gnd.n574 292.5
R730 gnd.n582 gnd.n581 292.5
R731 gnd.n581 gnd.n580 292.5
R732 gnd.n588 gnd.n587 292.5
R733 gnd.n587 gnd.n586 292.5
R734 gnd.n594 gnd.n593 292.5
R735 gnd.n593 gnd.n592 292.5
R736 gnd.n600 gnd.n599 292.5
R737 gnd.n599 gnd.n598 292.5
R738 gnd.n607 gnd.n606 292.5
R739 gnd.n606 gnd.n605 292.5
R740 gnd.n614 gnd.n613 292.5
R741 gnd.n613 gnd.n612 292.5
R742 gnd.n1002 gnd.n1001 292.5
R743 gnd.n1001 gnd.n1000 292.5
R744 gnd.n1007 gnd.n1006 292.5
R745 gnd.n1006 gnd.n1005 292.5
R746 gnd.n995 gnd.n994 292.5
R747 gnd.n994 gnd.n993 292.5
R748 gnd.n988 gnd.n987 292.5
R749 gnd.n987 gnd.n986 292.5
R750 gnd.n981 gnd.n980 292.5
R751 gnd.n980 gnd.n979 292.5
R752 gnd.n974 gnd.n973 292.5
R753 gnd.n973 gnd.n972 292.5
R754 gnd.n967 gnd.n966 292.5
R755 gnd.n966 gnd.n965 292.5
R756 gnd.n960 gnd.n959 292.5
R757 gnd.n959 gnd.n958 292.5
R758 gnd.n953 gnd.n952 292.5
R759 gnd.n952 gnd.n951 292.5
R760 gnd.n947 gnd.n946 292.5
R761 gnd.n946 gnd.n945 292.5
R762 gnd.n592 gnd.t112 263.38
R763 gnd.n894 gnd.t45 263.38
R764 gnd.n774 gnd.t59 263.38
R765 gnd.n653 gnd.t107 263.38
R766 gnd.n286 gnd.n285 255.63
R767 gnd.n7 gnd.n6 255.63
R768 gnd.n566 gnd.n565 253.487
R769 gnd.n12 gnd.t33 247.887
R770 gnd.n130 gnd.t110 247.887
R771 gnd.n409 gnd.t97 247.887
R772 gnd.n291 gnd.t93 247.887
R773 gnd.n979 gnd.t62 232.394
R774 gnd.n929 gnd.t103 232.394
R775 gnd.n853 gnd.t55 232.394
R776 gnd.n808 gnd.t48 232.394
R777 gnd.n733 gnd.t82 232.394
R778 gnd.n689 gnd.t56 232.394
R779 gnd.n60 gnd.t116 216.901
R780 gnd.n75 gnd.t19 216.901
R781 gnd.n354 gnd.t85 216.901
R782 gnd.n339 gnd.t118 216.901
R783 gnd.n965 gnd.t72 201.408
R784 gnd.n939 gnd.t53 201.408
R785 gnd.n844 gnd.t73 201.408
R786 gnd.n819 gnd.t2 201.408
R787 gnd.n724 gnd.t69 201.408
R788 gnd.n699 gnd.t109 201.408
R789 gnd.n26 gnd.t9 185.915
R790 gnd.n114 gnd.t100 185.915
R791 gnd.n393 gnd.t80 185.915
R792 gnd.n309 gnd.t11 185.915
R793 gnd.n580 gnd.t64 170.422
R794 gnd.n612 gnd.t60 170.422
R795 gnd.n904 gnd.t106 170.422
R796 gnd.n879 gnd.t38 170.422
R797 gnd.n783 gnd.t3 170.422
R798 gnd.n758 gnd.t1 170.422
R799 gnd.n664 gnd.t49 170.422
R800 gnd.n640 gnd.t40 170.422
R801 gnd.n154 gnd.t13 154.929
R802 gnd.n433 gnd.t21 154.929
R803 gnd.n569 gnd.t41 139.436
R804 gnd.n1005 gnd.t30 139.436
R805 gnd.n914 gnd.t43 139.436
R806 gnd.n869 gnd.t70 139.436
R807 gnd.n793 gnd.t29 139.436
R808 gnd.n749 gnd.t58 139.436
R809 gnd.n673 gnd.t115 139.436
R810 gnd.n632 gnd.t54 139.436
R811 gnd.n37 gnd.t83 123.943
R812 gnd.n98 gnd.t91 123.943
R813 gnd.n377 gnd.t113 123.943
R814 gnd.n316 gnd.t35 123.943
R815 gnd.n284 gnd.n283 118.219
R816 gnd.n625 gnd.n624 118.219
R817 gnd.n5 gnd.n4 118.219
R818 gnd.n564 gnd.n563 118.219
R819 gnd.n634 gnd.n630 118.219
R820 gnd.n630 gnd.n629 114.718
R821 gnd.n951 gnd.t4 108.45
R822 gnd.n945 gnd.t61 108.45
R823 gnd.n834 gnd.t66 108.45
R824 gnd.n829 gnd.t52 108.45
R825 gnd.n714 gnd.t46 108.45
R826 gnd.n709 gnd.t37 108.45
R827 gnd.n44 gnd.t76 92.957
R828 gnd.n91 gnd.t87 92.957
R829 gnd.n370 gnd.t17 92.957
R830 gnd.n323 gnd.t7 92.957
R831 gnd.n555 gnd.t28 77.464
R832 gnd.n993 gnd.t16 77.464
R833 gnd.n919 gnd.t57 77.464
R834 gnd.n864 gnd.t63 77.464
R835 gnd.n797 gnd.t51 77.464
R836 gnd.n741 gnd.t65 77.464
R837 gnd.n679 gnd.t104 77.464
R838 gnd.n628 gnd.t0 77.464
R839 gnd.n146 gnd.t78 61.971
R840 gnd.n425 gnd.t74 61.971
R841 gnd.n586 gnd.t23 46.478
R842 gnd.n605 gnd.t67 46.478
R843 gnd.n899 gnd.t71 46.478
R844 gnd.n884 gnd.t68 46.478
R845 gnd.n779 gnd.t47 46.478
R846 gnd.n764 gnd.t105 46.478
R847 gnd.n657 gnd.t44 46.478
R848 gnd.n644 gnd.t108 46.478
R849 gnd.n19 gnd.t31 30.985
R850 gnd.n122 gnd.t95 30.985
R851 gnd.n401 gnd.t5 30.985
R852 gnd.n298 gnd.t89 30.985
R853 gnd.n227 gnd.t34 28.876
R854 gnd.n501 gnd.t94 28.876
R855 gnd.n4 gnd.n3 25.6
R856 gnd.n3 gnd.n2 25.6
R857 gnd.n2 gnd.n1 25.6
R858 gnd.n1 gnd.n0 25.6
R859 gnd.n280 gnd.n279 25.6
R860 gnd.n281 gnd.n280 25.6
R861 gnd.n282 gnd.n281 25.6
R862 gnd.n283 gnd.n282 25.6
R863 gnd.n563 gnd.n562 25.6
R864 gnd.n562 gnd.n561 25.6
R865 gnd.n561 gnd.n560 25.6
R866 gnd.n560 gnd.n559 25.6
R867 gnd.n559 gnd.n558 25.6
R868 gnd.n937 gnd.n936 25.6
R869 gnd.n927 gnd.n926 25.6
R870 gnd.n857 gnd.n856 25.6
R871 gnd.n812 gnd.n811 25.6
R872 gnd.n802 gnd.n801 25.6
R873 gnd.n801 gnd.n800 25.6
R874 gnd.n787 gnd.n786 25.6
R875 gnd.n762 gnd.n761 25.6
R876 gnd.n747 gnd.n746 25.6
R877 gnd.n746 gnd.n745 25.6
R878 gnd.n745 gnd.n744 25.6
R879 gnd.n687 gnd.n686 25.6
R880 gnd.n677 gnd.n676 25.6
R881 gnd.n662 gnd.n661 25.6
R882 gnd.n661 gnd.n660 25.6
R883 gnd.n622 gnd.n621 25.6
R884 gnd.n623 gnd.n622 25.6
R885 gnd.n624 gnd.n623 25.6
R886 gnd.n942 gnd.n941 25.6
R887 gnd.n941 gnd.n935 25.6
R888 gnd.n935 gnd.n931 25.6
R889 gnd.n931 gnd.n925 25.6
R890 gnd.n925 gnd.n921 25.6
R891 gnd.n921 gnd.n916 25.6
R892 gnd.n916 gnd.n911 25.6
R893 gnd.n911 gnd.n906 25.6
R894 gnd.n906 gnd.n901 25.6
R895 gnd.n901 gnd.n896 25.6
R896 gnd.n896 gnd.n891 25.6
R897 gnd.n891 gnd.n886 25.6
R898 gnd.n886 gnd.n881 25.6
R899 gnd.n881 gnd.n876 25.6
R900 gnd.n876 gnd.n871 25.6
R901 gnd.n871 gnd.n866 25.6
R902 gnd.n866 gnd.n861 25.6
R903 gnd.n861 gnd.n855 25.6
R904 gnd.n855 gnd.n851 25.6
R905 gnd.n851 gnd.n846 25.6
R906 gnd.n846 gnd.n841 25.6
R907 gnd.n841 gnd.n836 25.6
R908 gnd.n836 gnd.n831 25.6
R909 gnd.n831 gnd.n826 25.6
R910 gnd.n826 gnd.n821 25.6
R911 gnd.n821 gnd.n816 25.6
R912 gnd.n816 gnd.n810 25.6
R913 gnd.n810 gnd.n806 25.6
R914 gnd.n806 gnd.n799 25.6
R915 gnd.n799 gnd.n795 25.6
R916 gnd.n795 gnd.n791 25.6
R917 gnd.n791 gnd.n785 25.6
R918 gnd.n785 gnd.n781 25.6
R919 gnd.n781 gnd.n776 25.6
R920 gnd.n776 gnd.n771 25.6
R921 gnd.n771 gnd.n766 25.6
R922 gnd.n766 gnd.n760 25.6
R923 gnd.n760 gnd.n756 25.6
R924 gnd.n756 gnd.n751 25.6
R925 gnd.n751 gnd.n743 25.6
R926 gnd.n743 gnd.n739 25.6
R927 gnd.n739 gnd.n735 25.6
R928 gnd.n735 gnd.n731 25.6
R929 gnd.n731 gnd.n726 25.6
R930 gnd.n726 gnd.n721 25.6
R931 gnd.n721 gnd.n716 25.6
R932 gnd.n716 gnd.n711 25.6
R933 gnd.n711 gnd.n706 25.6
R934 gnd.n706 gnd.n701 25.6
R935 gnd.n701 gnd.n696 25.6
R936 gnd.n696 gnd.n691 25.6
R937 gnd.n691 gnd.n685 25.6
R938 gnd.n685 gnd.n681 25.6
R939 gnd.n681 gnd.n675 25.6
R940 gnd.n675 gnd.n671 25.6
R941 gnd.n671 gnd.n666 25.6
R942 gnd.n666 gnd.n659 25.6
R943 gnd.n659 gnd.n655 25.6
R944 gnd.n655 gnd.n651 25.6
R945 gnd.n651 gnd.n646 25.6
R946 gnd.n646 gnd.n642 25.6
R947 gnd.n642 gnd.n638 25.6
R948 gnd.n638 gnd.n634 25.6
R949 gnd.n474 gnd.t25 23.571
R950 gnd.n474 gnd.t119 23.571
R951 gnd.n447 gnd.t98 23.571
R952 gnd.n447 gnd.t6 23.571
R953 gnd.n173 gnd.t96 23.571
R954 gnd.n173 gnd.t111 23.571
R955 gnd.n200 gnd.t117 23.571
R956 gnd.n200 gnd.t27 23.571
R957 gnd.n218 gnd.t32 23.571
R958 gnd.n218 gnd.t10 23.571
R959 gnd.n209 gnd.t84 23.571
R960 gnd.n209 gnd.t77 23.571
R961 gnd.n191 gnd.t20 23.571
R962 gnd.n191 gnd.t88 23.571
R963 gnd.n182 gnd.t92 23.571
R964 gnd.n182 gnd.t101 23.571
R965 gnd.n164 gnd.t79 23.571
R966 gnd.n164 gnd.t14 23.571
R967 gnd.n438 gnd.t22 23.571
R968 gnd.n438 gnd.t75 23.571
R969 gnd.n456 gnd.t81 23.571
R970 gnd.n456 gnd.t114 23.571
R971 gnd.n465 gnd.t18 23.571
R972 gnd.n465 gnd.t86 23.571
R973 gnd.n483 gnd.t8 23.571
R974 gnd.n483 gnd.t36 23.571
R975 gnd.n492 gnd.t12 23.571
R976 gnd.n492 gnd.t90 23.571
R977 gnd.n947 gnd.n942 18.394
R978 gnd.n972 gnd.t50 15.492
R979 gnd.n933 gnd.t99 15.492
R980 gnd.n849 gnd.t102 15.492
R981 gnd.n814 gnd.t15 15.492
R982 gnd.n729 gnd.t39 15.492
R983 gnd.n694 gnd.t42 15.492
R984 gnd.n232 gnd.n227 14.007
R985 gnd.n506 gnd.n501 14.007
R986 gnd.n480 gnd.n475 8.032
R987 gnd.n453 gnd.n448 8.032
R988 gnd.n179 gnd.n174 8.032
R989 gnd.n206 gnd.n201 8.032
R990 gnd.n224 gnd.n219 8.032
R991 gnd.n215 gnd.n210 8.032
R992 gnd.n197 gnd.n192 8.032
R993 gnd.n188 gnd.n183 8.032
R994 gnd.n170 gnd.n165 8.032
R995 gnd.n444 gnd.n439 8.032
R996 gnd.n462 gnd.n457 8.032
R997 gnd.n471 gnd.n466 8.032
R998 gnd.n489 gnd.n484 8.032
R999 gnd.n498 gnd.n493 8.032
R1000 gnd.n955 gnd.n948 4.658
R1001 gnd.n572 gnd.n571 4.65
R1002 gnd.n578 gnd.n577 4.65
R1003 gnd.n584 gnd.n583 4.65
R1004 gnd.n590 gnd.n589 4.65
R1005 gnd.n596 gnd.n595 4.65
R1006 gnd.n602 gnd.n601 4.65
R1007 gnd.n609 gnd.n608 4.65
R1008 gnd.n616 gnd.n615 4.65
R1009 gnd.n1009 gnd.n1008 4.65
R1010 gnd.n997 gnd.n996 4.65
R1011 gnd.n990 gnd.n989 4.65
R1012 gnd.n983 gnd.n982 4.65
R1013 gnd.n976 gnd.n975 4.65
R1014 gnd.n969 gnd.n968 4.65
R1015 gnd.n962 gnd.n961 4.65
R1016 gnd.n955 gnd.n954 4.65
R1017 gnd.n1008 gnd.n1007 4.608
R1018 gnd.n1008 gnd.n1002 4.096
R1019 gnd.n996 gnd.n995 4.096
R1020 gnd.n477 gnd.n476 3.85
R1021 gnd.n450 gnd.n449 3.85
R1022 gnd.n176 gnd.n175 3.85
R1023 gnd.n203 gnd.n202 3.85
R1024 gnd.n229 gnd.n228 3.85
R1025 gnd.n221 gnd.n220 3.85
R1026 gnd.n212 gnd.n211 3.85
R1027 gnd.n194 gnd.n193 3.85
R1028 gnd.n185 gnd.n184 3.85
R1029 gnd.n167 gnd.n166 3.85
R1030 gnd.n441 gnd.n440 3.85
R1031 gnd.n459 gnd.n458 3.85
R1032 gnd.n468 gnd.n467 3.85
R1033 gnd.n486 gnd.n485 3.85
R1034 gnd.n495 gnd.n494 3.85
R1035 gnd.n503 gnd.n502 3.85
R1036 gnd.n615 gnd.n614 3.584
R1037 gnd.n989 gnd.n988 3.584
R1038 gnd.n33 gnd.n28 3.572
R1039 gnd.n162 gnd.n161 3.572
R1040 gnd.n312 gnd.n311 3.572
R1041 gnd.n22 gnd.n21 3.175
R1042 gnd.n33 gnd.n32 3.175
R1043 gnd.n162 gnd.n156 3.175
R1044 gnd.n436 gnd.n435 3.175
R1045 gnd.n312 gnd.n307 3.175
R1046 gnd.n301 gnd.n300 3.175
R1047 gnd.n608 gnd.n607 3.072
R1048 gnd.n982 gnd.n981 3.072
R1049 gnd.n9 gnd.n8 3.033
R1050 gnd.n16 gnd.n15 3.033
R1051 gnd.n23 gnd.n22 3.033
R1052 gnd.n34 gnd.n33 3.033
R1053 gnd.n41 gnd.n40 3.033
R1054 gnd.n48 gnd.n47 3.033
R1055 gnd.n56 gnd.n55 3.033
R1056 gnd.n64 gnd.n63 3.033
R1057 gnd.n71 gnd.n70 3.033
R1058 gnd.n79 gnd.n78 3.033
R1059 gnd.n87 gnd.n86 3.033
R1060 gnd.n94 gnd.n93 3.033
R1061 gnd.n102 gnd.n101 3.033
R1062 gnd.n110 gnd.n109 3.033
R1063 gnd.n118 gnd.n117 3.033
R1064 gnd.n126 gnd.n125 3.033
R1065 gnd.n134 gnd.n133 3.033
R1066 gnd.n142 gnd.n141 3.033
R1067 gnd.n150 gnd.n149 3.033
R1068 gnd.n163 gnd.n162 3.033
R1069 gnd.n437 gnd.n436 3.033
R1070 gnd.n429 gnd.n428 3.033
R1071 gnd.n421 gnd.n420 3.033
R1072 gnd.n413 gnd.n412 3.033
R1073 gnd.n405 gnd.n404 3.033
R1074 gnd.n397 gnd.n396 3.033
R1075 gnd.n389 gnd.n388 3.033
R1076 gnd.n381 gnd.n380 3.033
R1077 gnd.n373 gnd.n372 3.033
R1078 gnd.n366 gnd.n365 3.033
R1079 gnd.n358 gnd.n357 3.033
R1080 gnd.n350 gnd.n349 3.033
R1081 gnd.n343 gnd.n342 3.033
R1082 gnd.n335 gnd.n334 3.033
R1083 gnd.n327 gnd.n326 3.033
R1084 gnd.n320 gnd.n319 3.033
R1085 gnd.n313 gnd.n312 3.033
R1086 gnd.n302 gnd.n301 3.033
R1087 gnd.n295 gnd.n294 3.033
R1088 gnd.n288 gnd.n287 3.033
R1089 gnd.n15 gnd.n14 2.778
R1090 gnd.n40 gnd.n39 2.778
R1091 gnd.n149 gnd.n148 2.778
R1092 gnd.n428 gnd.n427 2.778
R1093 gnd.n319 gnd.n318 2.778
R1094 gnd.n294 gnd.n293 2.778
R1095 gnd.n567 gnd.n557 2.569
R1096 gnd.n601 gnd.n600 2.56
R1097 gnd.n975 gnd.n974 2.56
R1098 gnd.n47 gnd.n46 2.381
R1099 gnd.n141 gnd.n140 2.381
R1100 gnd.n420 gnd.n419 2.381
R1101 gnd.n326 gnd.n325 2.381
R1102 gnd.n595 gnd.n594 2.048
R1103 gnd.n968 gnd.n967 2.048
R1104 gnd.n55 gnd.n54 1.984
R1105 gnd.n133 gnd.n132 1.984
R1106 gnd.n412 gnd.n411 1.984
R1107 gnd.n334 gnd.n333 1.984
R1108 gnd.n475 gnd.n474 1.601
R1109 gnd.n448 gnd.n447 1.601
R1110 gnd.n174 gnd.n173 1.601
R1111 gnd.n201 gnd.n200 1.601
R1112 gnd.n219 gnd.n218 1.601
R1113 gnd.n210 gnd.n209 1.601
R1114 gnd.n192 gnd.n191 1.601
R1115 gnd.n183 gnd.n182 1.601
R1116 gnd.n165 gnd.n164 1.601
R1117 gnd.n439 gnd.n438 1.601
R1118 gnd.n457 gnd.n456 1.601
R1119 gnd.n466 gnd.n465 1.601
R1120 gnd.n484 gnd.n483 1.601
R1121 gnd.n493 gnd.n492 1.601
R1122 gnd.n63 gnd.n62 1.587
R1123 gnd.n125 gnd.n124 1.587
R1124 gnd.n404 gnd.n403 1.587
R1125 gnd.n342 gnd.n341 1.587
R1126 gnd.n589 gnd.n588 1.536
R1127 gnd.n961 gnd.n960 1.536
R1128 gnd.n572 gnd.n567 1.435
R1129 gnd.n70 gnd.n69 1.19
R1130 gnd.n117 gnd.n116 1.19
R1131 gnd.n396 gnd.n395 1.19
R1132 gnd.n349 gnd.n348 1.19
R1133 gnd.n583 gnd.n582 1.024
R1134 gnd.n954 gnd.n953 1.024
R1135 gnd.n1011 gnd.n1010 0.911
R1136 gnd.n78 gnd.n77 0.793
R1137 gnd.n109 gnd.n108 0.793
R1138 gnd.n388 gnd.n387 0.793
R1139 gnd.n357 gnd.n356 0.793
R1140 gnd.n481 gnd.n480 0.617
R1141 gnd.n454 gnd.n453 0.617
R1142 gnd.n180 gnd.n179 0.617
R1143 gnd.n207 gnd.n206 0.617
R1144 gnd.n233 gnd.n232 0.617
R1145 gnd.n225 gnd.n224 0.617
R1146 gnd.n216 gnd.n215 0.617
R1147 gnd.n198 gnd.n197 0.617
R1148 gnd.n189 gnd.n188 0.617
R1149 gnd.n171 gnd.n170 0.617
R1150 gnd.n445 gnd.n444 0.617
R1151 gnd.n463 gnd.n462 0.617
R1152 gnd.n472 gnd.n471 0.617
R1153 gnd.n490 gnd.n489 0.617
R1154 gnd.n499 gnd.n498 0.617
R1155 gnd.n507 gnd.n506 0.617
R1156 gnd.n577 gnd.n576 0.512
R1157 gnd.n948 gnd.n947 0.512
R1158 gnd.n509 gnd.n508 0.454
R1159 gnd.n235 gnd.n234 0.454
R1160 gnd.n526 gnd.n482 0.443
R1161 gnd.n544 gnd.n455 0.443
R1162 gnd.n270 gnd.n181 0.443
R1163 gnd.n252 gnd.n208 0.443
R1164 gnd.n240 gnd.n226 0.443
R1165 gnd.n246 gnd.n217 0.443
R1166 gnd.n258 gnd.n199 0.443
R1167 gnd.n264 gnd.n190 0.443
R1168 gnd.n276 gnd.n172 0.443
R1169 gnd.n550 gnd.n446 0.443
R1170 gnd.n538 gnd.n464 0.443
R1171 gnd.n532 gnd.n473 0.443
R1172 gnd.n520 gnd.n491 0.443
R1173 gnd.n514 gnd.n500 0.443
R1174 gnd.n86 gnd.n85 0.396
R1175 gnd.n101 gnd.n100 0.396
R1176 gnd.n380 gnd.n379 0.396
R1177 gnd.n365 gnd.n364 0.396
R1178 gnd.n480 gnd.n479 0.098
R1179 gnd.n453 gnd.n452 0.098
R1180 gnd.n179 gnd.n178 0.098
R1181 gnd.n206 gnd.n205 0.098
R1182 gnd.n232 gnd.n231 0.098
R1183 gnd.n224 gnd.n223 0.098
R1184 gnd.n215 gnd.n214 0.098
R1185 gnd.n197 gnd.n196 0.098
R1186 gnd.n188 gnd.n187 0.098
R1187 gnd.n170 gnd.n169 0.098
R1188 gnd.n444 gnd.n443 0.098
R1189 gnd.n462 gnd.n461 0.098
R1190 gnd.n471 gnd.n470 0.098
R1191 gnd.n489 gnd.n488 0.098
R1192 gnd.n498 gnd.n497 0.098
R1193 gnd.n506 gnd.n505 0.098
R1194 gnd.n278 gnd.n277 0.044
R1195 gnd.n552 gnd.n551 0.044
R1196 gnd.n482 gnd.n481 0.039
R1197 gnd.n455 gnd.n454 0.039
R1198 gnd.n181 gnd.n180 0.039
R1199 gnd.n208 gnd.n207 0.039
R1200 gnd.n234 gnd.n233 0.039
R1201 gnd.n226 gnd.n225 0.039
R1202 gnd.n217 gnd.n216 0.039
R1203 gnd.n199 gnd.n198 0.039
R1204 gnd.n190 gnd.n189 0.039
R1205 gnd.n172 gnd.n171 0.039
R1206 gnd.n446 gnd.n445 0.039
R1207 gnd.n464 gnd.n463 0.039
R1208 gnd.n473 gnd.n472 0.039
R1209 gnd.n491 gnd.n490 0.039
R1210 gnd.n500 gnd.n499 0.039
R1211 gnd.n508 gnd.n507 0.039
R1212 gnd.n236 gnd.n235 0.033
R1213 gnd.n510 gnd.n509 0.033
R1214 gnd.n237 gnd.n236 0.022
R1215 gnd.n238 gnd.n237 0.022
R1216 gnd.n239 gnd.n238 0.022
R1217 gnd.n242 gnd.n241 0.022
R1218 gnd.n243 gnd.n242 0.022
R1219 gnd.n244 gnd.n243 0.022
R1220 gnd.n245 gnd.n244 0.022
R1221 gnd.n248 gnd.n247 0.022
R1222 gnd.n249 gnd.n248 0.022
R1223 gnd.n250 gnd.n249 0.022
R1224 gnd.n251 gnd.n250 0.022
R1225 gnd.n252 gnd.n251 0.022
R1226 gnd.n253 gnd.n252 0.022
R1227 gnd.n254 gnd.n253 0.022
R1228 gnd.n255 gnd.n254 0.022
R1229 gnd.n256 gnd.n255 0.022
R1230 gnd.n257 gnd.n256 0.022
R1231 gnd.n260 gnd.n259 0.022
R1232 gnd.n261 gnd.n260 0.022
R1233 gnd.n262 gnd.n261 0.022
R1234 gnd.n263 gnd.n262 0.022
R1235 gnd.n266 gnd.n265 0.022
R1236 gnd.n267 gnd.n266 0.022
R1237 gnd.n268 gnd.n267 0.022
R1238 gnd.n269 gnd.n268 0.022
R1239 gnd.n270 gnd.n269 0.022
R1240 gnd.n271 gnd.n270 0.022
R1241 gnd.n272 gnd.n271 0.022
R1242 gnd.n273 gnd.n272 0.022
R1243 gnd.n274 gnd.n273 0.022
R1244 gnd.n275 gnd.n274 0.022
R1245 gnd.n549 gnd.n548 0.022
R1246 gnd.n548 gnd.n547 0.022
R1247 gnd.n547 gnd.n546 0.022
R1248 gnd.n546 gnd.n545 0.022
R1249 gnd.n545 gnd.n544 0.022
R1250 gnd.n544 gnd.n543 0.022
R1251 gnd.n543 gnd.n542 0.022
R1252 gnd.n542 gnd.n541 0.022
R1253 gnd.n541 gnd.n540 0.022
R1254 gnd.n540 gnd.n539 0.022
R1255 gnd.n537 gnd.n536 0.022
R1256 gnd.n536 gnd.n535 0.022
R1257 gnd.n535 gnd.n534 0.022
R1258 gnd.n534 gnd.n533 0.022
R1259 gnd.n531 gnd.n530 0.022
R1260 gnd.n530 gnd.n529 0.022
R1261 gnd.n529 gnd.n528 0.022
R1262 gnd.n528 gnd.n527 0.022
R1263 gnd.n527 gnd.n526 0.022
R1264 gnd.n526 gnd.n525 0.022
R1265 gnd.n525 gnd.n524 0.022
R1266 gnd.n524 gnd.n523 0.022
R1267 gnd.n523 gnd.n522 0.022
R1268 gnd.n522 gnd.n521 0.022
R1269 gnd.n519 gnd.n518 0.022
R1270 gnd.n518 gnd.n517 0.022
R1271 gnd.n517 gnd.n516 0.022
R1272 gnd.n516 gnd.n515 0.022
R1273 gnd.n513 gnd.n512 0.022
R1274 gnd.n512 gnd.n511 0.022
R1275 gnd.n511 gnd.n510 0.022
R1276 gnd.n241 gnd.n240 0.015
R1277 gnd.n246 gnd.n245 0.015
R1278 gnd.n259 gnd.n258 0.015
R1279 gnd.n264 gnd.n263 0.015
R1280 gnd.n277 gnd.n276 0.015
R1281 gnd.n551 gnd.n550 0.015
R1282 gnd.n538 gnd.n537 0.015
R1283 gnd.n533 gnd.n532 0.015
R1284 gnd.n520 gnd.n519 0.015
R1285 gnd.n515 gnd.n514 0.015
R1286 gnd.n578 gnd.n572 0.008
R1287 gnd.n584 gnd.n578 0.008
R1288 gnd.n590 gnd.n584 0.008
R1289 gnd.n596 gnd.n590 0.008
R1290 gnd.n602 gnd.n596 0.008
R1291 gnd.n609 gnd.n602 0.008
R1292 gnd.n616 gnd.n609 0.008
R1293 gnd.n1009 gnd.n997 0.008
R1294 gnd.n997 gnd.n990 0.008
R1295 gnd.n990 gnd.n983 0.008
R1296 gnd.n983 gnd.n976 0.008
R1297 gnd.n976 gnd.n969 0.008
R1298 gnd.n969 gnd.n962 0.008
R1299 gnd.n962 gnd.n955 0.008
R1300 gnd.n478 gnd.n477 0.008
R1301 gnd.n451 gnd.n450 0.008
R1302 gnd.n177 gnd.n176 0.008
R1303 gnd.n204 gnd.n203 0.008
R1304 gnd.n230 gnd.n229 0.008
R1305 gnd.n222 gnd.n221 0.008
R1306 gnd.n213 gnd.n212 0.008
R1307 gnd.n195 gnd.n194 0.008
R1308 gnd.n186 gnd.n185 0.008
R1309 gnd.n168 gnd.n167 0.008
R1310 gnd.n442 gnd.n441 0.008
R1311 gnd.n460 gnd.n459 0.008
R1312 gnd.n469 gnd.n468 0.008
R1313 gnd.n487 gnd.n486 0.008
R1314 gnd.n496 gnd.n495 0.008
R1315 gnd.n504 gnd.n503 0.008
R1316 gnd.n240 gnd.n239 0.007
R1317 gnd.n247 gnd.n246 0.007
R1318 gnd.n258 gnd.n257 0.007
R1319 gnd.n265 gnd.n264 0.007
R1320 gnd.n276 gnd.n275 0.007
R1321 gnd.n550 gnd.n549 0.007
R1322 gnd.n539 gnd.n538 0.007
R1323 gnd.n532 gnd.n531 0.007
R1324 gnd.n521 gnd.n520 0.007
R1325 gnd.n514 gnd.n513 0.007
R1326 gnd gnd.n1011 0.006
R1327 gnd.n278 gnd.n163 0.005
R1328 gnd.n552 gnd.n437 0.005
R1329 gnd.n10 gnd.n9 0.005
R1330 gnd.n16 gnd.n10 0.005
R1331 gnd.n17 gnd.n16 0.005
R1332 gnd.n23 gnd.n17 0.005
R1333 gnd.n24 gnd.n23 0.005
R1334 gnd.n34 gnd.n24 0.005
R1335 gnd.n35 gnd.n34 0.005
R1336 gnd.n41 gnd.n35 0.005
R1337 gnd.n42 gnd.n41 0.005
R1338 gnd.n48 gnd.n42 0.005
R1339 gnd.n49 gnd.n48 0.005
R1340 gnd.n56 gnd.n49 0.005
R1341 gnd.n57 gnd.n56 0.005
R1342 gnd.n64 gnd.n57 0.005
R1343 gnd.n65 gnd.n64 0.005
R1344 gnd.n71 gnd.n65 0.005
R1345 gnd.n72 gnd.n71 0.005
R1346 gnd.n79 gnd.n72 0.005
R1347 gnd.n80 gnd.n79 0.005
R1348 gnd.n87 gnd.n80 0.005
R1349 gnd.n88 gnd.n87 0.005
R1350 gnd.n94 gnd.n88 0.005
R1351 gnd.n95 gnd.n94 0.005
R1352 gnd.n102 gnd.n95 0.005
R1353 gnd.n103 gnd.n102 0.005
R1354 gnd.n110 gnd.n103 0.005
R1355 gnd.n111 gnd.n110 0.005
R1356 gnd.n118 gnd.n111 0.005
R1357 gnd.n119 gnd.n118 0.005
R1358 gnd.n126 gnd.n119 0.005
R1359 gnd.n127 gnd.n126 0.005
R1360 gnd.n134 gnd.n127 0.005
R1361 gnd.n135 gnd.n134 0.005
R1362 gnd.n142 gnd.n135 0.005
R1363 gnd.n143 gnd.n142 0.005
R1364 gnd.n150 gnd.n143 0.005
R1365 gnd.n151 gnd.n150 0.005
R1366 gnd.n163 gnd.n151 0.005
R1367 gnd.n437 gnd.n430 0.005
R1368 gnd.n430 gnd.n429 0.005
R1369 gnd.n429 gnd.n422 0.005
R1370 gnd.n422 gnd.n421 0.005
R1371 gnd.n421 gnd.n414 0.005
R1372 gnd.n414 gnd.n413 0.005
R1373 gnd.n413 gnd.n406 0.005
R1374 gnd.n406 gnd.n405 0.005
R1375 gnd.n405 gnd.n398 0.005
R1376 gnd.n398 gnd.n397 0.005
R1377 gnd.n397 gnd.n390 0.005
R1378 gnd.n390 gnd.n389 0.005
R1379 gnd.n389 gnd.n382 0.005
R1380 gnd.n382 gnd.n381 0.005
R1381 gnd.n381 gnd.n374 0.005
R1382 gnd.n374 gnd.n373 0.005
R1383 gnd.n373 gnd.n367 0.005
R1384 gnd.n367 gnd.n366 0.005
R1385 gnd.n366 gnd.n359 0.005
R1386 gnd.n359 gnd.n358 0.005
R1387 gnd.n358 gnd.n351 0.005
R1388 gnd.n351 gnd.n350 0.005
R1389 gnd.n350 gnd.n344 0.005
R1390 gnd.n344 gnd.n343 0.005
R1391 gnd.n343 gnd.n336 0.005
R1392 gnd.n336 gnd.n335 0.005
R1393 gnd.n335 gnd.n328 0.005
R1394 gnd.n328 gnd.n327 0.005
R1395 gnd.n327 gnd.n321 0.005
R1396 gnd.n321 gnd.n320 0.005
R1397 gnd.n320 gnd.n314 0.005
R1398 gnd.n314 gnd.n313 0.005
R1399 gnd.n313 gnd.n303 0.005
R1400 gnd.n303 gnd.n302 0.005
R1401 gnd.n302 gnd.n296 0.005
R1402 gnd.n296 gnd.n295 0.005
R1403 gnd.n295 gnd.n289 0.005
R1404 gnd.n289 gnd.n288 0.005
R1405 gnd.n1010 gnd.n1009 0.005
R1406 gnd.n1011 gnd.n553 0.004
R1407 gnd.n1010 gnd.n616 0.003
R1408 gnd.n479 gnd.n478 0.001
R1409 gnd.n452 gnd.n451 0.001
R1410 gnd.n178 gnd.n177 0.001
R1411 gnd.n205 gnd.n204 0.001
R1412 gnd.n231 gnd.n230 0.001
R1413 gnd.n223 gnd.n222 0.001
R1414 gnd.n214 gnd.n213 0.001
R1415 gnd.n196 gnd.n195 0.001
R1416 gnd.n187 gnd.n186 0.001
R1417 gnd.n169 gnd.n168 0.001
R1418 gnd.n443 gnd.n442 0.001
R1419 gnd.n461 gnd.n460 0.001
R1420 gnd.n470 gnd.n469 0.001
R1421 gnd.n488 gnd.n487 0.001
R1422 gnd.n497 gnd.n496 0.001
R1423 gnd.n505 gnd.n504 0.001
R1424 gnd.n553 gnd.n278 0.001
R1425 gnd.n553 gnd.n552 0.001
R1426 gate.n30 gate.t8 208.42
R1427 gate.n84 gate.t1 207.82
R1428 gate.n28 gate.t4 170.306
R1429 gate.n26 gate.t10 170.306
R1430 gate.n32 gate.t26 170.306
R1431 gate.n24 gate.t6 170.306
R1432 gate.n36 gate.t3 170.306
R1433 gate.n22 gate.t14 170.306
R1434 gate.n40 gate.t12 170.306
R1435 gate.n20 gate.t20 170.306
R1436 gate.n44 gate.t15 170.306
R1437 gate.n18 gate.t0 170.306
R1438 gate.n48 gate.t28 170.306
R1439 gate.n16 gate.t7 170.306
R1440 gate.n52 gate.t19 170.306
R1441 gate.n14 gate.t23 170.306
R1442 gate.n56 gate.t24 170.306
R1443 gate.n12 gate.t18 170.306
R1444 gate.n60 gate.t21 170.306
R1445 gate.n10 gate.t13 170.306
R1446 gate.n64 gate.t16 170.306
R1447 gate.n8 gate.t2 170.306
R1448 gate.n68 gate.t5 170.306
R1449 gate.n6 gate.t27 170.306
R1450 gate.n72 gate.t22 170.306
R1451 gate.n4 gate.t25 170.306
R1452 gate.n76 gate.t29 170.306
R1453 gate.n2 gate.t11 170.306
R1454 gate.n80 gate.t17 170.306
R1455 gate.n0 gate.t9 170.306
R1456 gate.n27 gate.n26 8.764
R1457 gate.n25 gate.n24 8.764
R1458 gate.n23 gate.n22 8.764
R1459 gate.n21 gate.n20 8.764
R1460 gate.n19 gate.n18 8.764
R1461 gate.n17 gate.n16 8.764
R1462 gate.n15 gate.n14 8.764
R1463 gate.n13 gate.n12 8.764
R1464 gate.n11 gate.n10 8.764
R1465 gate.n9 gate.n8 8.764
R1466 gate.n7 gate.n6 8.764
R1467 gate.n5 gate.n4 8.764
R1468 gate.n3 gate.n2 8.764
R1469 gate.n1 gate.n0 8.764
R1470 gate.n81 gate.n80 8.764
R1471 gate.n77 gate.n76 8.764
R1472 gate.n73 gate.n72 8.764
R1473 gate.n69 gate.n68 8.764
R1474 gate.n65 gate.n64 8.764
R1475 gate.n61 gate.n60 8.764
R1476 gate.n57 gate.n56 8.764
R1477 gate.n53 gate.n52 8.764
R1478 gate.n49 gate.n48 8.764
R1479 gate.n45 gate.n44 8.764
R1480 gate.n41 gate.n40 8.764
R1481 gate.n37 gate.n36 8.764
R1482 gate.n33 gate.n32 8.764
R1483 gate.n29 gate.n28 8.764
R1484 gate.n83 gate.n1 4.65
R1485 gate.n82 gate.n81 4.65
R1486 gate.n79 gate.n3 4.65
R1487 gate.n78 gate.n77 4.65
R1488 gate.n75 gate.n5 4.65
R1489 gate.n74 gate.n73 4.65
R1490 gate.n71 gate.n7 4.65
R1491 gate.n70 gate.n69 4.65
R1492 gate.n67 gate.n9 4.65
R1493 gate.n66 gate.n65 4.65
R1494 gate.n63 gate.n11 4.65
R1495 gate.n62 gate.n61 4.65
R1496 gate.n59 gate.n13 4.65
R1497 gate.n58 gate.n57 4.65
R1498 gate.n55 gate.n15 4.65
R1499 gate.n54 gate.n53 4.65
R1500 gate.n51 gate.n17 4.65
R1501 gate.n50 gate.n49 4.65
R1502 gate.n47 gate.n19 4.65
R1503 gate.n46 gate.n45 4.65
R1504 gate.n43 gate.n21 4.65
R1505 gate.n42 gate.n41 4.65
R1506 gate.n39 gate.n23 4.65
R1507 gate.n38 gate.n37 4.65
R1508 gate.n35 gate.n25 4.65
R1509 gate.n34 gate.n33 4.65
R1510 gate.n31 gate.n27 4.65
R1511 gate.n30 gate.n29 4.65
R1512 gate.n84 gate.n83 0.6
R1513 gate.n82 gate.n79 0.6
R1514 gate.n78 gate.n75 0.6
R1515 gate.n74 gate.n71 0.6
R1516 gate.n70 gate.n67 0.6
R1517 gate.n66 gate.n63 0.6
R1518 gate.n62 gate.n59 0.6
R1519 gate.n58 gate.n55 0.6
R1520 gate.n54 gate.n51 0.6
R1521 gate.n50 gate.n47 0.6
R1522 gate.n46 gate.n43 0.6
R1523 gate.n42 gate.n39 0.6
R1524 gate.n38 gate.n35 0.6
R1525 gate.n34 gate.n31 0.6
R1526 gate gate.n84 0.526
R1527 gate.n83 gate.n82 0.2
R1528 gate.n79 gate.n78 0.2
R1529 gate.n75 gate.n74 0.2
R1530 gate.n71 gate.n70 0.2
R1531 gate.n67 gate.n66 0.2
R1532 gate.n63 gate.n62 0.2
R1533 gate.n59 gate.n58 0.2
R1534 gate.n55 gate.n54 0.2
R1535 gate.n51 gate.n50 0.2
R1536 gate.n47 gate.n46 0.2
R1537 gate.n43 gate.n42 0.2
R1538 gate.n39 gate.n38 0.2
R1539 gate.n35 gate.n34 0.2
R1540 gate.n31 gate.n30 0.2
R1541 out.n63 out.t21 28.876
R1542 out.n141 out.t28 28.876
R1543 out.n54 out.t19 23.571
R1544 out.n54 out.t25 23.571
R1545 out.n45 out.t23 23.571
R1546 out.n45 out.t3 23.571
R1547 out.n36 out.t15 23.571
R1548 out.n36 out.t26 23.571
R1549 out.n27 out.t9 23.571
R1550 out.n27 out.t17 23.571
R1551 out.n18 out.t29 23.571
R1552 out.n18 out.t14 23.571
R1553 out.n9 out.t22 23.571
R1554 out.n9 out.t1 23.571
R1555 out.n0 out.t6 23.571
R1556 out.n0 out.t10 23.571
R1557 out.n78 out.t11 23.571
R1558 out.n78 out.t5 23.571
R1559 out.n87 out.t16 23.571
R1560 out.n87 out.t8 23.571
R1561 out.n96 out.t27 23.571
R1562 out.n96 out.t13 23.571
R1563 out.n105 out.t2 23.571
R1564 out.n105 out.t24 23.571
R1565 out.n114 out.t4 23.571
R1566 out.n114 out.t7 23.571
R1567 out.n123 out.t18 23.571
R1568 out.n123 out.t0 23.571
R1569 out.n132 out.t20 23.571
R1570 out.n132 out.t12 23.571
R1571 out.n146 out.n141 14.006
R1572 out.n68 out.n63 14.006
R1573 out.n60 out.n55 8.032
R1574 out.n51 out.n46 8.032
R1575 out.n42 out.n37 8.032
R1576 out.n33 out.n28 8.032
R1577 out.n24 out.n19 8.032
R1578 out.n15 out.n10 8.032
R1579 out.n6 out.n1 8.032
R1580 out.n84 out.n79 8.032
R1581 out.n93 out.n88 8.032
R1582 out.n102 out.n97 8.032
R1583 out.n111 out.n106 8.032
R1584 out.n120 out.n115 8.032
R1585 out.n129 out.n124 8.032
R1586 out.n138 out.n133 8.032
R1587 out.n65 out.n64 3.85
R1588 out.n57 out.n56 3.85
R1589 out.n48 out.n47 3.85
R1590 out.n39 out.n38 3.85
R1591 out.n30 out.n29 3.85
R1592 out.n21 out.n20 3.85
R1593 out.n12 out.n11 3.85
R1594 out.n3 out.n2 3.85
R1595 out.n81 out.n80 3.85
R1596 out.n90 out.n89 3.85
R1597 out.n99 out.n98 3.85
R1598 out.n108 out.n107 3.85
R1599 out.n117 out.n116 3.85
R1600 out.n126 out.n125 3.85
R1601 out.n135 out.n134 3.85
R1602 out.n143 out.n142 3.85
R1603 out.n55 out.n54 1.601
R1604 out.n46 out.n45 1.601
R1605 out.n37 out.n36 1.601
R1606 out.n28 out.n27 1.601
R1607 out.n19 out.n18 1.601
R1608 out.n10 out.n9 1.601
R1609 out.n1 out.n0 1.601
R1610 out.n79 out.n78 1.601
R1611 out.n88 out.n87 1.601
R1612 out.n97 out.n96 1.601
R1613 out.n106 out.n105 1.601
R1614 out.n115 out.n114 1.601
R1615 out.n124 out.n123 1.601
R1616 out.n133 out.n132 1.601
R1617 out.n71 out.n70 1.49
R1618 out.n149 out.n148 1.49
R1619 out.n71 out.n62 1.369
R1620 out.n72 out.n53 1.369
R1621 out.n73 out.n44 1.369
R1622 out.n74 out.n35 1.369
R1623 out.n75 out.n26 1.369
R1624 out.n76 out.n17 1.369
R1625 out.n77 out.n8 1.369
R1626 out.n155 out.n86 1.369
R1627 out.n154 out.n95 1.369
R1628 out.n153 out.n104 1.369
R1629 out.n152 out.n113 1.369
R1630 out.n151 out.n122 1.369
R1631 out.n150 out.n131 1.369
R1632 out.n149 out.n140 1.369
R1633 out.n69 out.n68 0.619
R1634 out.n61 out.n60 0.618
R1635 out.n52 out.n51 0.618
R1636 out.n43 out.n42 0.618
R1637 out.n34 out.n33 0.618
R1638 out.n25 out.n24 0.618
R1639 out.n16 out.n15 0.618
R1640 out.n7 out.n6 0.618
R1641 out.n85 out.n84 0.618
R1642 out.n94 out.n93 0.618
R1643 out.n103 out.n102 0.618
R1644 out.n112 out.n111 0.618
R1645 out.n121 out.n120 0.618
R1646 out.n130 out.n129 0.618
R1647 out.n139 out.n138 0.618
R1648 out.n147 out.n146 0.618
R1649 out.n150 out.n149 0.121
R1650 out.n151 out.n150 0.121
R1651 out.n152 out.n151 0.121
R1652 out.n153 out.n152 0.121
R1653 out.n154 out.n153 0.121
R1654 out.n155 out.n154 0.121
R1655 out.n77 out.n76 0.121
R1656 out.n76 out.n75 0.121
R1657 out.n75 out.n74 0.121
R1658 out.n74 out.n73 0.121
R1659 out.n73 out.n72 0.121
R1660 out.n72 out.n71 0.121
R1661 out.n68 out.n67 0.098
R1662 out.n60 out.n59 0.098
R1663 out.n51 out.n50 0.098
R1664 out.n42 out.n41 0.098
R1665 out.n33 out.n32 0.098
R1666 out.n24 out.n23 0.098
R1667 out.n15 out.n14 0.098
R1668 out.n6 out.n5 0.098
R1669 out.n84 out.n83 0.098
R1670 out.n93 out.n92 0.098
R1671 out.n102 out.n101 0.098
R1672 out.n111 out.n110 0.098
R1673 out.n120 out.n119 0.098
R1674 out.n129 out.n128 0.098
R1675 out.n138 out.n137 0.098
R1676 out.n146 out.n145 0.098
R1677 out.n156 out.n155 0.06
R1678 out.n156 out.n77 0.06
R1679 out.n70 out.n69 0.037
R1680 out.n62 out.n61 0.037
R1681 out.n53 out.n52 0.037
R1682 out.n44 out.n43 0.037
R1683 out.n35 out.n34 0.037
R1684 out.n26 out.n25 0.037
R1685 out.n17 out.n16 0.037
R1686 out.n8 out.n7 0.037
R1687 out.n86 out.n85 0.037
R1688 out.n95 out.n94 0.037
R1689 out.n104 out.n103 0.037
R1690 out.n113 out.n112 0.037
R1691 out.n122 out.n121 0.037
R1692 out.n131 out.n130 0.037
R1693 out.n140 out.n139 0.037
R1694 out.n148 out.n147 0.037
R1695 out out.n156 0.033
R1696 out.n66 out.n65 0.008
R1697 out.n58 out.n57 0.008
R1698 out.n49 out.n48 0.008
R1699 out.n40 out.n39 0.008
R1700 out.n31 out.n30 0.008
R1701 out.n22 out.n21 0.008
R1702 out.n13 out.n12 0.008
R1703 out.n4 out.n3 0.008
R1704 out.n82 out.n81 0.008
R1705 out.n91 out.n90 0.008
R1706 out.n100 out.n99 0.008
R1707 out.n109 out.n108 0.008
R1708 out.n118 out.n117 0.008
R1709 out.n127 out.n126 0.008
R1710 out.n136 out.n135 0.008
R1711 out.n144 out.n143 0.008
R1712 out.n67 out.n66 0.001
R1713 out.n59 out.n58 0.001
R1714 out.n50 out.n49 0.001
R1715 out.n41 out.n40 0.001
R1716 out.n32 out.n31 0.001
R1717 out.n23 out.n22 0.001
R1718 out.n14 out.n13 0.001
R1719 out.n5 out.n4 0.001
R1720 out.n83 out.n82 0.001
R1721 out.n92 out.n91 0.001
R1722 out.n101 out.n100 0.001
R1723 out.n110 out.n109 0.001
R1724 out.n119 out.n118 0.001
R1725 out.n128 out.n127 0.001
R1726 out.n137 out.n136 0.001
R1727 out.n145 out.n144 0.001
R1728 in.n0 in.t12 208.341
R1729 in.n14 in.t11 208.341
R1730 in.n13 in.t15 207.82
R1731 in.n12 in.t22 207.82
R1732 in.n11 in.t23 207.82
R1733 in.n10 in.t16 207.82
R1734 in.n9 in.t26 207.82
R1735 in.n8 in.t6 207.82
R1736 in.n7 in.t18 207.82
R1737 in.n6 in.t27 207.82
R1738 in.n5 in.t1 207.82
R1739 in.n4 in.t0 207.82
R1740 in.n3 in.t4 207.82
R1741 in.n2 in.t8 207.82
R1742 in.n1 in.t9 207.82
R1743 in.n0 in.t13 207.82
R1744 in.n14 in.t10 207.82
R1745 in.n15 in.t7 207.82
R1746 in.n16 in.t5 207.82
R1747 in.n17 in.t3 207.82
R1748 in.n18 in.t2 207.82
R1749 in.n19 in.t20 207.82
R1750 in.n20 in.t19 207.82
R1751 in.n21 in.t29 207.82
R1752 in.n22 in.t17 207.82
R1753 in.n23 in.t25 207.82
R1754 in.n24 in.t24 207.82
R1755 in.n25 in.t28 207.82
R1756 in.n26 in.t21 207.82
R1757 in.n27 in.t14 207.82
R1758 in.n28 in.n13 0.74
R1759 in.n1 in.n0 0.521
R1760 in.n2 in.n1 0.521
R1761 in.n3 in.n2 0.521
R1762 in.n4 in.n3 0.521
R1763 in.n5 in.n4 0.521
R1764 in.n6 in.n5 0.521
R1765 in.n7 in.n6 0.521
R1766 in.n8 in.n7 0.521
R1767 in.n9 in.n8 0.521
R1768 in.n10 in.n9 0.521
R1769 in.n11 in.n10 0.521
R1770 in.n12 in.n11 0.521
R1771 in.n13 in.n12 0.521
R1772 in.n15 in.n14 0.521
R1773 in.n16 in.n15 0.521
R1774 in.n17 in.n16 0.521
R1775 in.n18 in.n17 0.521
R1776 in.n19 in.n18 0.521
R1777 in.n20 in.n19 0.521
R1778 in.n21 in.n20 0.521
R1779 in.n22 in.n21 0.521
R1780 in.n23 in.n22 0.521
R1781 in.n24 in.n23 0.521
R1782 in.n25 in.n24 0.521
R1783 in.n26 in.n25 0.521
R1784 in.n27 in.n26 0.521
R1785 in.n28 in.n27 0.48
R1786 in.n34 in.n30 0.261
R1787 in.n33 in.n31 0.233
R1788 in.n33 in.n32 0.124
R1789 in.n30 in.n29 0.088
R1790 in.n34 in.n33 0.088
R1791 in.n35 in.n34 0.077
R1792 in.n29 in.n28 0.027
R1793 in.n35 in 0.001
C0 gate in 0.02963fF
C1 out Vctrl 1.44433fF
C2 a_n2543_2314# Vctrl 1.96910fF
C3 out Vdd 7.69784fF
C4 Vdd a_n2543_2314# 13.20780fF
C5 out in 0.00147fF
C6 gate out 0.89442fF
C7 in a_n2543_2314# 2.82331fF
C8 gate a_n2543_2314# 3.07244fF
C9 out a_n2543_2314# 12.68150fF
C10 Vdd Vctrl 1.91398fF
C11 gate Vctrl 0.58769fF
C12 gate Vdd 0.49363fF
