.subckt VGA_final RF_in Gnd RF_out Vdd_1v8 Vgg_1v2 Vctrl
*.PININFO RF_in:B Gnd:B RF_out:B Vdd_1v8:B Vgg_1v2:B Vctrl:B
x1 Vdd_1v8 Vdd_1v8 Vdd_1v8 Vctrl_in gate1_in Gnd VGA_gainCellv3
XC1 gate1_in RF_in sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC2 Gnd gate1_in sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC3 Gnd gate1_in sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC4 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC5 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC6 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC7 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC8 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XC9 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 W=15 L=15 MF=1 m=1
XM1 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
R1 Vgg_1v2 gate1_in sky130_fd_pr__res_generic_po W=2 L=10.53 mult=1 m=1
XM3 gate1_in Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 gate1_in Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM5 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM6 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
R2 Vctrl Vctrl_in sky130_fd_pr__res_generic_po W=2 L=10.53 mult=1 m=1
XM7 Vctrl_in Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM8 Vctrl_in Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM9 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM10 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt L=1 W=112.2 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
x2 RF_out Vdd_1v8 Gnd MOM_capacitor
.ends

* expanding   symbol:
*+  /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/VGA_core/VGA_gainCellv3.sym # of pins=6
* sym_path:
*+ /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/VGA_core/VGA_gainCellv3.sym
* sch_path:
*+ /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/VGA_core/VGA_gainCellv3.sch
.subckt VGA_gainCellv3  out Vdd gate Vctrl in gnd
*.PININFO in:B out:B gate:B Vdd:B Vctrl:B gnd:B
XM1 net1 in gnd gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=25.2 nf=30 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out gate net1 gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=25.2 nf=30 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 Vdd Vctrl net1 gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=25.2 nf=30 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM5 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM6 gnd gnd net1 gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM7 gnd gnd net1 gnd sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XC1 Vctrl gnd sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
XC2 Vdd gnd sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
D1 gnd in sky130_fd_pr__diode_pw2nd_05v5 area=202.5m
D2 gnd gate sky130_fd_pr__diode_pw2nd_05v5 area=202.5m
D3 gnd Vctrl sky130_fd_pr__diode_pw2nd_05v5 area=202.5m
.ends


* expanding   symbol:
*+  /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/MOM_capacitor.sym # of pins=3
* sym_path: /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/MOM_capacitor.sym
* sch_path: /home/leonardo/sky130_projects/SSCS_PICO_tapeout/VGA_tapeout/xschem/MOM_capacitor.sch
.subckt MOM_capacitor  out in gnd
*.PININFO in:B out:B gnd:B
.ends

** flattened .save nodes
.end
