* SPICE3 file created from core_v3.ext - technology: sky130A

X0 source.t27 bias1_inputa.t0 a_85_n463.t27 bulk.t348 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs0 bias1_input.t0 bias1_inputa.t0 434.216
X1 bulk bulk.t309 bulk bulk.t310 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 bulk.t308 bulk.t305 bulk.t307 bulk.t306 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 bulk bulk.t300 bulk bulk.t301 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 source.t26 bias1_inputa.t1 a_85_n463.t28 bulk.t347 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs4 bias1_input.t1 bias1_inputa.t1 434.216
X5 bulk bulk.t295 bulk bulk.t296 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 bulk.t294 bulk.t291 bulk.t293 bulk.t292 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 bulk bulk.t286 bulk bulk.t287 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 bulk bulk.t281 bulk bulk.t282 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_85_n463.t18 bias1_inputa.t2 source.t25 bulk.t346 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs9 bias1_input.t2 bias1_inputa.t2 434.216
X10 a_85_n463.t15 bias1_inputa.t3 source.t24 bulk.t345 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs10 bias1_input.t3 bias1_inputa.t3 434.216
X11 a_85_n463.t6 bias2a.t0 tank_out.t27 bulk.t316 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs11 bias2.t0 bias2a.t0 402.18
X12 source.t23 bias1_inputa.t4 a_85_n463.t12 bulk.t344 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs12 bias1_input.t4 bias1_inputa.t4 434.216
X13 tank_out.t26 bias2.t1 a_85_n463.t5 bulk.t315 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs13 bias2.t1 bias2a.t1 402.18
X14 a_85_n463.t9 bias2a.t2 tank_out.t25 bulk.t319 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs14 bias2.t2 bias2a.t2 402.18
X15 tank_out.t24 bias2a.t3 a_85_n463.t44 bulk.t354 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs15 bias2.t3 bias2a.t3 402.18
X16 a_85_n463.t40 bias2a.t4 tank_out.t23 bulk.t350 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs16 bias2.t4 bias2a.t4 402.18
X17 a_85_n463.t46 bias2a.t5 tank_out.t22 bulk.t356 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs17 bias2.t5 bias2a.t5 402.18
X18 tank_out.t21 bias2a.t6 a_85_n463.t41 bulk.t351 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs18 bias2.t6 bias2a.t6 402.18
X19 tank_out.t20 bias2a.t7 a_85_n463.t50 bulk.t360 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs19 bias2.t7 bias2a.t7 402.18
X20 source.t22 bias1_inputa.t5 a_85_n463.t36 bulk.t343 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs20 bias1_input.t5 bias1_inputa.t5 434.216
X21 source.t21 bias1_inputa.t6 a_85_n463.t34 bulk.t342 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs21 bias1_input.t6 bias1_inputa.t6 434.216
X22 a_85_n463.t37 bias1_inputa.t7 source.t20 bulk.t341 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs22 bias1_input.t7 bias1_inputa.t7 434.216
X23 a_85_n463.t23 bias1_inputa.t8 source.t19 bulk.t340 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs23 bias1_input.t8 bias1_inputa.t8 434.216
X24 a_85_n463.t47 bias2a.t8 tank_out.t19 bulk.t357 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs24 bias2.t8 bias2a.t8 402.18
X25 tank_out.t18 bias2a.t9 a_85_n463.t8 bulk.t318 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs25 bias2.t9 bias2a.t9 402.18
X26 a_85_n463.t21 bias1_inputa.t9 source.t18 bulk.t339 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs26 bias1_input.t9 bias1_inputa.t9 434.216
X27 a_85_n463.t55 bias2a.t10 tank_out.t17 bulk.t365 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs27 bias2.t10 bias2a.t10 402.18
X28 tank_out.t16 bias2a.t11 a_85_n463.t3 bulk.t3 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs28 bias2.t11 bias2a.t11 402.18
X29 a_85_n463.t54 bias2a.t12 tank_out.t15 bulk.t364 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs29 bias2.t12 bias2a.t12 402.18
X30 bulk bulk.t276 bulk bulk.t277 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_85_n463.t53 bias2a.t13 tank_out.t14 bulk.t363 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs31 bias2.t13 bias2a.t13 402.18
X32 tank_out.t13 bias2a.t14 a_85_n463.t48 bulk.t358 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs32 bias2.t14 bias2a.t14 402.18
X33 a_85_n463.t52 bias2a.t15 tank_out.t12 bulk.t362 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs33 bias2.t15 bias2a.t15 402.18
X34 source.t17 bias1_inputa.t10 a_85_n463.t30 bulk.t338 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs34 bias1_input.t10 bias1_inputa.t10 434.216
X35 tank_out.t11 bias2a.t16 a_85_n463.t51 bulk.t361 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs35 bias2.t16 bias2a.t16 402.18
X36 source.t16 bias1_inputa.t11 a_85_n463.t14 bulk.t337 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs36 bias1_input.t11 bias1_inputa.t11 434.216
X37 bulk.t275 bulk.t272 bulk.t274 bulk.t273 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 source.t15 bias1_inputa.t12 a_85_n463.t33 bulk.t336 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs38 bias1_input.t12 bias1_inputa.t12 434.216
X39 tank_out.t10 bias2a.t17 a_85_n463.t42 bulk.t352 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs39 bias2.t17 bias2a.t17 402.18
X40 bulk bulk.t267 bulk bulk.t268 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 tank_out.t9 bias2a.t18 a_85_n463.t45 bulk.t355 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs41 bias2.t18 bias2a.t18 402.18
X42 a_85_n463.t43 bias2a.t19 tank_out.t8 bulk.t353 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs42 bias2.t19 bias2a.t19 402.18
X43 bulk bulk.t262 bulk bulk.t263 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 bulk bulk.t257 bulk bulk.t258 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_85_n463.t31 bias1_inputa.t13 source.t14 bulk.t335 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs45 bias1_input.t13 bias1_inputa.t13 434.216
X46 bulk bulk.t252 bulk bulk.t253 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 bulk.t251 bulk.t248 bulk.t250 bulk.t249 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_85_n463.t38 bias1_inputa.t14 source.t13 bulk.t334 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs48 bias1_input.t14 bias1_inputa.t14 434.216
X49 bulk bulk.t243 bulk bulk.t244 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 source.t12 bias1_inputa.t15 a_85_n463.t17 bulk.t333 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs50 bias1_input.t15 bias1_inputa.t15 434.216
X51 bulk bulk.t238 bulk bulk.t239 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 bulk bulk.t233 bulk bulk.t234 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 bulk bulk.t228 bulk bulk.t229 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 bulk bulk.t223 bulk bulk.t224 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 bulk bulk.t218 bulk bulk.t219 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 bulk bulk.t213 bulk bulk.t214 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 bulk bulk.t208 bulk bulk.t209 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 bulk bulk.t203 bulk bulk.t204 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 bulk bulk.t198 bulk bulk.t199 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 bulk.t197 bulk.t194 bulk.t196 bulk.t195 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 bulk bulk.t189 bulk bulk.t190 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 source.t11 bias1_inputa.t16 a_85_n463.t22 bulk.t332 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs62 bias1_input.t16 bias1_inputa.t16 434.216
X63 source.t10 bias1_inputa.t17 a_85_n463.t25 bulk.t331 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs63 bias1_input.t17 bias1_inputa.t17 434.216
X64 a_85_n463.t32 bias1_inputa.t18 source.t9 bulk.t330 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs64 bias1_input.t18 bias1_inputa.t18 434.216
X65 bulk bulk.t184 bulk bulk.t185 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 bulk bulk.t179 bulk bulk.t180 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 bulk bulk.t174 bulk bulk.t175 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 bulk bulk.t169 bulk bulk.t170 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 a_85_n463.t29 bias1_inputa.t19 source.t8 bulk.t329 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs69 bias1_input.t19 bias1_inputa.t19 434.216
X70 bulk bulk.t164 bulk bulk.t165 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 bulk.t163 bulk.t160 bulk.t162 bulk.t161 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 bulk.t159 bulk.t156 bulk.t158 bulk.t157 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 bulk bulk.t151 bulk bulk.t152 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 bulk bulk.t146 bulk bulk.t147 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 bulk bulk.t141 bulk bulk.t142 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 bulk bulk.t136 bulk bulk.t137 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 bulk bulk.t131 bulk bulk.t132 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 bulk bulk.t126 bulk bulk.t127 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 bulk bulk.t121 bulk bulk.t122 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 bulk bulk.t116 bulk bulk.t117 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 bulk bulk.t111 bulk bulk.t112 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 bulk bulk.t106 bulk bulk.t107 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 a_85_n463.t11 bias1_inputa.t20 source.t7 bulk.t328 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs83 bias1_input.t20 bias1_inputa.t20 434.216
X84 a_85_n463.t26 bias1_inputa.t21 source.t6 bulk.t327 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs84 bias1_input.t21 bias1_inputa.t21 434.216
X85 source.t5 bias1_inputa.t22 a_85_n463.t13 bulk.t326 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs85 bias1_input.t22 bias1_inputa.t22 434.216
X86 bulk bulk.t101 bulk bulk.t102 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 bulk bulk.t96 bulk bulk.t97 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 bulk.t95 bulk.t92 bulk.t94 bulk.t93 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X89 bulk bulk.t87 bulk bulk.t88 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X90 bulk bulk.t82 bulk bulk.t83 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 a_85_n463.t19 bias1_inputa.t23 source.t4 bulk.t325 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs91 bias1_input.t23 bias1_inputa.t23 434.216
X92 a_85_n463.t20 bias1_inputa.t24 source.t3 bulk.t324 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs92 bias1_input.t24 bias1_inputa.t24 434.216
X93 bulk bulk.t77 bulk bulk.t78 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 bulk bulk.t72 bulk bulk.t73 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 bulk bulk.t67 bulk bulk.t68 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 bulk bulk.t62 bulk bulk.t63 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 bulk.t61 bulk.t58 bulk.t60 bulk.t59 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 bulk bulk.t53 bulk bulk.t54 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 source.t2 bias1_inputa.t25 a_85_n463.t16 bulk.t323 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs99 bias1_input.t25 bias1_inputa.t25 434.216
X100 bulk bulk.t48 bulk bulk.t49 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 source.t1 bias1_inputa.t26 a_85_n463.t35 bulk.t322 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs101 bias1_input.t26 bias1_inputa.t26 434.216
X102 a_85_n463.t2 bias2a.t20 tank_out.t7 bulk.t2 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs102 bias2.t20 bias2a.t20 402.18
X103 tank_out.t6 bias2a.t21 a_85_n463.t4 bulk.t314 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs103 bias2.t21 bias2a.t21 402.18
X104 bulk bulk.t43 bulk bulk.t44 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 a_85_n463.t39 bias2a.t22 tank_out.t5 bulk.t349 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs105 bias2.t22 bias2a.t22 402.18
X106 bulk bulk.t38 bulk bulk.t39 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 bulk bulk.t33 bulk bulk.t34 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X108 a_85_n463.t24 bias1_inputa.t27 source.t0 bulk.t321 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs108 bias1_input.t27 bias1_inputa.t27 434.216
X109 a_85_n463.t10 bias2a.t23 tank_out.t4 bulk.t320 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs109 bias2.t23 bias2a.t23 402.18
X110 tank_out.t3 bias2a.t24 a_85_n463.t0 bulk.t0 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs110 bias2.t24 bias2a.t24 402.18
X111 bulk bulk.t28 bulk bulk.t29 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 tank_out.t2 bias2a.t25 a_85_n463.t49 bulk.t359 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs112 bias2.t25 bias2a.t25 402.18
X113 a_85_n463.t7 bias2a.t26 tank_out.t1 bulk.t317 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs113 bias2.t26 bias2a.t26 402.18
X114 bulk bulk.t23 bulk bulk.t24 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 bulk bulk.t18 bulk bulk.t19 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 tank_out.t0 bias2a.t27 a_85_n463.t1 bulk.t1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
Rnqs116 bias2.t27 bias2a.t27 402.18
X117 bulk.t17 bulk.t14 bulk.t16 bulk.t15 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 bulk bulk.t9 bulk bulk.t10 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 bulk bulk.t4 bulk bulk.t5 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 bias1_input source 3.75508fF
C1 bias2 tank_out 5.19660fF
C2 bias2 bias1_input 1.73261fF
C3 tank_out bias1_input 0.00402fF
C4 bias2 source 0.00402fF
C5 tank_out source 0.47754fF
R0 bias1_input.n89 bias1_input.t10 286.107
R1 bias1_input.n90 bias1_input.t0 286.107
R2 bias1_input.n91 bias1_input.t15 286.107
R3 bias1_input.n92 bias1_input.t4 286.107
R4 bias1_input.n93 bias1_input.t16 286.107
R5 bias1_input.n94 bias1_input.t5 286.107
R6 bias1_input.n95 bias1_input.t25 286.107
R7 bias1_input.n96 bias1_input.t11 286.107
R8 bias1_input.n97 bias1_input.t22 286.107
R9 bias1_input.n98 bias1_input.t17 286.107
R10 bias1_input.n99 bias1_input.t6 286.107
R11 bias1_input.n100 bias1_input.t26 286.107
R12 bias1_input.n101 bias1_input.t12 286.107
R13 bias1_input.n102 bias1_input.t1 286.107
R14 bias1_input.n43 bias1_input.t24 233.526
R15 bias1_input.n42 bias1_input.t3 233.526
R16 bias1_input.n41 bias1_input.t14 233.526
R17 bias1_input.n40 bias1_input.t21 233.526
R18 bias1_input.n39 bias1_input.t8 233.526
R19 bias1_input.n38 bias1_input.t19 233.526
R20 bias1_input.n37 bias1_input.t2 233.526
R21 bias1_input.n36 bias1_input.t13 233.526
R22 bias1_input.n35 bias1_input.t20 233.526
R23 bias1_input.n34 bias1_input.t9 233.526
R24 bias1_input.n33 bias1_input.t27 233.526
R25 bias1_input.n32 bias1_input.t7 233.526
R26 bias1_input.n31 bias1_input.t18 233.526
R27 bias1_input.n30 bias1_input.t23 233.526
R28 bias1_input.n112 bias1_input.n111 1.143
R29 bias1_input.n52 bias1_input.n51 1.143
R30 bias1_input.n65 bias1_input.n64 1.137
R31 bias1_input.n5 bias1_input.n4 1.137
R32 bias1_input.n47 bias1_input.n46 1.137
R33 bias1_input.n20 bias1_input.n19 1.137
R34 bias1_input.n14 bias1_input.n13 1.137
R35 bias1_input.n80 bias1_input.n79 1.137
R36 bias1_input.n107 bias1_input.n106 1.137
R37 bias1_input.n74 bias1_input.n73 1.137
R38 bias1_input.n45 bias1_input.n44 0.963
R39 bias1_input.n104 bias1_input.n103 0.963
R40 bias1_input.n53 bias1_input.n52 0.687
R41 bias1_input.n113 bias1_input.n112 0.687
R42 bias1_input.n44 bias1_input.n43 0.293
R43 bias1_input.n90 bias1_input.n89 0.203
R44 bias1_input.n91 bias1_input.n90 0.203
R45 bias1_input.n92 bias1_input.n91 0.203
R46 bias1_input.n93 bias1_input.n92 0.203
R47 bias1_input.n94 bias1_input.n93 0.203
R48 bias1_input.n95 bias1_input.n94 0.203
R49 bias1_input.n96 bias1_input.n95 0.203
R50 bias1_input.n97 bias1_input.n96 0.203
R51 bias1_input.n98 bias1_input.n97 0.203
R52 bias1_input.n99 bias1_input.n98 0.203
R53 bias1_input.n100 bias1_input.n99 0.203
R54 bias1_input.n101 bias1_input.n100 0.203
R55 bias1_input.n102 bias1_input.n101 0.203
R56 bias1_input.n31 bias1_input.n30 0.203
R57 bias1_input.n32 bias1_input.n31 0.203
R58 bias1_input.n33 bias1_input.n32 0.203
R59 bias1_input.n34 bias1_input.n33 0.203
R60 bias1_input.n35 bias1_input.n34 0.203
R61 bias1_input.n36 bias1_input.n35 0.203
R62 bias1_input.n37 bias1_input.n36 0.203
R63 bias1_input.n38 bias1_input.n37 0.203
R64 bias1_input.n39 bias1_input.n38 0.203
R65 bias1_input.n40 bias1_input.n39 0.203
R66 bias1_input.n41 bias1_input.n40 0.203
R67 bias1_input.n42 bias1_input.n41 0.203
R68 bias1_input.n43 bias1_input.n42 0.203
R69 bias1_input.n103 bias1_input.n102 0.191
R70 bias1_input bias1_input.n120 0.087
R71 bias1_input.n27 bias1_input.n26 0.048
R72 bias1_input.n86 bias1_input.n85 0.048
R73 bias1_input.n44 bias1_input.n29 0.026
R74 bias1_input.n103 bias1_input.n88 0.026
R75 bias1_input.n25 bias1_input.n24 0.024
R76 bias1_input.n84 bias1_input.n83 0.024
R77 bias1_input.n3 bias1_input.n2 0.024
R78 bias1_input.n62 bias1_input.n61 0.024
R79 bias1_input.n46 bias1_input.n45 0.021
R80 bias1_input.n106 bias1_input.n104 0.021
R81 bias1_input.n11 bias1_input.n10 0.019
R82 bias1_input.n71 bias1_input.n70 0.019
R83 bias1_input.n28 bias1_input.n27 0.015
R84 bias1_input.n87 bias1_input.n86 0.015
R85 bias1_input.n12 bias1_input.n11 0.015
R86 bias1_input.n72 bias1_input.n71 0.015
R87 bias1_input.n51 bias1_input.n50 0.013
R88 bias1_input.n46 bias1_input.n23 0.013
R89 bias1_input.n19 bias1_input.n18 0.013
R90 bias1_input.n79 bias1_input.n78 0.013
R91 bias1_input.n106 bias1_input.n105 0.013
R92 bias1_input.n111 bias1_input.n110 0.013
R93 bias1_input.n29 bias1_input.n28 0.011
R94 bias1_input.n88 bias1_input.n87 0.011
R95 bias1_input.n13 bias1_input.n12 0.011
R96 bias1_input.n73 bias1_input.n72 0.011
R97 bias1_input.n7 bias1_input.n6 0.009
R98 bias1_input.n5 bias1_input.n0 0.009
R99 bias1_input.n65 bias1_input.n60 0.009
R100 bias1_input.n67 bias1_input.n66 0.009
R101 bias1_input.n18 bias1_input.n17 0.008
R102 bias1_input.n78 bias1_input.n77 0.008
R103 bias1_input.n22 bias1_input.n21 0.007
R104 bias1_input.n9 bias1_input.n8 0.007
R105 bias1_input.n69 bias1_input.n68 0.007
R106 bias1_input.n82 bias1_input.n81 0.007
R107 bias1_input.n14 bias1_input.n9 0.006
R108 bias1_input.n74 bias1_input.n69 0.006
R109 bias1_input.n4 bias1_input.n1 0.005
R110 bias1_input.n64 bias1_input.n63 0.005
R111 bias1_input.n48 bias1_input.n47 0.005
R112 bias1_input.n20 bias1_input.n16 0.005
R113 bias1_input.n15 bias1_input.n14 0.005
R114 bias1_input.n75 bias1_input.n74 0.005
R115 bias1_input.n80 bias1_input.n76 0.005
R116 bias1_input.n108 bias1_input.n107 0.005
R117 bias1_input.n55 bias1_input.n54 0.005
R118 bias1_input.n56 bias1_input.n55 0.005
R119 bias1_input.n58 bias1_input.n57 0.005
R120 bias1_input.n59 bias1_input.n58 0.005
R121 bias1_input.n119 bias1_input.n118 0.005
R122 bias1_input.n118 bias1_input.n117 0.005
R123 bias1_input.n116 bias1_input.n115 0.005
R124 bias1_input.n115 bias1_input.n114 0.005
R125 bias1_input.n26 bias1_input.n25 0.003
R126 bias1_input.n85 bias1_input.n84 0.003
R127 bias1_input.n4 bias1_input.n3 0.003
R128 bias1_input.n64 bias1_input.n62 0.003
R129 bias1_input.n49 bias1_input.n48 0.003
R130 bias1_input.n47 bias1_input.n22 0.003
R131 bias1_input.n21 bias1_input.n20 0.003
R132 bias1_input.n16 bias1_input.n15 0.003
R133 bias1_input.n76 bias1_input.n75 0.003
R134 bias1_input.n81 bias1_input.n80 0.003
R135 bias1_input.n107 bias1_input.n82 0.003
R136 bias1_input.n109 bias1_input.n108 0.003
R137 bias1_input.n54 bias1_input.n53 0.003
R138 bias1_input.n57 bias1_input.n56 0.003
R139 bias1_input.n117 bias1_input.n116 0.003
R140 bias1_input.n114 bias1_input.n113 0.003
R141 bias1_input.n52 bias1_input.n49 0.002
R142 bias1_input.n112 bias1_input.n109 0.002
R143 bias1_input.n8 bias1_input.n7 0.002
R144 bias1_input.n68 bias1_input.n67 0.002
R145 bias1_input.n6 bias1_input.n5 0.001
R146 bias1_input.n66 bias1_input.n65 0.001
R147 bias1_input.n120 bias1_input.n59 0.001
R148 bias1_input.n120 bias1_input.n119 0.001
R149 a_85_n463.n20 a_85_n463.t1 19.8
R150 a_85_n463.n20 a_85_n463.t10 19.8
R151 a_85_n463.n33 a_85_n463.t49 19.8
R152 a_85_n463.n33 a_85_n463.t2 19.8
R153 a_85_n463.n46 a_85_n463.t4 19.8
R154 a_85_n463.n46 a_85_n463.t39 19.8
R155 a_85_n463.n59 a_85_n463.t5 19.8
R156 a_85_n463.n59 a_85_n463.t46 19.8
R157 a_85_n463.n72 a_85_n463.t50 19.8
R158 a_85_n463.n72 a_85_n463.t9 19.8
R159 a_85_n463.n85 a_85_n463.t41 19.8
R160 a_85_n463.n85 a_85_n463.t6 19.8
R161 a_85_n463.n98 a_85_n463.t44 19.8
R162 a_85_n463.n98 a_85_n463.t40 19.8
R163 a_85_n463.n111 a_85_n463.t45 19.8
R164 a_85_n463.n111 a_85_n463.t43 19.8
R165 a_85_n463.n124 a_85_n463.t42 19.8
R166 a_85_n463.n124 a_85_n463.t53 19.8
R167 a_85_n463.n137 a_85_n463.t51 19.8
R168 a_85_n463.n137 a_85_n463.t55 19.8
R169 a_85_n463.n150 a_85_n463.t48 19.8
R170 a_85_n463.n150 a_85_n463.t47 19.8
R171 a_85_n463.n163 a_85_n463.t3 19.8
R172 a_85_n463.n163 a_85_n463.t52 19.8
R173 a_85_n463.n176 a_85_n463.t8 19.8
R174 a_85_n463.n176 a_85_n463.t54 19.8
R175 a_85_n463.n441 a_85_n463.t28 19.8
R176 a_85_n463.n426 a_85_n463.t33 19.8
R177 a_85_n463.n426 a_85_n463.t20 19.8
R178 a_85_n463.n411 a_85_n463.t35 19.8
R179 a_85_n463.n411 a_85_n463.t15 19.8
R180 a_85_n463.n396 a_85_n463.t34 19.8
R181 a_85_n463.n396 a_85_n463.t38 19.8
R182 a_85_n463.n381 a_85_n463.t25 19.8
R183 a_85_n463.n381 a_85_n463.t26 19.8
R184 a_85_n463.n366 a_85_n463.t13 19.8
R185 a_85_n463.n366 a_85_n463.t23 19.8
R186 a_85_n463.n351 a_85_n463.t14 19.8
R187 a_85_n463.n351 a_85_n463.t29 19.8
R188 a_85_n463.n336 a_85_n463.t16 19.8
R189 a_85_n463.n336 a_85_n463.t18 19.8
R190 a_85_n463.n321 a_85_n463.t36 19.8
R191 a_85_n463.n321 a_85_n463.t31 19.8
R192 a_85_n463.n306 a_85_n463.t22 19.8
R193 a_85_n463.n306 a_85_n463.t11 19.8
R194 a_85_n463.n291 a_85_n463.t12 19.8
R195 a_85_n463.n291 a_85_n463.t21 19.8
R196 a_85_n463.n276 a_85_n463.t17 19.8
R197 a_85_n463.n276 a_85_n463.t24 19.8
R198 a_85_n463.n229 a_85_n463.t27 19.8
R199 a_85_n463.n229 a_85_n463.t37 19.8
R200 a_85_n463.n244 a_85_n463.t30 19.8
R201 a_85_n463.n244 a_85_n463.t32 19.8
R202 a_85_n463.n259 a_85_n463.t19 19.8
R203 a_85_n463.t0 a_85_n463.n465 19.8
R204 a_85_n463.n465 a_85_n463.t7 19.8
R205 a_85_n463.n442 a_85_n463.n441 8.5
R206 a_85_n463.n427 a_85_n463.n426 8.5
R207 a_85_n463.n412 a_85_n463.n411 8.5
R208 a_85_n463.n397 a_85_n463.n396 8.5
R209 a_85_n463.n382 a_85_n463.n381 8.5
R210 a_85_n463.n367 a_85_n463.n366 8.5
R211 a_85_n463.n352 a_85_n463.n351 8.5
R212 a_85_n463.n337 a_85_n463.n336 8.5
R213 a_85_n463.n322 a_85_n463.n321 8.5
R214 a_85_n463.n307 a_85_n463.n306 8.5
R215 a_85_n463.n292 a_85_n463.n291 8.5
R216 a_85_n463.n277 a_85_n463.n276 8.5
R217 a_85_n463.n230 a_85_n463.n229 8.5
R218 a_85_n463.n245 a_85_n463.n244 8.5
R219 a_85_n463.n260 a_85_n463.n259 8.5
R220 a_85_n463.n21 a_85_n463.n20 8.5
R221 a_85_n463.n34 a_85_n463.n33 8.5
R222 a_85_n463.n47 a_85_n463.n46 8.5
R223 a_85_n463.n60 a_85_n463.n59 8.5
R224 a_85_n463.n73 a_85_n463.n72 8.5
R225 a_85_n463.n86 a_85_n463.n85 8.5
R226 a_85_n463.n99 a_85_n463.n98 8.5
R227 a_85_n463.n112 a_85_n463.n111 8.5
R228 a_85_n463.n125 a_85_n463.n124 8.5
R229 a_85_n463.n138 a_85_n463.n137 8.5
R230 a_85_n463.n151 a_85_n463.n150 8.5
R231 a_85_n463.n164 a_85_n463.n163 8.5
R232 a_85_n463.n177 a_85_n463.n176 8.5
R233 a_85_n463.n465 a_85_n463.n215 8.5
R234 a_85_n463.n465 a_85_n463.n464 8.499
R235 a_85_n463.n25 a_85_n463.n24 7.529
R236 a_85_n463.n38 a_85_n463.n37 7.529
R237 a_85_n463.n51 a_85_n463.n50 7.529
R238 a_85_n463.n64 a_85_n463.n63 7.529
R239 a_85_n463.n77 a_85_n463.n76 7.529
R240 a_85_n463.n90 a_85_n463.n89 7.529
R241 a_85_n463.n103 a_85_n463.n102 7.529
R242 a_85_n463.n116 a_85_n463.n115 7.529
R243 a_85_n463.n129 a_85_n463.n128 7.529
R244 a_85_n463.n142 a_85_n463.n141 7.529
R245 a_85_n463.n155 a_85_n463.n154 7.529
R246 a_85_n463.n168 a_85_n463.n167 7.529
R247 a_85_n463.n181 a_85_n463.n180 7.529
R248 a_85_n463.n437 a_85_n463.n436 7.529
R249 a_85_n463.n422 a_85_n463.n421 7.529
R250 a_85_n463.n407 a_85_n463.n406 7.529
R251 a_85_n463.n392 a_85_n463.n391 7.529
R252 a_85_n463.n377 a_85_n463.n376 7.529
R253 a_85_n463.n362 a_85_n463.n361 7.529
R254 a_85_n463.n347 a_85_n463.n346 7.529
R255 a_85_n463.n332 a_85_n463.n331 7.529
R256 a_85_n463.n317 a_85_n463.n316 7.529
R257 a_85_n463.n302 a_85_n463.n301 7.529
R258 a_85_n463.n287 a_85_n463.n286 7.529
R259 a_85_n463.n272 a_85_n463.n271 7.529
R260 a_85_n463.n225 a_85_n463.n224 7.529
R261 a_85_n463.n240 a_85_n463.n239 7.529
R262 a_85_n463.n255 a_85_n463.n254 7.529
R263 a_85_n463.n462 a_85_n463.n461 7.529
R264 a_85_n463.n434 a_85_n463.n433 4.543
R265 a_85_n463.n419 a_85_n463.n418 4.543
R266 a_85_n463.n404 a_85_n463.n403 4.543
R267 a_85_n463.n389 a_85_n463.n388 4.543
R268 a_85_n463.n374 a_85_n463.n373 4.543
R269 a_85_n463.n359 a_85_n463.n358 4.543
R270 a_85_n463.n344 a_85_n463.n343 4.543
R271 a_85_n463.n329 a_85_n463.n328 4.543
R272 a_85_n463.n314 a_85_n463.n313 4.543
R273 a_85_n463.n299 a_85_n463.n298 4.543
R274 a_85_n463.n284 a_85_n463.n283 4.543
R275 a_85_n463.n269 a_85_n463.n268 4.543
R276 a_85_n463.n222 a_85_n463.n221 4.543
R277 a_85_n463.n237 a_85_n463.n236 4.543
R278 a_85_n463.n252 a_85_n463.n251 4.543
R279 a_85_n463.n463 a_85_n463.n218 4.517
R280 a_85_n463.n12 a_85_n463.n19 4.5
R281 a_85_n463.n12 a_85_n463.n25 4.5
R282 a_85_n463.n12 a_85_n463.n15 4.5
R283 a_85_n463.n11 a_85_n463.n32 4.5
R284 a_85_n463.n11 a_85_n463.n38 4.5
R285 a_85_n463.n11 a_85_n463.n28 4.5
R286 a_85_n463.n10 a_85_n463.n45 4.5
R287 a_85_n463.n10 a_85_n463.n51 4.5
R288 a_85_n463.n10 a_85_n463.n41 4.5
R289 a_85_n463.n9 a_85_n463.n58 4.5
R290 a_85_n463.n9 a_85_n463.n64 4.5
R291 a_85_n463.n9 a_85_n463.n54 4.5
R292 a_85_n463.n8 a_85_n463.n71 4.5
R293 a_85_n463.n8 a_85_n463.n77 4.5
R294 a_85_n463.n8 a_85_n463.n67 4.5
R295 a_85_n463.n7 a_85_n463.n84 4.5
R296 a_85_n463.n7 a_85_n463.n90 4.5
R297 a_85_n463.n7 a_85_n463.n80 4.5
R298 a_85_n463.n6 a_85_n463.n97 4.5
R299 a_85_n463.n6 a_85_n463.n103 4.5
R300 a_85_n463.n6 a_85_n463.n93 4.5
R301 a_85_n463.n5 a_85_n463.n110 4.5
R302 a_85_n463.n5 a_85_n463.n116 4.5
R303 a_85_n463.n5 a_85_n463.n106 4.5
R304 a_85_n463.n4 a_85_n463.n123 4.5
R305 a_85_n463.n4 a_85_n463.n129 4.5
R306 a_85_n463.n4 a_85_n463.n119 4.5
R307 a_85_n463.n3 a_85_n463.n136 4.5
R308 a_85_n463.n3 a_85_n463.n142 4.5
R309 a_85_n463.n3 a_85_n463.n132 4.5
R310 a_85_n463.n2 a_85_n463.n149 4.5
R311 a_85_n463.n2 a_85_n463.n155 4.5
R312 a_85_n463.n2 a_85_n463.n145 4.5
R313 a_85_n463.n1 a_85_n463.n162 4.5
R314 a_85_n463.n1 a_85_n463.n168 4.5
R315 a_85_n463.n1 a_85_n463.n158 4.5
R316 a_85_n463.n0 a_85_n463.n175 4.5
R317 a_85_n463.n0 a_85_n463.n181 4.5
R318 a_85_n463.n0 a_85_n463.n171 4.5
R319 a_85_n463.n183 a_85_n463.n443 4.5
R320 a_85_n463.n182 a_85_n463.n440 4.5
R321 a_85_n463.n434 a_85_n463.n437 4.5
R322 a_85_n463.n185 a_85_n463.n428 4.5
R323 a_85_n463.n184 a_85_n463.n425 4.5
R324 a_85_n463.n419 a_85_n463.n422 4.5
R325 a_85_n463.n187 a_85_n463.n413 4.5
R326 a_85_n463.n186 a_85_n463.n410 4.5
R327 a_85_n463.n404 a_85_n463.n407 4.5
R328 a_85_n463.n189 a_85_n463.n398 4.5
R329 a_85_n463.n188 a_85_n463.n395 4.5
R330 a_85_n463.n389 a_85_n463.n392 4.5
R331 a_85_n463.n191 a_85_n463.n383 4.5
R332 a_85_n463.n190 a_85_n463.n380 4.5
R333 a_85_n463.n374 a_85_n463.n377 4.5
R334 a_85_n463.n193 a_85_n463.n368 4.5
R335 a_85_n463.n192 a_85_n463.n365 4.5
R336 a_85_n463.n359 a_85_n463.n362 4.5
R337 a_85_n463.n195 a_85_n463.n353 4.5
R338 a_85_n463.n194 a_85_n463.n350 4.5
R339 a_85_n463.n344 a_85_n463.n347 4.5
R340 a_85_n463.n197 a_85_n463.n338 4.5
R341 a_85_n463.n196 a_85_n463.n335 4.5
R342 a_85_n463.n329 a_85_n463.n332 4.5
R343 a_85_n463.n199 a_85_n463.n323 4.5
R344 a_85_n463.n198 a_85_n463.n320 4.5
R345 a_85_n463.n314 a_85_n463.n317 4.5
R346 a_85_n463.n201 a_85_n463.n308 4.5
R347 a_85_n463.n200 a_85_n463.n305 4.5
R348 a_85_n463.n299 a_85_n463.n302 4.5
R349 a_85_n463.n203 a_85_n463.n293 4.5
R350 a_85_n463.n202 a_85_n463.n290 4.5
R351 a_85_n463.n284 a_85_n463.n287 4.5
R352 a_85_n463.n205 a_85_n463.n278 4.5
R353 a_85_n463.n204 a_85_n463.n275 4.5
R354 a_85_n463.n269 a_85_n463.n272 4.5
R355 a_85_n463.n207 a_85_n463.n231 4.5
R356 a_85_n463.n206 a_85_n463.n228 4.5
R357 a_85_n463.n222 a_85_n463.n225 4.5
R358 a_85_n463.n209 a_85_n463.n246 4.5
R359 a_85_n463.n208 a_85_n463.n243 4.5
R360 a_85_n463.n237 a_85_n463.n240 4.5
R361 a_85_n463.n211 a_85_n463.n261 4.5
R362 a_85_n463.n210 a_85_n463.n258 4.5
R363 a_85_n463.n252 a_85_n463.n255 4.5
R364 a_85_n463.n460 a_85_n463.n462 4.5
R365 a_85_n463.n19 a_85_n463.n18 3.764
R366 a_85_n463.n32 a_85_n463.n31 3.764
R367 a_85_n463.n45 a_85_n463.n44 3.764
R368 a_85_n463.n58 a_85_n463.n57 3.764
R369 a_85_n463.n71 a_85_n463.n70 3.764
R370 a_85_n463.n84 a_85_n463.n83 3.764
R371 a_85_n463.n97 a_85_n463.n96 3.764
R372 a_85_n463.n110 a_85_n463.n109 3.764
R373 a_85_n463.n123 a_85_n463.n122 3.764
R374 a_85_n463.n136 a_85_n463.n135 3.764
R375 a_85_n463.n149 a_85_n463.n148 3.764
R376 a_85_n463.n162 a_85_n463.n161 3.764
R377 a_85_n463.n175 a_85_n463.n174 3.764
R378 a_85_n463.n440 a_85_n463.n439 3.764
R379 a_85_n463.n425 a_85_n463.n424 3.764
R380 a_85_n463.n410 a_85_n463.n409 3.764
R381 a_85_n463.n395 a_85_n463.n394 3.764
R382 a_85_n463.n380 a_85_n463.n379 3.764
R383 a_85_n463.n365 a_85_n463.n364 3.764
R384 a_85_n463.n350 a_85_n463.n349 3.764
R385 a_85_n463.n335 a_85_n463.n334 3.764
R386 a_85_n463.n320 a_85_n463.n319 3.764
R387 a_85_n463.n305 a_85_n463.n304 3.764
R388 a_85_n463.n290 a_85_n463.n289 3.764
R389 a_85_n463.n275 a_85_n463.n274 3.764
R390 a_85_n463.n228 a_85_n463.n227 3.764
R391 a_85_n463.n243 a_85_n463.n242 3.764
R392 a_85_n463.n258 a_85_n463.n257 3.764
R393 a_85_n463.n217 a_85_n463.n216 3.764
R394 a_85_n463.n15 a_85_n463.n13 3.388
R395 a_85_n463.n28 a_85_n463.n26 3.388
R396 a_85_n463.n41 a_85_n463.n39 3.388
R397 a_85_n463.n54 a_85_n463.n52 3.388
R398 a_85_n463.n67 a_85_n463.n65 3.388
R399 a_85_n463.n80 a_85_n463.n78 3.388
R400 a_85_n463.n93 a_85_n463.n91 3.388
R401 a_85_n463.n106 a_85_n463.n104 3.388
R402 a_85_n463.n119 a_85_n463.n117 3.388
R403 a_85_n463.n132 a_85_n463.n130 3.388
R404 a_85_n463.n145 a_85_n463.n143 3.388
R405 a_85_n463.n158 a_85_n463.n156 3.388
R406 a_85_n463.n171 a_85_n463.n169 3.388
R407 a_85_n463.n433 a_85_n463.n431 3.388
R408 a_85_n463.n418 a_85_n463.n416 3.388
R409 a_85_n463.n403 a_85_n463.n401 3.388
R410 a_85_n463.n388 a_85_n463.n386 3.388
R411 a_85_n463.n373 a_85_n463.n371 3.388
R412 a_85_n463.n358 a_85_n463.n356 3.388
R413 a_85_n463.n343 a_85_n463.n341 3.388
R414 a_85_n463.n328 a_85_n463.n326 3.388
R415 a_85_n463.n313 a_85_n463.n311 3.388
R416 a_85_n463.n298 a_85_n463.n296 3.388
R417 a_85_n463.n283 a_85_n463.n281 3.388
R418 a_85_n463.n268 a_85_n463.n266 3.388
R419 a_85_n463.n221 a_85_n463.n219 3.388
R420 a_85_n463.n236 a_85_n463.n234 3.388
R421 a_85_n463.n251 a_85_n463.n249 3.388
R422 a_85_n463.n215 a_85_n463.n214 3.388
R423 a_85_n463.n15 a_85_n463.n14 3.011
R424 a_85_n463.n25 a_85_n463.n23 3.011
R425 a_85_n463.n28 a_85_n463.n27 3.011
R426 a_85_n463.n38 a_85_n463.n36 3.011
R427 a_85_n463.n41 a_85_n463.n40 3.011
R428 a_85_n463.n51 a_85_n463.n49 3.011
R429 a_85_n463.n54 a_85_n463.n53 3.011
R430 a_85_n463.n64 a_85_n463.n62 3.011
R431 a_85_n463.n67 a_85_n463.n66 3.011
R432 a_85_n463.n77 a_85_n463.n75 3.011
R433 a_85_n463.n80 a_85_n463.n79 3.011
R434 a_85_n463.n90 a_85_n463.n88 3.011
R435 a_85_n463.n93 a_85_n463.n92 3.011
R436 a_85_n463.n103 a_85_n463.n101 3.011
R437 a_85_n463.n106 a_85_n463.n105 3.011
R438 a_85_n463.n116 a_85_n463.n114 3.011
R439 a_85_n463.n119 a_85_n463.n118 3.011
R440 a_85_n463.n129 a_85_n463.n127 3.011
R441 a_85_n463.n132 a_85_n463.n131 3.011
R442 a_85_n463.n142 a_85_n463.n140 3.011
R443 a_85_n463.n145 a_85_n463.n144 3.011
R444 a_85_n463.n155 a_85_n463.n153 3.011
R445 a_85_n463.n158 a_85_n463.n157 3.011
R446 a_85_n463.n168 a_85_n463.n166 3.011
R447 a_85_n463.n171 a_85_n463.n170 3.011
R448 a_85_n463.n181 a_85_n463.n179 3.011
R449 a_85_n463.n433 a_85_n463.n432 3.011
R450 a_85_n463.n437 a_85_n463.n435 3.011
R451 a_85_n463.n418 a_85_n463.n417 3.011
R452 a_85_n463.n422 a_85_n463.n420 3.011
R453 a_85_n463.n403 a_85_n463.n402 3.011
R454 a_85_n463.n407 a_85_n463.n405 3.011
R455 a_85_n463.n388 a_85_n463.n387 3.011
R456 a_85_n463.n392 a_85_n463.n390 3.011
R457 a_85_n463.n373 a_85_n463.n372 3.011
R458 a_85_n463.n377 a_85_n463.n375 3.011
R459 a_85_n463.n358 a_85_n463.n357 3.011
R460 a_85_n463.n362 a_85_n463.n360 3.011
R461 a_85_n463.n343 a_85_n463.n342 3.011
R462 a_85_n463.n347 a_85_n463.n345 3.011
R463 a_85_n463.n328 a_85_n463.n327 3.011
R464 a_85_n463.n332 a_85_n463.n330 3.011
R465 a_85_n463.n313 a_85_n463.n312 3.011
R466 a_85_n463.n317 a_85_n463.n315 3.011
R467 a_85_n463.n298 a_85_n463.n297 3.011
R468 a_85_n463.n302 a_85_n463.n300 3.011
R469 a_85_n463.n283 a_85_n463.n282 3.011
R470 a_85_n463.n287 a_85_n463.n285 3.011
R471 a_85_n463.n268 a_85_n463.n267 3.011
R472 a_85_n463.n272 a_85_n463.n270 3.011
R473 a_85_n463.n221 a_85_n463.n220 3.011
R474 a_85_n463.n225 a_85_n463.n223 3.011
R475 a_85_n463.n236 a_85_n463.n235 3.011
R476 a_85_n463.n240 a_85_n463.n238 3.011
R477 a_85_n463.n251 a_85_n463.n250 3.011
R478 a_85_n463.n255 a_85_n463.n253 3.011
R479 a_85_n463.n214 a_85_n463.n213 3.011
R480 a_85_n463.n213 a_85_n463.n212 2.635
R481 a_85_n463.n22 a_85_n463.n21 1.505
R482 a_85_n463.n35 a_85_n463.n34 1.505
R483 a_85_n463.n48 a_85_n463.n47 1.505
R484 a_85_n463.n61 a_85_n463.n60 1.505
R485 a_85_n463.n74 a_85_n463.n73 1.505
R486 a_85_n463.n87 a_85_n463.n86 1.505
R487 a_85_n463.n100 a_85_n463.n99 1.505
R488 a_85_n463.n113 a_85_n463.n112 1.505
R489 a_85_n463.n126 a_85_n463.n125 1.505
R490 a_85_n463.n139 a_85_n463.n138 1.505
R491 a_85_n463.n152 a_85_n463.n151 1.505
R492 a_85_n463.n165 a_85_n463.n164 1.505
R493 a_85_n463.n178 a_85_n463.n177 1.505
R494 a_85_n463.n443 a_85_n463.n442 1.505
R495 a_85_n463.n428 a_85_n463.n427 1.505
R496 a_85_n463.n413 a_85_n463.n412 1.505
R497 a_85_n463.n398 a_85_n463.n397 1.505
R498 a_85_n463.n383 a_85_n463.n382 1.505
R499 a_85_n463.n368 a_85_n463.n367 1.505
R500 a_85_n463.n353 a_85_n463.n352 1.505
R501 a_85_n463.n338 a_85_n463.n337 1.505
R502 a_85_n463.n323 a_85_n463.n322 1.505
R503 a_85_n463.n308 a_85_n463.n307 1.505
R504 a_85_n463.n293 a_85_n463.n292 1.505
R505 a_85_n463.n278 a_85_n463.n277 1.505
R506 a_85_n463.n231 a_85_n463.n230 1.505
R507 a_85_n463.n246 a_85_n463.n245 1.505
R508 a_85_n463.n261 a_85_n463.n260 1.505
R509 a_85_n463.n464 a_85_n463.n463 1.505
R510 a_85_n463.n460 a_85_n463.n459 1.131
R511 a_85_n463.n444 a_85_n463.n183 0.955
R512 a_85_n463.n429 a_85_n463.n185 0.955
R513 a_85_n463.n414 a_85_n463.n187 0.955
R514 a_85_n463.n399 a_85_n463.n189 0.955
R515 a_85_n463.n384 a_85_n463.n191 0.955
R516 a_85_n463.n369 a_85_n463.n193 0.955
R517 a_85_n463.n354 a_85_n463.n195 0.955
R518 a_85_n463.n339 a_85_n463.n197 0.955
R519 a_85_n463.n324 a_85_n463.n199 0.955
R520 a_85_n463.n309 a_85_n463.n201 0.955
R521 a_85_n463.n294 a_85_n463.n203 0.955
R522 a_85_n463.n279 a_85_n463.n205 0.955
R523 a_85_n463.n232 a_85_n463.n207 0.955
R524 a_85_n463.n247 a_85_n463.n209 0.955
R525 a_85_n463.n262 a_85_n463.n211 0.955
R526 a_85_n463.n172 a_85_n463.n445 0.656
R527 a_85_n463.n16 a_85_n463.n263 0.656
R528 a_85_n463.n446 a_85_n463.n430 0.523
R529 a_85_n463.n447 a_85_n463.n415 0.523
R530 a_85_n463.n448 a_85_n463.n400 0.523
R531 a_85_n463.n449 a_85_n463.n385 0.523
R532 a_85_n463.n450 a_85_n463.n370 0.523
R533 a_85_n463.n451 a_85_n463.n355 0.523
R534 a_85_n463.n452 a_85_n463.n340 0.523
R535 a_85_n463.n453 a_85_n463.n325 0.523
R536 a_85_n463.n454 a_85_n463.n310 0.523
R537 a_85_n463.n455 a_85_n463.n295 0.523
R538 a_85_n463.n456 a_85_n463.n280 0.523
R539 a_85_n463.n265 a_85_n463.n233 0.523
R540 a_85_n463.n264 a_85_n463.n248 0.523
R541 a_85_n463.n458 a_85_n463.n457 0.379
R542 a_85_n463.n18 a_85_n463.n17 0.376
R543 a_85_n463.n31 a_85_n463.n30 0.376
R544 a_85_n463.n44 a_85_n463.n43 0.376
R545 a_85_n463.n57 a_85_n463.n56 0.376
R546 a_85_n463.n70 a_85_n463.n69 0.376
R547 a_85_n463.n83 a_85_n463.n82 0.376
R548 a_85_n463.n96 a_85_n463.n95 0.376
R549 a_85_n463.n109 a_85_n463.n108 0.376
R550 a_85_n463.n122 a_85_n463.n121 0.376
R551 a_85_n463.n135 a_85_n463.n134 0.376
R552 a_85_n463.n148 a_85_n463.n147 0.376
R553 a_85_n463.n161 a_85_n463.n160 0.376
R554 a_85_n463.n174 a_85_n463.n173 0.376
R555 a_85_n463.n439 a_85_n463.n438 0.376
R556 a_85_n463.n424 a_85_n463.n423 0.376
R557 a_85_n463.n409 a_85_n463.n408 0.376
R558 a_85_n463.n394 a_85_n463.n393 0.376
R559 a_85_n463.n379 a_85_n463.n378 0.376
R560 a_85_n463.n364 a_85_n463.n363 0.376
R561 a_85_n463.n349 a_85_n463.n348 0.376
R562 a_85_n463.n334 a_85_n463.n333 0.376
R563 a_85_n463.n319 a_85_n463.n318 0.376
R564 a_85_n463.n304 a_85_n463.n303 0.376
R565 a_85_n463.n289 a_85_n463.n288 0.376
R566 a_85_n463.n274 a_85_n463.n273 0.376
R567 a_85_n463.n227 a_85_n463.n226 0.376
R568 a_85_n463.n242 a_85_n463.n241 0.376
R569 a_85_n463.n257 a_85_n463.n256 0.376
R570 a_85_n463.n218 a_85_n463.n217 0.376
R571 a_85_n463.n264 a_85_n463.n16 0.133
R572 a_85_n463.n29 a_85_n463.n264 0.133
R573 a_85_n463.n265 a_85_n463.n29 0.133
R574 a_85_n463.n457 a_85_n463.n265 0.133
R575 a_85_n463.n457 a_85_n463.n456 0.133
R576 a_85_n463.n456 a_85_n463.n42 0.133
R577 a_85_n463.n42 a_85_n463.n455 0.133
R578 a_85_n463.n455 a_85_n463.n55 0.133
R579 a_85_n463.n55 a_85_n463.n454 0.133
R580 a_85_n463.n454 a_85_n463.n68 0.133
R581 a_85_n463.n68 a_85_n463.n453 0.133
R582 a_85_n463.n453 a_85_n463.n81 0.133
R583 a_85_n463.n81 a_85_n463.n452 0.133
R584 a_85_n463.n452 a_85_n463.n94 0.133
R585 a_85_n463.n94 a_85_n463.n451 0.133
R586 a_85_n463.n451 a_85_n463.n107 0.133
R587 a_85_n463.n107 a_85_n463.n450 0.133
R588 a_85_n463.n450 a_85_n463.n120 0.133
R589 a_85_n463.n120 a_85_n463.n449 0.133
R590 a_85_n463.n449 a_85_n463.n133 0.133
R591 a_85_n463.n133 a_85_n463.n448 0.133
R592 a_85_n463.n448 a_85_n463.n146 0.133
R593 a_85_n463.n146 a_85_n463.n447 0.133
R594 a_85_n463.n447 a_85_n463.n159 0.133
R595 a_85_n463.n159 a_85_n463.n446 0.133
R596 a_85_n463.n446 a_85_n463.n172 0.133
R597 a_85_n463.n463 a_85_n463.n460 4.63
R598 a_85_n463.n182 a_85_n463.n434 0.087
R599 a_85_n463.n184 a_85_n463.n419 0.087
R600 a_85_n463.n186 a_85_n463.n404 0.087
R601 a_85_n463.n188 a_85_n463.n389 0.087
R602 a_85_n463.n190 a_85_n463.n374 0.087
R603 a_85_n463.n192 a_85_n463.n359 0.087
R604 a_85_n463.n194 a_85_n463.n344 0.087
R605 a_85_n463.n196 a_85_n463.n329 0.087
R606 a_85_n463.n198 a_85_n463.n314 0.087
R607 a_85_n463.n200 a_85_n463.n299 0.087
R608 a_85_n463.n202 a_85_n463.n284 0.087
R609 a_85_n463.n204 a_85_n463.n269 0.087
R610 a_85_n463.n206 a_85_n463.n222 0.087
R611 a_85_n463.n208 a_85_n463.n237 0.087
R612 a_85_n463.n210 a_85_n463.n252 0.087
R613 a_85_n463.n211 a_85_n463.n210 0.046
R614 a_85_n463.n209 a_85_n463.n208 0.046
R615 a_85_n463.n207 a_85_n463.n206 0.046
R616 a_85_n463.n205 a_85_n463.n204 0.046
R617 a_85_n463.n203 a_85_n463.n202 0.046
R618 a_85_n463.n201 a_85_n463.n200 0.046
R619 a_85_n463.n199 a_85_n463.n198 0.046
R620 a_85_n463.n197 a_85_n463.n196 0.046
R621 a_85_n463.n195 a_85_n463.n194 0.046
R622 a_85_n463.n193 a_85_n463.n192 0.046
R623 a_85_n463.n191 a_85_n463.n190 0.046
R624 a_85_n463.n189 a_85_n463.n188 0.046
R625 a_85_n463.n187 a_85_n463.n186 0.046
R626 a_85_n463.n185 a_85_n463.n184 0.046
R627 a_85_n463.n183 a_85_n463.n182 0.046
R628 a_85_n463.n459 a_85_n463.n458 0.045
R629 a_85_n463.n445 a_85_n463.n444 0.041
R630 a_85_n463.n430 a_85_n463.n429 0.041
R631 a_85_n463.n415 a_85_n463.n414 0.041
R632 a_85_n463.n400 a_85_n463.n399 0.041
R633 a_85_n463.n385 a_85_n463.n384 0.041
R634 a_85_n463.n370 a_85_n463.n369 0.041
R635 a_85_n463.n355 a_85_n463.n354 0.041
R636 a_85_n463.n340 a_85_n463.n339 0.041
R637 a_85_n463.n325 a_85_n463.n324 0.041
R638 a_85_n463.n310 a_85_n463.n309 0.041
R639 a_85_n463.n295 a_85_n463.n294 0.041
R640 a_85_n463.n280 a_85_n463.n279 0.041
R641 a_85_n463.n233 a_85_n463.n232 0.041
R642 a_85_n463.n248 a_85_n463.n247 0.041
R643 a_85_n463.n263 a_85_n463.n262 0.041
R644 a_85_n463.n0 a_85_n463.n178 4.543
R645 a_85_n463.n1 a_85_n463.n165 4.543
R646 a_85_n463.n2 a_85_n463.n152 4.543
R647 a_85_n463.n3 a_85_n463.n139 4.543
R648 a_85_n463.n4 a_85_n463.n126 4.543
R649 a_85_n463.n5 a_85_n463.n113 4.543
R650 a_85_n463.n6 a_85_n463.n100 4.543
R651 a_85_n463.n7 a_85_n463.n87 4.543
R652 a_85_n463.n8 a_85_n463.n74 4.543
R653 a_85_n463.n9 a_85_n463.n61 4.543
R654 a_85_n463.n10 a_85_n463.n48 4.543
R655 a_85_n463.n11 a_85_n463.n35 4.543
R656 a_85_n463.n12 a_85_n463.n22 4.543
R657 a_85_n463.n0 a_85_n463.n172 1.643
R658 a_85_n463.n12 a_85_n463.n16 1.642
R659 a_85_n463.n11 a_85_n463.n29 1.642
R660 a_85_n463.n10 a_85_n463.n42 1.642
R661 a_85_n463.n9 a_85_n463.n55 1.642
R662 a_85_n463.n8 a_85_n463.n68 1.642
R663 a_85_n463.n7 a_85_n463.n81 1.642
R664 a_85_n463.n6 a_85_n463.n94 1.642
R665 a_85_n463.n5 a_85_n463.n107 1.642
R666 a_85_n463.n4 a_85_n463.n120 1.642
R667 a_85_n463.n3 a_85_n463.n133 1.642
R668 a_85_n463.n2 a_85_n463.n146 1.642
R669 a_85_n463.n1 a_85_n463.n159 1.642
R670 source.n402 source.t4 19.8
R671 source.n402 source.t17 19.8
R672 source.n372 source.t9 19.8
R673 source.n372 source.t27 19.8
R674 source.n342 source.t20 19.8
R675 source.n342 source.t12 19.8
R676 source.n312 source.t0 19.8
R677 source.n312 source.t23 19.8
R678 source.n282 source.t18 19.8
R679 source.n282 source.t11 19.8
R680 source.n252 source.t7 19.8
R681 source.n252 source.t22 19.8
R682 source.n222 source.t14 19.8
R683 source.n222 source.t2 19.8
R684 source.n6 source.t25 19.8
R685 source.n6 source.t16 19.8
R686 source.n36 source.t8 19.8
R687 source.n36 source.t5 19.8
R688 source.n66 source.t19 19.8
R689 source.n66 source.t10 19.8
R690 source.n96 source.t6 19.8
R691 source.n96 source.t21 19.8
R692 source.n126 source.t13 19.8
R693 source.n126 source.t1 19.8
R694 source.n156 source.t24 19.8
R695 source.n156 source.t15 19.8
R696 source.n183 source.t3 19.8
R697 source.n183 source.t26 19.8
R698 source.n403 source.n402 8.5
R699 source.n373 source.n372 8.5
R700 source.n343 source.n342 8.5
R701 source.n313 source.n312 8.5
R702 source.n283 source.n282 8.5
R703 source.n253 source.n252 8.5
R704 source.n223 source.n222 8.5
R705 source.n7 source.n6 8.5
R706 source.n37 source.n36 8.5
R707 source.n67 source.n66 8.5
R708 source.n97 source.n96 8.5
R709 source.n127 source.n126 8.5
R710 source.n157 source.n156 8.5
R711 source.n184 source.n183 8.5
R712 source.n414 source.n413 7.529
R713 source.n384 source.n383 7.529
R714 source.n354 source.n353 7.529
R715 source.n324 source.n323 7.529
R716 source.n294 source.n293 7.529
R717 source.n264 source.n263 7.529
R718 source.n234 source.n233 7.529
R719 source.n18 source.n17 7.529
R720 source.n48 source.n47 7.529
R721 source.n78 source.n77 7.529
R722 source.n108 source.n107 7.529
R723 source.n138 source.n137 7.529
R724 source.n168 source.n167 7.529
R725 source.n195 source.n194 7.529
R726 source.n409 source.n401 4.5
R727 source.n406 source.n404 4.5
R728 source.n415 source.n414 4.5
R729 source.n418 source.n398 4.5
R730 source.n379 source.n371 4.5
R731 source.n376 source.n374 4.5
R732 source.n385 source.n384 4.5
R733 source.n388 source.n368 4.5
R734 source.n349 source.n341 4.5
R735 source.n346 source.n344 4.5
R736 source.n355 source.n354 4.5
R737 source.n358 source.n338 4.5
R738 source.n319 source.n311 4.5
R739 source.n316 source.n314 4.5
R740 source.n325 source.n324 4.5
R741 source.n328 source.n308 4.5
R742 source.n289 source.n281 4.5
R743 source.n286 source.n284 4.5
R744 source.n295 source.n294 4.5
R745 source.n298 source.n278 4.5
R746 source.n259 source.n251 4.5
R747 source.n256 source.n254 4.5
R748 source.n265 source.n264 4.5
R749 source.n268 source.n248 4.5
R750 source.n229 source.n221 4.5
R751 source.n226 source.n224 4.5
R752 source.n235 source.n234 4.5
R753 source.n238 source.n218 4.5
R754 source.n13 source.n5 4.5
R755 source.n10 source.n8 4.5
R756 source.n19 source.n18 4.5
R757 source.n22 source.n2 4.5
R758 source.n43 source.n35 4.5
R759 source.n40 source.n38 4.5
R760 source.n49 source.n48 4.5
R761 source.n52 source.n32 4.5
R762 source.n73 source.n65 4.5
R763 source.n70 source.n68 4.5
R764 source.n79 source.n78 4.5
R765 source.n82 source.n62 4.5
R766 source.n103 source.n95 4.5
R767 source.n100 source.n98 4.5
R768 source.n109 source.n108 4.5
R769 source.n112 source.n92 4.5
R770 source.n133 source.n125 4.5
R771 source.n130 source.n128 4.5
R772 source.n139 source.n138 4.5
R773 source.n142 source.n122 4.5
R774 source.n163 source.n155 4.5
R775 source.n160 source.n158 4.5
R776 source.n169 source.n168 4.5
R777 source.n172 source.n152 4.5
R778 source.n187 source.n185 4.5
R779 source.n190 source.n182 4.5
R780 source.n196 source.n195 4.5
R781 source.n202 source.n201 4.5
R782 source.n401 source.n400 3.764
R783 source.n371 source.n370 3.764
R784 source.n341 source.n340 3.764
R785 source.n311 source.n310 3.764
R786 source.n281 source.n280 3.764
R787 source.n251 source.n250 3.764
R788 source.n221 source.n220 3.764
R789 source.n5 source.n4 3.764
R790 source.n35 source.n34 3.764
R791 source.n65 source.n64 3.764
R792 source.n95 source.n94 3.764
R793 source.n125 source.n124 3.764
R794 source.n155 source.n154 3.764
R795 source.n182 source.n181 3.764
R796 source.n398 source.n396 3.388
R797 source.n368 source.n366 3.388
R798 source.n338 source.n336 3.388
R799 source.n308 source.n306 3.388
R800 source.n278 source.n276 3.388
R801 source.n248 source.n246 3.388
R802 source.n218 source.n216 3.388
R803 source.n2 source.n0 3.388
R804 source.n32 source.n30 3.388
R805 source.n62 source.n60 3.388
R806 source.n92 source.n90 3.388
R807 source.n122 source.n120 3.388
R808 source.n152 source.n150 3.388
R809 source.n201 source.n199 3.388
R810 source.n398 source.n397 3.011
R811 source.n414 source.n412 3.011
R812 source.n368 source.n367 3.011
R813 source.n384 source.n382 3.011
R814 source.n338 source.n337 3.011
R815 source.n354 source.n352 3.011
R816 source.n308 source.n307 3.011
R817 source.n324 source.n322 3.011
R818 source.n278 source.n277 3.011
R819 source.n294 source.n292 3.011
R820 source.n248 source.n247 3.011
R821 source.n264 source.n262 3.011
R822 source.n218 source.n217 3.011
R823 source.n234 source.n232 3.011
R824 source.n2 source.n1 3.011
R825 source.n18 source.n16 3.011
R826 source.n32 source.n31 3.011
R827 source.n48 source.n46 3.011
R828 source.n62 source.n61 3.011
R829 source.n78 source.n76 3.011
R830 source.n92 source.n91 3.011
R831 source.n108 source.n106 3.011
R832 source.n122 source.n121 3.011
R833 source.n138 source.n136 3.011
R834 source.n152 source.n151 3.011
R835 source.n168 source.n166 3.011
R836 source.n201 source.n200 3.011
R837 source.n195 source.n193 3.011
R838 source.n404 source.n403 1.505
R839 source.n374 source.n373 1.505
R840 source.n344 source.n343 1.505
R841 source.n314 source.n313 1.505
R842 source.n284 source.n283 1.505
R843 source.n254 source.n253 1.505
R844 source.n224 source.n223 1.505
R845 source.n8 source.n7 1.505
R846 source.n38 source.n37 1.505
R847 source.n68 source.n67 1.505
R848 source.n98 source.n97 1.505
R849 source.n128 source.n127 1.505
R850 source.n158 source.n157 1.505
R851 source.n185 source.n184 1.505
R852 source.n204 source.n203 0.95
R853 source.n420 source.n419 0.949
R854 source.n390 source.n389 0.949
R855 source.n360 source.n359 0.949
R856 source.n330 source.n329 0.949
R857 source.n300 source.n299 0.949
R858 source.n270 source.n269 0.949
R859 source.n240 source.n239 0.949
R860 source.n24 source.n23 0.949
R861 source.n54 source.n53 0.949
R862 source.n84 source.n83 0.949
R863 source.n114 source.n113 0.949
R864 source.n144 source.n143 0.949
R865 source.n174 source.n173 0.949
R866 source.n426 source.n425 0.399
R867 source.n210 source.n209 0.399
R868 source.n400 source.n399 0.376
R869 source.n370 source.n369 0.376
R870 source.n340 source.n339 0.376
R871 source.n310 source.n309 0.376
R872 source.n280 source.n279 0.376
R873 source.n250 source.n249 0.376
R874 source.n220 source.n219 0.376
R875 source.n4 source.n3 0.376
R876 source.n34 source.n33 0.376
R877 source.n64 source.n63 0.376
R878 source.n94 source.n93 0.376
R879 source.n124 source.n123 0.376
R880 source.n154 source.n153 0.376
R881 source.n181 source.n180 0.376
R882 source.n426 source.n395 0.369
R883 source.n427 source.n365 0.369
R884 source.n428 source.n335 0.369
R885 source.n429 source.n305 0.369
R886 source.n430 source.n275 0.369
R887 source.n431 source.n245 0.369
R888 source.n215 source.n29 0.369
R889 source.n214 source.n59 0.369
R890 source.n213 source.n89 0.369
R891 source.n212 source.n119 0.369
R892 source.n211 source.n149 0.369
R893 source.n210 source.n179 0.369
R894 source.n425 source.n424 0.045
R895 source.n395 source.n394 0.045
R896 source.n365 source.n364 0.045
R897 source.n335 source.n334 0.045
R898 source.n305 source.n304 0.045
R899 source.n275 source.n274 0.045
R900 source.n245 source.n244 0.045
R901 source.n29 source.n28 0.045
R902 source.n59 source.n58 0.045
R903 source.n89 source.n88 0.045
R904 source.n119 source.n118 0.045
R905 source.n149 source.n148 0.045
R906 source.n179 source.n178 0.045
R907 source.n209 source.n208 0.045
R908 source.n424 source.n423 0.044
R909 source.n394 source.n393 0.044
R910 source.n364 source.n363 0.044
R911 source.n334 source.n333 0.044
R912 source.n304 source.n303 0.044
R913 source.n274 source.n273 0.044
R914 source.n244 source.n243 0.044
R915 source.n28 source.n27 0.044
R916 source.n58 source.n57 0.044
R917 source.n88 source.n87 0.044
R918 source.n118 source.n117 0.044
R919 source.n148 source.n147 0.044
R920 source.n178 source.n177 0.044
R921 source.n208 source.n207 0.044
R922 source.n410 source.n409 0.041
R923 source.n423 source.n422 0.041
R924 source.n380 source.n379 0.041
R925 source.n393 source.n392 0.041
R926 source.n350 source.n349 0.041
R927 source.n363 source.n362 0.041
R928 source.n320 source.n319 0.041
R929 source.n333 source.n332 0.041
R930 source.n290 source.n289 0.041
R931 source.n303 source.n302 0.041
R932 source.n260 source.n259 0.041
R933 source.n273 source.n272 0.041
R934 source.n230 source.n229 0.041
R935 source.n243 source.n242 0.041
R936 source.n14 source.n13 0.041
R937 source.n27 source.n26 0.041
R938 source.n44 source.n43 0.041
R939 source.n57 source.n56 0.041
R940 source.n74 source.n73 0.041
R941 source.n87 source.n86 0.041
R942 source.n104 source.n103 0.041
R943 source.n117 source.n116 0.041
R944 source.n134 source.n133 0.041
R945 source.n147 source.n146 0.041
R946 source.n164 source.n163 0.041
R947 source.n177 source.n176 0.041
R948 source.n191 source.n190 0.041
R949 source.n207 source.n206 0.041
R950 source.n415 source.n411 0.039
R951 source.n421 source.n420 0.039
R952 source.n385 source.n381 0.039
R953 source.n391 source.n390 0.039
R954 source.n355 source.n351 0.039
R955 source.n361 source.n360 0.039
R956 source.n325 source.n321 0.039
R957 source.n331 source.n330 0.039
R958 source.n295 source.n291 0.039
R959 source.n301 source.n300 0.039
R960 source.n265 source.n261 0.039
R961 source.n271 source.n270 0.039
R962 source.n235 source.n231 0.039
R963 source.n241 source.n240 0.039
R964 source.n19 source.n15 0.039
R965 source.n25 source.n24 0.039
R966 source.n49 source.n45 0.039
R967 source.n55 source.n54 0.039
R968 source.n79 source.n75 0.039
R969 source.n85 source.n84 0.039
R970 source.n109 source.n105 0.039
R971 source.n115 source.n114 0.039
R972 source.n139 source.n135 0.039
R973 source.n145 source.n144 0.039
R974 source.n169 source.n165 0.039
R975 source.n175 source.n174 0.039
R976 source.n196 source.n192 0.039
R977 source.n205 source.n204 0.039
R978 source.n427 source.n426 0.03
R979 source.n428 source.n427 0.03
R980 source.n429 source.n428 0.03
R981 source.n430 source.n429 0.03
R982 source.n431 source.n430 0.03
R983 source.n215 source.n214 0.03
R984 source.n214 source.n213 0.03
R985 source.n213 source.n212 0.03
R986 source.n212 source.n211 0.03
R987 source.n211 source.n210 0.03
R988 source.n407 source.n406 0.023
R989 source.n377 source.n376 0.023
R990 source.n347 source.n346 0.023
R991 source.n317 source.n316 0.023
R992 source.n287 source.n286 0.023
R993 source.n257 source.n256 0.023
R994 source.n227 source.n226 0.023
R995 source.n11 source.n10 0.023
R996 source.n41 source.n40 0.023
R997 source.n71 source.n70 0.023
R998 source.n101 source.n100 0.023
R999 source.n131 source.n130 0.023
R1000 source.n161 source.n160 0.023
R1001 source.n188 source.n187 0.023
R1002 source.n409 source.n408 0.019
R1003 source.n379 source.n378 0.019
R1004 source.n349 source.n348 0.019
R1005 source.n319 source.n318 0.019
R1006 source.n289 source.n288 0.019
R1007 source.n259 source.n258 0.019
R1008 source.n229 source.n228 0.019
R1009 source.n13 source.n12 0.019
R1010 source.n43 source.n42 0.019
R1011 source.n73 source.n72 0.019
R1012 source.n103 source.n102 0.019
R1013 source.n133 source.n132 0.019
R1014 source.n163 source.n162 0.019
R1015 source.n190 source.n189 0.019
R1016 source.n418 source.n417 0.015
R1017 source.n416 source.n415 0.015
R1018 source.n388 source.n387 0.015
R1019 source.n386 source.n385 0.015
R1020 source.n358 source.n357 0.015
R1021 source.n356 source.n355 0.015
R1022 source.n328 source.n327 0.015
R1023 source.n326 source.n325 0.015
R1024 source.n298 source.n297 0.015
R1025 source.n296 source.n295 0.015
R1026 source.n268 source.n267 0.015
R1027 source.n266 source.n265 0.015
R1028 source.n238 source.n237 0.015
R1029 source.n236 source.n235 0.015
R1030 source.n22 source.n21 0.015
R1031 source.n20 source.n19 0.015
R1032 source.n52 source.n51 0.015
R1033 source.n50 source.n49 0.015
R1034 source.n82 source.n81 0.015
R1035 source.n80 source.n79 0.015
R1036 source.n112 source.n111 0.015
R1037 source.n110 source.n109 0.015
R1038 source.n142 source.n141 0.015
R1039 source.n140 source.n139 0.015
R1040 source.n172 source.n171 0.015
R1041 source.n170 source.n169 0.015
R1042 source.n202 source.n198 0.015
R1043 source.n197 source.n196 0.015
R1044 source.n432 source.n215 0.015
R1045 source.n432 source.n431 0.014
R1046 source.n417 source.n416 0.013
R1047 source.n387 source.n386 0.013
R1048 source.n357 source.n356 0.013
R1049 source.n327 source.n326 0.013
R1050 source.n297 source.n296 0.013
R1051 source.n267 source.n266 0.013
R1052 source.n237 source.n236 0.013
R1053 source.n21 source.n20 0.013
R1054 source.n51 source.n50 0.013
R1055 source.n81 source.n80 0.013
R1056 source.n111 source.n110 0.013
R1057 source.n141 source.n140 0.013
R1058 source.n171 source.n170 0.013
R1059 source.n198 source.n197 0.013
R1060 source.n203 source.n202 0.008
R1061 source.n419 source.n418 0.007
R1062 source.n389 source.n388 0.007
R1063 source.n359 source.n358 0.007
R1064 source.n329 source.n328 0.007
R1065 source.n299 source.n298 0.007
R1066 source.n269 source.n268 0.007
R1067 source.n239 source.n238 0.007
R1068 source.n23 source.n22 0.007
R1069 source.n53 source.n52 0.007
R1070 source.n83 source.n82 0.007
R1071 source.n113 source.n112 0.007
R1072 source.n143 source.n142 0.007
R1073 source.n173 source.n172 0.007
R1074 source.n411 source.n410 0.007
R1075 source.n406 source.n405 0.007
R1076 source.n422 source.n421 0.007
R1077 source.n381 source.n380 0.007
R1078 source.n376 source.n375 0.007
R1079 source.n392 source.n391 0.007
R1080 source.n351 source.n350 0.007
R1081 source.n346 source.n345 0.007
R1082 source.n362 source.n361 0.007
R1083 source.n321 source.n320 0.007
R1084 source.n316 source.n315 0.007
R1085 source.n332 source.n331 0.007
R1086 source.n291 source.n290 0.007
R1087 source.n286 source.n285 0.007
R1088 source.n302 source.n301 0.007
R1089 source.n261 source.n260 0.007
R1090 source.n256 source.n255 0.007
R1091 source.n272 source.n271 0.007
R1092 source.n231 source.n230 0.007
R1093 source.n226 source.n225 0.007
R1094 source.n242 source.n241 0.007
R1095 source.n15 source.n14 0.007
R1096 source.n10 source.n9 0.007
R1097 source.n26 source.n25 0.007
R1098 source.n45 source.n44 0.007
R1099 source.n40 source.n39 0.007
R1100 source.n56 source.n55 0.007
R1101 source.n75 source.n74 0.007
R1102 source.n70 source.n69 0.007
R1103 source.n86 source.n85 0.007
R1104 source.n105 source.n104 0.007
R1105 source.n100 source.n99 0.007
R1106 source.n116 source.n115 0.007
R1107 source.n135 source.n134 0.007
R1108 source.n130 source.n129 0.007
R1109 source.n146 source.n145 0.007
R1110 source.n165 source.n164 0.007
R1111 source.n160 source.n159 0.007
R1112 source.n176 source.n175 0.007
R1113 source.n192 source.n191 0.007
R1114 source.n187 source.n186 0.007
R1115 source.n206 source.n205 0.007
R1116 source source.n432 0.002
R1117 source.n408 source.n407 0.001
R1118 source.n378 source.n377 0.001
R1119 source.n348 source.n347 0.001
R1120 source.n318 source.n317 0.001
R1121 source.n288 source.n287 0.001
R1122 source.n258 source.n257 0.001
R1123 source.n228 source.n227 0.001
R1124 source.n12 source.n11 0.001
R1125 source.n42 source.n41 0.001
R1126 source.n72 source.n71 0.001
R1127 source.n102 source.n101 0.001
R1128 source.n132 source.n131 0.001
R1129 source.n162 source.n161 0.001
R1130 source.n189 source.n188 0.001
R1131 bulk.t292 bulk.t1 6442.86
R1132 bulk.t195 bulk.t364 6442.86
R1133 bulk.t273 bulk.t325 6442.86
R1134 bulk.t59 bulk.t347 6442.86
R1135 bulk.t15 bulk.t263 6442.86
R1136 bulk.t161 bulk.t249 6442.86
R1137 bulk.t157 bulk.t190 6442.86
R1138 bulk.t306 bulk.t93 6442.86
R1139 bulk.n66 bulk.t292 2671.43
R1140 bulk.n344 bulk.t273 2671.43
R1141 bulk.n375 bulk.t15 2671.43
R1142 bulk.n41 bulk.t157 2671.43
R1143 bulk.n10 bulk.t195 2584.13
R1144 bulk.n279 bulk.t59 2584.13
R1145 bulk.n521 bulk.t161 2584.13
R1146 bulk.n225 bulk.t306 2584.13
R1147 bulk.t1 bulk.t320 1676.19
R1148 bulk.t320 bulk.t359 1676.19
R1149 bulk.t359 bulk.t2 1676.19
R1150 bulk.t2 bulk.t0 1676.19
R1151 bulk.t0 bulk.t317 1676.19
R1152 bulk.t317 bulk.t314 1676.19
R1153 bulk.t314 bulk.t349 1676.19
R1154 bulk.t349 bulk.t315 1676.19
R1155 bulk.t315 bulk.t356 1676.19
R1156 bulk.t356 bulk.t360 1676.19
R1157 bulk.t360 bulk.t319 1676.19
R1158 bulk.t319 bulk.t351 1676.19
R1159 bulk.t351 bulk.t316 1676.19
R1160 bulk.t350 bulk.t354 1676.19
R1161 bulk.t355 bulk.t350 1676.19
R1162 bulk.t353 bulk.t355 1676.19
R1163 bulk.t352 bulk.t353 1676.19
R1164 bulk.t363 bulk.t352 1676.19
R1165 bulk.t361 bulk.t363 1676.19
R1166 bulk.t365 bulk.t361 1676.19
R1167 bulk.t358 bulk.t365 1676.19
R1168 bulk.t357 bulk.t358 1676.19
R1169 bulk.t3 bulk.t357 1676.19
R1170 bulk.t362 bulk.t3 1676.19
R1171 bulk.t318 bulk.t362 1676.19
R1172 bulk.t364 bulk.t318 1676.19
R1173 bulk.t325 bulk.t338 1676.19
R1174 bulk.t338 bulk.t330 1676.19
R1175 bulk.t330 bulk.t348 1676.19
R1176 bulk.t348 bulk.t341 1676.19
R1177 bulk.t341 bulk.t333 1676.19
R1178 bulk.t333 bulk.t321 1676.19
R1179 bulk.t321 bulk.t344 1676.19
R1180 bulk.t344 bulk.t339 1676.19
R1181 bulk.t339 bulk.t332 1676.19
R1182 bulk.t332 bulk.t328 1676.19
R1183 bulk.t328 bulk.t343 1676.19
R1184 bulk.t343 bulk.t335 1676.19
R1185 bulk.t335 bulk.t323 1676.19
R1186 bulk.t337 bulk.t346 1676.19
R1187 bulk.t329 bulk.t337 1676.19
R1188 bulk.t326 bulk.t329 1676.19
R1189 bulk.t340 bulk.t326 1676.19
R1190 bulk.t331 bulk.t340 1676.19
R1191 bulk.t327 bulk.t331 1676.19
R1192 bulk.t342 bulk.t327 1676.19
R1193 bulk.t334 bulk.t342 1676.19
R1194 bulk.t322 bulk.t334 1676.19
R1195 bulk.t345 bulk.t322 1676.19
R1196 bulk.t336 bulk.t345 1676.19
R1197 bulk.t324 bulk.t336 1676.19
R1198 bulk.t347 bulk.t324 1676.19
R1199 bulk.t263 bulk.t296 1676.19
R1200 bulk.t296 bulk.t24 1676.19
R1201 bulk.t24 bulk.t165 1676.19
R1202 bulk.t165 bulk.t199 1676.19
R1203 bulk.t199 bulk.t268 1676.19
R1204 bulk.t268 bulk.t310 1676.19
R1205 bulk.t310 bulk.t44 1676.19
R1206 bulk.t44 bulk.t142 1676.19
R1207 bulk.t142 bulk.t175 1676.19
R1208 bulk.t175 bulk.t229 1676.19
R1209 bulk.t229 bulk.t287 1676.19
R1210 bulk.t287 bulk.t10 1676.19
R1211 bulk.t10 bulk.t152 1676.19
R1212 bulk.t253 bulk.t185 1676.19
R1213 bulk.t258 bulk.t253 1676.19
R1214 bulk.t277 bulk.t258 1676.19
R1215 bulk.t19 bulk.t277 1676.19
R1216 bulk.t301 bulk.t19 1676.19
R1217 bulk.t34 bulk.t301 1676.19
R1218 bulk.t170 bulk.t34 1676.19
R1219 bulk.t214 bulk.t170 1676.19
R1220 bulk.t282 bulk.t214 1676.19
R1221 bulk.t5 bulk.t282 1676.19
R1222 bulk.t54 bulk.t5 1676.19
R1223 bulk.t180 bulk.t54 1676.19
R1224 bulk.t249 bulk.t180 1676.19
R1225 bulk.t190 bulk.t224 1676.19
R1226 bulk.t224 bulk.t204 1676.19
R1227 bulk.t204 bulk.t239 1676.19
R1228 bulk.t239 bulk.t219 1676.19
R1229 bulk.t219 bulk.t209 1676.19
R1230 bulk.t209 bulk.t244 1676.19
R1231 bulk.t244 bulk.t234 1676.19
R1232 bulk.t234 bulk.t127 1676.19
R1233 bulk.t127 bulk.t112 1676.19
R1234 bulk.t112 bulk.t107 1676.19
R1235 bulk.t107 bulk.t132 1676.19
R1236 bulk.t132 bulk.t117 1676.19
R1237 bulk.t117 bulk.t147 1676.19
R1238 bulk.t122 bulk.t137 1676.19
R1239 bulk.t39 bulk.t122 1676.19
R1240 bulk.t29 bulk.t39 1676.19
R1241 bulk.t49 bulk.t29 1676.19
R1242 bulk.t68 bulk.t49 1676.19
R1243 bulk.t63 bulk.t68 1676.19
R1244 bulk.t83 bulk.t63 1676.19
R1245 bulk.t73 bulk.t83 1676.19
R1246 bulk.t97 bulk.t73 1676.19
R1247 bulk.t88 bulk.t97 1676.19
R1248 bulk.t78 bulk.t88 1676.19
R1249 bulk.t102 bulk.t78 1676.19
R1250 bulk.t93 bulk.t102 1676.19
R1251 bulk.n504 bulk.t248 286.107
R1252 bulk.n496 bulk.t53 286.107
R1253 bulk.n488 bulk.t281 286.107
R1254 bulk.n480 bulk.t169 286.107
R1255 bulk.n472 bulk.t300 286.107
R1256 bulk.n464 bulk.t276 286.107
R1257 bulk.n456 bulk.t252 286.107
R1258 bulk.n448 bulk.t151 286.107
R1259 bulk.n440 bulk.t286 286.107
R1260 bulk.n432 bulk.t174 286.107
R1261 bulk.n424 bulk.t43 286.107
R1262 bulk.n416 bulk.t267 286.107
R1263 bulk.n408 bulk.t164 286.107
R1264 bulk.n400 bulk.t295 286.107
R1265 bulk.n109 bulk.t223 286.107
R1266 bulk.n117 bulk.t238 286.107
R1267 bulk.n125 bulk.t208 286.107
R1268 bulk.n133 bulk.t233 286.107
R1269 bulk.n141 bulk.t111 286.107
R1270 bulk.n149 bulk.t131 286.107
R1271 bulk.n157 bulk.t146 286.107
R1272 bulk.n165 bulk.t121 286.107
R1273 bulk.n173 bulk.t28 286.107
R1274 bulk.n181 bulk.t67 286.107
R1275 bulk.n189 bulk.t82 286.107
R1276 bulk.n197 bulk.t96 286.107
R1277 bulk.n205 bulk.t77 286.107
R1278 bulk.n213 bulk.t92 286.107
R1279 bulk.n532 bulk.t160 233.526
R1280 bulk.n564 bulk.t58 233.526
R1281 bulk.n250 bulk.t194 233.526
R1282 bulk.n219 bulk.t305 233.526
R1283 bulk.n500 bulk.t179 233.526
R1284 bulk.n492 bulk.t4 233.526
R1285 bulk.n484 bulk.t213 233.526
R1286 bulk.n476 bulk.t33 233.526
R1287 bulk.n468 bulk.t18 233.526
R1288 bulk.n460 bulk.t257 233.526
R1289 bulk.n452 bulk.t184 233.526
R1290 bulk.n444 bulk.t9 233.526
R1291 bulk.n436 bulk.t228 233.526
R1292 bulk.n428 bulk.t141 233.526
R1293 bulk.n420 bulk.t309 233.526
R1294 bulk.n412 bulk.t198 233.526
R1295 bulk.n404 bulk.t23 233.526
R1296 bulk.n396 bulk.t262 233.526
R1297 bulk.n34 bulk.t156 233.526
R1298 bulk.n209 bulk.t101 233.526
R1299 bulk.n201 bulk.t87 233.526
R1300 bulk.n193 bulk.t72 233.526
R1301 bulk.n185 bulk.t62 233.526
R1302 bulk.n177 bulk.t48 233.526
R1303 bulk.n169 bulk.t38 233.526
R1304 bulk.n161 bulk.t136 233.526
R1305 bulk.n153 bulk.t116 233.526
R1306 bulk.n145 bulk.t106 233.526
R1307 bulk.n137 bulk.t126 233.526
R1308 bulk.n129 bulk.t243 233.526
R1309 bulk.n121 bulk.t218 233.526
R1310 bulk.n113 bulk.t203 233.526
R1311 bulk.n105 bulk.t189 233.526
R1312 bulk.n335 bulk.t272 233.526
R1313 bulk.n87 bulk.t291 233.526
R1314 bulk.n368 bulk.t14 233.526
R1315 bulk.n280 bulk.n279 220.689
R1316 bulk.n345 bulk.n344 220.689
R1317 bulk.n226 bulk.n225 165.517
R1318 bulk.n42 bulk.n41 165.517
R1319 bulk.n522 bulk.n521 82.758
R1320 bulk.n376 bulk.n375 82.758
R1321 bulk.n11 bulk.n10 27.586
R1322 bulk.n67 bulk.n66 27.586
R1323 bulk.n505 bulk.t251 26.241
R1324 bulk.n214 bulk.t95 26.241
R1325 bulk.n257 bulk.t196 23.906
R1326 bulk.n552 bulk.t60 23.906
R1327 bulk.n343 bulk.t275 23.906
R1328 bulk.n71 bulk.t294 23.906
R1329 bulk.n394 bulk.t17 23.841
R1330 bulk.n506 bulk.t162 23.841
R1331 bulk.n103 bulk.t159 23.841
R1332 bulk.n215 bulk.t307 23.841
R1333 bulk.n398 bulk.n397 19.8
R1334 bulk.n402 bulk.n401 19.8
R1335 bulk.n406 bulk.n405 19.8
R1336 bulk.n410 bulk.n409 19.8
R1337 bulk.n414 bulk.n413 19.8
R1338 bulk.n418 bulk.n417 19.8
R1339 bulk.n422 bulk.n421 19.8
R1340 bulk.n426 bulk.n425 19.8
R1341 bulk.n430 bulk.n429 19.8
R1342 bulk.n434 bulk.n433 19.8
R1343 bulk.n438 bulk.n437 19.8
R1344 bulk.n442 bulk.n441 19.8
R1345 bulk.n446 bulk.n445 19.8
R1346 bulk.n450 bulk.n449 19.8
R1347 bulk.n454 bulk.n453 19.8
R1348 bulk.n458 bulk.n457 19.8
R1349 bulk.n462 bulk.n461 19.8
R1350 bulk.n466 bulk.n465 19.8
R1351 bulk.n470 bulk.n469 19.8
R1352 bulk.n474 bulk.n473 19.8
R1353 bulk.n478 bulk.n477 19.8
R1354 bulk.n482 bulk.n481 19.8
R1355 bulk.n486 bulk.n485 19.8
R1356 bulk.n490 bulk.n489 19.8
R1357 bulk.n494 bulk.n493 19.8
R1358 bulk.n498 bulk.n497 19.8
R1359 bulk.n502 bulk.n501 19.8
R1360 bulk.n502 bulk.t250 19.8
R1361 bulk.n107 bulk.n106 19.8
R1362 bulk.n111 bulk.n110 19.8
R1363 bulk.n115 bulk.n114 19.8
R1364 bulk.n119 bulk.n118 19.8
R1365 bulk.n123 bulk.n122 19.8
R1366 bulk.n127 bulk.n126 19.8
R1367 bulk.n131 bulk.n130 19.8
R1368 bulk.n135 bulk.n134 19.8
R1369 bulk.n139 bulk.n138 19.8
R1370 bulk.n143 bulk.n142 19.8
R1371 bulk.n147 bulk.n146 19.8
R1372 bulk.n151 bulk.n150 19.8
R1373 bulk.n155 bulk.n154 19.8
R1374 bulk.n159 bulk.n158 19.8
R1375 bulk.n163 bulk.n162 19.8
R1376 bulk.n167 bulk.n166 19.8
R1377 bulk.n171 bulk.n170 19.8
R1378 bulk.n175 bulk.n174 19.8
R1379 bulk.n179 bulk.n178 19.8
R1380 bulk.n183 bulk.n182 19.8
R1381 bulk.n187 bulk.n186 19.8
R1382 bulk.n191 bulk.n190 19.8
R1383 bulk.n195 bulk.n194 19.8
R1384 bulk.n199 bulk.n198 19.8
R1385 bulk.n203 bulk.n202 19.8
R1386 bulk.n207 bulk.n206 19.8
R1387 bulk.n211 bulk.n210 19.8
R1388 bulk.n211 bulk.t94 19.8
R1389 bulk.n558 bulk.t61 17.4
R1390 bulk.n260 bulk.t197 17.4
R1391 bulk.n527 bulk.t163 17.4
R1392 bulk.n26 bulk.t308 17.4
R1393 bulk.n76 bulk.t293 17.4
R1394 bulk.n350 bulk.t274 17.4
R1395 bulk.n371 bulk.t16 17.4
R1396 bulk.n37 bulk.t158 17.4
R1397 bulk.n278 bulk.n277 13.361
R1398 bulk.n9 bulk.n8 13.361
R1399 bulk.n295 bulk.n294 13.361
R1400 bulk.n29 bulk.n28 13.361
R1401 bulk.n74 bulk.n73 13.361
R1402 bulk.n309 bulk.n308 13.361
R1403 bulk.n297 bulk.n296 13.361
R1404 bulk.n31 bulk.n30 13.361
R1405 bulk.n373 bulk.n372 9.3
R1406 bulk.n390 bulk.n389 9.3
R1407 bulk.n340 bulk.n339 9.3
R1408 bulk.n352 bulk.n351 9.3
R1409 bulk.n78 bulk.n77 9.3
R1410 bulk.n63 bulk.n62 9.3
R1411 bulk.n39 bulk.n38 9.3
R1412 bulk.n99 bulk.n47 9.3
R1413 bulk.n529 bulk.n528 9.3
R1414 bulk.n517 bulk.n516 9.3
R1415 bulk.n254 bulk.n253 9.3
R1416 bulk.n262 bulk.n261 9.3
R1417 bulk.n560 bulk.n559 9.3
R1418 bulk.n549 bulk.n548 9.3
R1419 bulk.n223 bulk.n222 9.3
R1420 bulk.n233 bulk.n27 9.3
R1421 bulk.n261 bulk.n260 8.5
R1422 bulk.n27 bulk.n26 8.5
R1423 bulk.n77 bulk.n76 8.5
R1424 bulk.n372 bulk.n371 8.5
R1425 bulk.n351 bulk.n350 8.5
R1426 bulk.n38 bulk.n37 8.499
R1427 bulk.n528 bulk.n527 8.499
R1428 bulk.n559 bulk.n558 8.499
R1429 bulk.n399 bulk.n398 6.441
R1430 bulk.n403 bulk.n402 6.441
R1431 bulk.n407 bulk.n406 6.441
R1432 bulk.n411 bulk.n410 6.441
R1433 bulk.n415 bulk.n414 6.441
R1434 bulk.n419 bulk.n418 6.441
R1435 bulk.n423 bulk.n422 6.441
R1436 bulk.n427 bulk.n426 6.441
R1437 bulk.n431 bulk.n430 6.441
R1438 bulk.n435 bulk.n434 6.441
R1439 bulk.n439 bulk.n438 6.441
R1440 bulk.n443 bulk.n442 6.441
R1441 bulk.n447 bulk.n446 6.441
R1442 bulk.n451 bulk.n450 6.441
R1443 bulk.n455 bulk.n454 6.441
R1444 bulk.n459 bulk.n458 6.441
R1445 bulk.n463 bulk.n462 6.441
R1446 bulk.n467 bulk.n466 6.441
R1447 bulk.n471 bulk.n470 6.441
R1448 bulk.n475 bulk.n474 6.441
R1449 bulk.n479 bulk.n478 6.441
R1450 bulk.n483 bulk.n482 6.441
R1451 bulk.n487 bulk.n486 6.441
R1452 bulk.n491 bulk.n490 6.441
R1453 bulk.n495 bulk.n494 6.441
R1454 bulk.n499 bulk.n498 6.441
R1455 bulk.n503 bulk.n502 6.441
R1456 bulk.n108 bulk.n107 6.441
R1457 bulk.n112 bulk.n111 6.441
R1458 bulk.n116 bulk.n115 6.441
R1459 bulk.n120 bulk.n119 6.441
R1460 bulk.n124 bulk.n123 6.441
R1461 bulk.n128 bulk.n127 6.441
R1462 bulk.n132 bulk.n131 6.441
R1463 bulk.n136 bulk.n135 6.441
R1464 bulk.n140 bulk.n139 6.441
R1465 bulk.n144 bulk.n143 6.441
R1466 bulk.n148 bulk.n147 6.441
R1467 bulk.n152 bulk.n151 6.441
R1468 bulk.n156 bulk.n155 6.441
R1469 bulk.n160 bulk.n159 6.441
R1470 bulk.n164 bulk.n163 6.441
R1471 bulk.n168 bulk.n167 6.441
R1472 bulk.n172 bulk.n171 6.441
R1473 bulk.n176 bulk.n175 6.441
R1474 bulk.n180 bulk.n179 6.441
R1475 bulk.n184 bulk.n183 6.441
R1476 bulk.n188 bulk.n187 6.441
R1477 bulk.n192 bulk.n191 6.441
R1478 bulk.n196 bulk.n195 6.441
R1479 bulk.n200 bulk.n199 6.441
R1480 bulk.n204 bulk.n203 6.441
R1481 bulk.n208 bulk.n207 6.441
R1482 bulk.n212 bulk.n211 6.441
R1483 bulk.n40 bulk.n31 4.558
R1484 bulk.n391 bulk.n380 4.558
R1485 bulk.n374 bulk.n297 4.558
R1486 bulk.n349 bulk.n309 4.558
R1487 bulk.n341 bulk.n313 4.558
R1488 bulk.n65 bulk.n64 4.558
R1489 bulk.n75 bulk.n74 4.558
R1490 bulk.n100 bulk.n46 4.558
R1491 bulk.n224 bulk.n216 4.558
R1492 bulk.n526 bulk.n295 4.558
R1493 bulk.n518 bulk.n507 4.558
R1494 bulk.n255 bulk.n14 4.558
R1495 bulk.n259 bulk.n9 4.558
R1496 bulk.n557 bulk.n278 4.558
R1497 bulk.n550 bulk.n283 4.558
R1498 bulk.n232 bulk.n29 4.558
R1499 bulk.n530 bulk.n293 1.161
R1500 bulk.n511 bulk.n509 1.161
R1501 bulk.n237 bulk.n236 1.161
R1502 bulk.n240 bulk.n239 1.161
R1503 bulk.n245 bulk.n244 1.161
R1504 bulk.n248 bulk.n247 1.161
R1505 bulk.n266 bulk.n265 1.161
R1506 bulk.n273 bulk.n272 1.161
R1507 bulk.n545 bulk.n287 1.161
R1508 bulk.n538 bulk.n289 1.161
R1509 bulk.n537 bulk.n291 1.161
R1510 bulk.n94 bulk.n49 1.161
R1511 bulk.n93 bulk.n51 1.161
R1512 bulk.n90 bulk.n55 1.161
R1513 bulk.n89 bulk.n57 1.161
R1514 bulk.n326 bulk.n325 1.161
R1515 bulk.n357 bulk.n356 1.161
R1516 bulk.n363 bulk.n362 1.161
R1517 bulk.n366 bulk.n365 1.161
R1518 bulk.n384 bulk.n383 1.159
R1519 bulk.n332 bulk.n331 1.159
R1520 bulk.n333 bulk.n320 1.159
R1521 bulk.n35 bulk.n33 1.159
R1522 bulk.n220 bulk.n218 1.159
R1523 bulk.n242 bulk.n22 1.159
R1524 bulk.n270 bulk.n1 1.159
R1525 bulk.n562 bulk.n276 1.159
R1526 bulk.n546 bulk.n285 1.159
R1527 bulk.n91 bulk.n53 1.159
R1528 bulk.n337 bulk.n315 1.159
R1529 bulk.n354 bulk.n307 1.159
R1530 bulk.n370 bulk.n299 1.159
R1531 bulk.n387 bulk.n386 1.142
R1532 bulk.n378 bulk.n377 1.142
R1533 bulk.n302 bulk.n301 1.142
R1534 bulk.n305 bulk.n304 1.142
R1535 bulk.n347 bulk.n346 1.142
R1536 bulk.n312 bulk.n311 1.142
R1537 bulk.n318 bulk.n317 1.142
R1538 bulk.n323 bulk.n322 1.142
R1539 bulk.n60 bulk.n59 1.142
R1540 bulk.n69 bulk.n68 1.142
R1541 bulk.n81 bulk.n80 1.142
R1542 bulk.n85 bulk.n84 1.142
R1543 bulk.n97 bulk.n96 1.142
R1544 bulk.n44 bulk.n43 1.142
R1545 bulk.n514 bulk.n513 1.142
R1546 bulk.n524 bulk.n523 1.142
R1547 bulk.n535 bulk.n534 1.142
R1548 bulk.n541 bulk.n540 1.142
R1549 bulk.n282 bulk.n281 1.142
R1550 bulk.n555 bulk.n554 1.142
R1551 bulk.n567 bulk.n566 1.142
R1552 bulk.n4 bulk.n3 1.142
R1553 bulk.n7 bulk.n6 1.142
R1554 bulk.n13 bulk.n12 1.142
R1555 bulk.n17 bulk.n16 1.142
R1556 bulk.n20 bulk.n19 1.142
R1557 bulk.n25 bulk.n24 1.142
R1558 bulk.n228 bulk.n227 1.142
R1559 bulk.n386 bulk.n385 1.142
R1560 bulk.n377 bulk.n376 1.142
R1561 bulk.n299 bulk.n298 1.142
R1562 bulk.n301 bulk.n300 1.142
R1563 bulk.n365 bulk.n364 1.142
R1564 bulk.n362 bulk.n361 1.142
R1565 bulk.n304 bulk.n303 1.142
R1566 bulk.n356 bulk.n355 1.142
R1567 bulk.n307 bulk.n306 1.142
R1568 bulk.n346 bulk.n345 1.142
R1569 bulk.n311 bulk.n310 1.142
R1570 bulk.n315 bulk.n314 1.142
R1571 bulk.n317 bulk.n316 1.142
R1572 bulk.n320 bulk.n319 1.142
R1573 bulk.n331 bulk.n330 1.142
R1574 bulk.n322 bulk.n321 1.142
R1575 bulk.n325 bulk.n324 1.142
R1576 bulk.n59 bulk.n58 1.142
R1577 bulk.n68 bulk.n67 1.142
R1578 bulk.n80 bulk.n79 1.142
R1579 bulk.n84 bulk.n83 1.142
R1580 bulk.n57 bulk.n56 1.142
R1581 bulk.n55 bulk.n54 1.142
R1582 bulk.n53 bulk.n52 1.142
R1583 bulk.n51 bulk.n50 1.142
R1584 bulk.n49 bulk.n48 1.142
R1585 bulk.n96 bulk.n95 1.142
R1586 bulk.n43 bulk.n42 1.142
R1587 bulk.n513 bulk.n512 1.142
R1588 bulk.n523 bulk.n522 1.142
R1589 bulk.n293 bulk.n292 1.142
R1590 bulk.n534 bulk.n533 1.142
R1591 bulk.n291 bulk.n290 1.142
R1592 bulk.n289 bulk.n288 1.142
R1593 bulk.n540 bulk.n539 1.142
R1594 bulk.n287 bulk.n286 1.142
R1595 bulk.n285 bulk.n284 1.142
R1596 bulk.n281 bulk.n280 1.142
R1597 bulk.n554 bulk.n553 1.142
R1598 bulk.n276 bulk.n275 1.142
R1599 bulk.n566 bulk.n565 1.142
R1600 bulk.n272 bulk.n271 1.142
R1601 bulk.n1 bulk.n0 1.142
R1602 bulk.n3 bulk.n2 1.142
R1603 bulk.n265 bulk.n264 1.142
R1604 bulk.n6 bulk.n5 1.142
R1605 bulk.n12 bulk.n11 1.142
R1606 bulk.n16 bulk.n15 1.142
R1607 bulk.n19 bulk.n18 1.142
R1608 bulk.n247 bulk.n246 1.142
R1609 bulk.n244 bulk.n243 1.142
R1610 bulk.n22 bulk.n21 1.142
R1611 bulk.n239 bulk.n238 1.142
R1612 bulk.n236 bulk.n235 1.142
R1613 bulk.n24 bulk.n23 1.142
R1614 bulk.n227 bulk.n226 1.142
R1615 bulk.n104 bulk.n103 0.069
R1616 bulk.n215 bulk.n214 0.069
R1617 bulk.n395 bulk.n394 0.069
R1618 bulk.n506 bulk.n505 0.069
R1619 bulk.n383 bulk.n382 0.053
R1620 bulk.n33 bulk.n32 0.053
R1621 bulk.n509 bulk.n508 0.053
R1622 bulk.n218 bulk.n217 0.053
R1623 bulk.n366 bulk.n363 0.026
R1624 bulk.n90 bulk.n89 0.026
R1625 bulk.n94 bulk.n93 0.026
R1626 bulk.n538 bulk.n537 0.026
R1627 bulk.n248 bulk.n245 0.026
R1628 bulk.n240 bulk.n237 0.026
R1629 bulk.n367 bulk.n366 0.025
R1630 bulk.n327 bulk.n326 0.025
R1631 bulk.n267 bulk.n266 0.025
R1632 bulk.n384 bulk.n381 0.025
R1633 bulk.n537 bulk.n536 0.025
R1634 bulk.n536 bulk.n535 0.024
R1635 bulk.n245 bulk.n242 0.023
R1636 bulk.n273 bulk.n270 0.023
R1637 bulk.n546 bulk.n545 0.023
R1638 bulk.n91 bulk.n90 0.023
R1639 bulk.n357 bulk.n354 0.023
R1640 bulk.n266 bulk.n263 0.022
R1641 bulk.n542 bulk.n538 0.022
R1642 bulk.n98 bulk.n94 0.022
R1643 bulk.n363 bulk.n360 0.022
R1644 bulk.n515 bulk.n511 0.022
R1645 bulk.n252 bulk.n17 0.021
R1646 bulk.n267 bulk.n4 0.021
R1647 bulk.n82 bulk.n81 0.021
R1648 bulk.n327 bulk.n323 0.021
R1649 bulk.n334 bulk.n318 0.021
R1650 bulk.n367 bulk.n302 0.021
R1651 bulk.n334 bulk.n333 0.021
R1652 bulk.n237 bulk.n234 0.021
R1653 bulk.n252 bulk.n251 0.021
R1654 bulk.n86 bulk.n82 0.021
R1655 bulk.n531 bulk.n530 0.02
R1656 bulk.n70 bulk.n69 0.019
R1657 bulk.n258 bulk.n13 0.019
R1658 bulk.n342 bulk.n312 0.017
R1659 bulk.n551 bulk.n282 0.017
R1660 bulk.n556 bulk.n555 0.017
R1661 bulk.n234 bulk.n25 0.017
R1662 bulk.n388 bulk.n387 0.017
R1663 bulk.n360 bulk.n305 0.017
R1664 bulk.n348 bulk.n347 0.017
R1665 bulk.n61 bulk.n60 0.017
R1666 bulk.n86 bulk.n85 0.017
R1667 bulk.n98 bulk.n97 0.017
R1668 bulk.n515 bulk.n514 0.017
R1669 bulk.n542 bulk.n541 0.017
R1670 bulk.n263 bulk.n7 0.017
R1671 bulk.n251 bulk.n20 0.017
R1672 bulk.n379 bulk.n378 0.017
R1673 bulk.n45 bulk.n44 0.017
R1674 bulk.n525 bulk.n524 0.017
R1675 bulk.n568 bulk.n567 0.017
R1676 bulk.n229 bulk.n228 0.017
R1677 bulk.n511 bulk.n510 0.016
R1678 bulk.n388 bulk.n384 0.012
R1679 bulk.n333 bulk.n332 0.012
R1680 bulk.n105 bulk.n104 0.012
R1681 bulk.n108 bulk.n105 0.012
R1682 bulk.n109 bulk.n108 0.012
R1683 bulk.n112 bulk.n109 0.012
R1684 bulk.n113 bulk.n112 0.012
R1685 bulk.n116 bulk.n113 0.012
R1686 bulk.n117 bulk.n116 0.012
R1687 bulk.n120 bulk.n117 0.012
R1688 bulk.n121 bulk.n120 0.012
R1689 bulk.n124 bulk.n121 0.012
R1690 bulk.n125 bulk.n124 0.012
R1691 bulk.n128 bulk.n125 0.012
R1692 bulk.n129 bulk.n128 0.012
R1693 bulk.n132 bulk.n129 0.012
R1694 bulk.n133 bulk.n132 0.012
R1695 bulk.n136 bulk.n133 0.012
R1696 bulk.n137 bulk.n136 0.012
R1697 bulk.n140 bulk.n137 0.012
R1698 bulk.n141 bulk.n140 0.012
R1699 bulk.n144 bulk.n141 0.012
R1700 bulk.n145 bulk.n144 0.012
R1701 bulk.n148 bulk.n145 0.012
R1702 bulk.n149 bulk.n148 0.012
R1703 bulk.n152 bulk.n149 0.012
R1704 bulk.n153 bulk.n152 0.012
R1705 bulk.n156 bulk.n153 0.012
R1706 bulk.n157 bulk.n156 0.012
R1707 bulk.n160 bulk.n157 0.012
R1708 bulk.n161 bulk.n160 0.012
R1709 bulk.n164 bulk.n161 0.012
R1710 bulk.n165 bulk.n164 0.012
R1711 bulk.n168 bulk.n165 0.012
R1712 bulk.n169 bulk.n168 0.012
R1713 bulk.n172 bulk.n169 0.012
R1714 bulk.n173 bulk.n172 0.012
R1715 bulk.n176 bulk.n173 0.012
R1716 bulk.n177 bulk.n176 0.012
R1717 bulk.n180 bulk.n177 0.012
R1718 bulk.n181 bulk.n180 0.012
R1719 bulk.n184 bulk.n181 0.012
R1720 bulk.n185 bulk.n184 0.012
R1721 bulk.n188 bulk.n185 0.012
R1722 bulk.n189 bulk.n188 0.012
R1723 bulk.n192 bulk.n189 0.012
R1724 bulk.n193 bulk.n192 0.012
R1725 bulk.n196 bulk.n193 0.012
R1726 bulk.n197 bulk.n196 0.012
R1727 bulk.n200 bulk.n197 0.012
R1728 bulk.n201 bulk.n200 0.012
R1729 bulk.n204 bulk.n201 0.012
R1730 bulk.n205 bulk.n204 0.012
R1731 bulk.n208 bulk.n205 0.012
R1732 bulk.n209 bulk.n208 0.012
R1733 bulk.n212 bulk.n209 0.012
R1734 bulk.n213 bulk.n212 0.012
R1735 bulk.n214 bulk.n213 0.012
R1736 bulk.n396 bulk.n395 0.012
R1737 bulk.n399 bulk.n396 0.012
R1738 bulk.n400 bulk.n399 0.012
R1739 bulk.n403 bulk.n400 0.012
R1740 bulk.n404 bulk.n403 0.012
R1741 bulk.n407 bulk.n404 0.012
R1742 bulk.n408 bulk.n407 0.012
R1743 bulk.n411 bulk.n408 0.012
R1744 bulk.n412 bulk.n411 0.012
R1745 bulk.n415 bulk.n412 0.012
R1746 bulk.n416 bulk.n415 0.012
R1747 bulk.n419 bulk.n416 0.012
R1748 bulk.n420 bulk.n419 0.012
R1749 bulk.n423 bulk.n420 0.012
R1750 bulk.n424 bulk.n423 0.012
R1751 bulk.n427 bulk.n424 0.012
R1752 bulk.n428 bulk.n427 0.012
R1753 bulk.n431 bulk.n428 0.012
R1754 bulk.n432 bulk.n431 0.012
R1755 bulk.n435 bulk.n432 0.012
R1756 bulk.n436 bulk.n435 0.012
R1757 bulk.n439 bulk.n436 0.012
R1758 bulk.n440 bulk.n439 0.012
R1759 bulk.n443 bulk.n440 0.012
R1760 bulk.n444 bulk.n443 0.012
R1761 bulk.n447 bulk.n444 0.012
R1762 bulk.n448 bulk.n447 0.012
R1763 bulk.n451 bulk.n448 0.012
R1764 bulk.n452 bulk.n451 0.012
R1765 bulk.n455 bulk.n452 0.012
R1766 bulk.n456 bulk.n455 0.012
R1767 bulk.n459 bulk.n456 0.012
R1768 bulk.n460 bulk.n459 0.012
R1769 bulk.n463 bulk.n460 0.012
R1770 bulk.n464 bulk.n463 0.012
R1771 bulk.n467 bulk.n464 0.012
R1772 bulk.n468 bulk.n467 0.012
R1773 bulk.n471 bulk.n468 0.012
R1774 bulk.n472 bulk.n471 0.012
R1775 bulk.n475 bulk.n472 0.012
R1776 bulk.n476 bulk.n475 0.012
R1777 bulk.n479 bulk.n476 0.012
R1778 bulk.n480 bulk.n479 0.012
R1779 bulk.n483 bulk.n480 0.012
R1780 bulk.n484 bulk.n483 0.012
R1781 bulk.n487 bulk.n484 0.012
R1782 bulk.n488 bulk.n487 0.012
R1783 bulk.n491 bulk.n488 0.012
R1784 bulk.n492 bulk.n491 0.012
R1785 bulk.n495 bulk.n492 0.012
R1786 bulk.n496 bulk.n495 0.012
R1787 bulk.n499 bulk.n496 0.012
R1788 bulk.n500 bulk.n499 0.012
R1789 bulk.n503 bulk.n500 0.012
R1790 bulk.n504 bulk.n503 0.012
R1791 bulk.n505 bulk.n504 0.012
R1792 bulk.n358 bulk.n357 0.011
R1793 bulk.n89 bulk.n88 0.011
R1794 bulk.n93 bulk.n92 0.011
R1795 bulk.n545 bulk.n544 0.011
R1796 bulk.n274 bulk.n273 0.011
R1797 bulk.n249 bulk.n248 0.011
R1798 bulk.n241 bulk.n240 0.011
R1799 bulk.n335 bulk.n334 0.01
R1800 bulk.n35 bulk.n34 0.01
R1801 bulk.n220 bulk.n219 0.01
R1802 bulk.n530 bulk.n529 0.01
R1803 bulk.n82 bulk.n78 0.008
R1804 bulk.n254 bulk.n252 0.008
R1805 bulk.n328 bulk.n327 0.007
R1806 bulk.n268 bulk.n267 0.007
R1807 bulk.n562 bulk.n561 0.007
R1808 bulk.n338 bulk.n337 0.007
R1809 bulk.n373 bulk.n370 0.007
R1810 bulk.n332 bulk.n329 0.007
R1811 bulk.n370 bulk.n369 0.007
R1812 bulk.n354 bulk.n353 0.007
R1813 bulk.n337 bulk.n336 0.007
R1814 bulk.n92 bulk.n91 0.007
R1815 bulk.n547 bulk.n546 0.007
R1816 bulk.n563 bulk.n562 0.007
R1817 bulk.n270 bulk.n269 0.007
R1818 bulk.n242 bulk.n241 0.007
R1819 bulk.n221 bulk.n220 0.007
R1820 bulk.n36 bulk.n35 0.007
R1821 bulk.n368 bulk.n367 0.006
R1822 bulk.n348 bulk.n343 0.006
R1823 bulk.n536 bulk.n532 0.006
R1824 bulk.n556 bulk.n552 0.005
R1825 bulk.n552 bulk.n551 0.005
R1826 bulk.n343 bulk.n342 0.005
R1827 bulk.n259 bulk.n258 0.005
R1828 bulk.n70 bulk.n65 0.005
R1829 bulk.n369 bulk.n368 0.005
R1830 bulk.n75 bulk.n72 0.005
R1831 bulk.n329 bulk.n328 0.004
R1832 bulk.n269 bulk.n268 0.004
R1833 bulk.n568 bulk.n564 0.004
R1834 bulk.n256 bulk.n255 0.004
R1835 bulk.n63 bulk.n61 0.004
R1836 bulk.n360 bulk.n359 0.004
R1837 bulk.n263 bulk.n262 0.004
R1838 bulk.n543 bulk.n542 0.004
R1839 bulk.n103 bulk.n102 0.003
R1840 bulk.n230 bulk.n215 0.003
R1841 bulk.n102 bulk.n45 0.003
R1842 bulk.n101 bulk.n100 0.003
R1843 bulk.n88 bulk.n87 0.003
R1844 bulk.n340 bulk.n338 0.003
R1845 bulk.n379 bulk.n374 0.003
R1846 bulk.n393 bulk.n392 0.003
R1847 bulk.n394 bulk.n393 0.003
R1848 bulk.n520 bulk.n506 0.003
R1849 bulk.n230 bulk.n229 0.003
R1850 bulk.n232 bulk.n231 0.003
R1851 bulk.n250 bulk.n249 0.003
R1852 bulk bulk.n568 0.003
R1853 bulk.n561 bulk.n560 0.003
R1854 bulk.n526 bulk.n525 0.003
R1855 bulk.n520 bulk.n519 0.003
R1856 bulk.n87 bulk.n86 0.003
R1857 bulk.n251 bulk.n250 0.003
R1858 bulk.n40 bulk.n39 0.002
R1859 bulk.n78 bulk.n75 0.002
R1860 bulk.n352 bulk.n349 0.002
R1861 bulk.n353 bulk.n352 0.002
R1862 bulk.n359 bulk.n358 0.002
R1863 bulk.n391 bulk.n390 0.002
R1864 bulk.n224 bulk.n223 0.002
R1865 bulk.n255 bulk.n254 0.002
R1866 bulk.n550 bulk.n549 0.002
R1867 bulk.n549 bulk.n547 0.002
R1868 bulk.n544 bulk.n543 0.002
R1869 bulk.n518 bulk.n517 0.002
R1870 bulk.n390 bulk.n388 0.002
R1871 bulk.n517 bulk.n515 0.002
R1872 bulk.n72 bulk.n71 0.001
R1873 bulk.n532 bulk.n531 0.001
R1874 bulk.n257 bulk.n256 0.001
R1875 bulk.n39 bulk.n36 0.001
R1876 bulk.n45 bulk.n40 0.001
R1877 bulk.n102 bulk.n101 0.001
R1878 bulk.n100 bulk.n99 0.001
R1879 bulk.n65 bulk.n63 0.001
R1880 bulk.n336 bulk.n335 0.001
R1881 bulk.n341 bulk.n340 0.001
R1882 bulk.n374 bulk.n373 0.001
R1883 bulk.n393 bulk.n379 0.001
R1884 bulk.n392 bulk.n391 0.001
R1885 bulk.n223 bulk.n221 0.001
R1886 bulk.n229 bulk.n224 0.001
R1887 bulk.n231 bulk.n230 0.001
R1888 bulk.n233 bulk.n232 0.001
R1889 bulk.n262 bulk.n259 0.001
R1890 bulk bulk.n274 0.001
R1891 bulk.n564 bulk.n563 0.001
R1892 bulk.n560 bulk.n557 0.001
R1893 bulk.n529 bulk.n526 0.001
R1894 bulk.n525 bulk.n520 0.001
R1895 bulk.n519 bulk.n518 0.001
R1896 bulk.n71 bulk.n70 0.001
R1897 bulk.n258 bulk.n257 0.001
R1898 bulk.n349 bulk.n348 0.001
R1899 bulk.n99 bulk.n98 0.001
R1900 bulk.n342 bulk.n341 0.001
R1901 bulk.n551 bulk.n550 0.001
R1902 bulk.n557 bulk.n556 0.001
R1903 bulk.n234 bulk.n233 0.001
R1904 bias2.n0 bias2.t23 286.107
R1905 bias2.n1 bias2.t20 286.107
R1906 bias2.n2 bias2.t26 286.107
R1907 bias2.n3 bias2.t22 286.107
R1908 bias2.n4 bias2.t5 286.107
R1909 bias2.n5 bias2.t2 286.107
R1910 bias2.n6 bias2.t0 286.107
R1911 bias2.n7 bias2.t4 286.107
R1912 bias2.n8 bias2.t19 286.107
R1913 bias2.n9 bias2.t13 286.107
R1914 bias2.n10 bias2.t10 286.107
R1915 bias2.n11 bias2.t8 286.107
R1916 bias2.n12 bias2.t15 286.107
R1917 bias2.n13 bias2.t12 286.107
R1918 bias2.n27 bias2.t9 233.526
R1919 bias2.n26 bias2.t11 233.526
R1920 bias2.n25 bias2.t14 233.526
R1921 bias2.n24 bias2.t16 233.526
R1922 bias2.n23 bias2.t17 233.526
R1923 bias2.n22 bias2.t18 233.526
R1924 bias2.n21 bias2.t3 233.526
R1925 bias2.n20 bias2.t6 233.526
R1926 bias2.n19 bias2.t7 233.526
R1927 bias2.n18 bias2.t1 233.526
R1928 bias2.n17 bias2.t21 233.526
R1929 bias2.n16 bias2.t24 233.526
R1930 bias2.n15 bias2.t25 233.526
R1931 bias2.n14 bias2.t27 233.526
R1932 bias2.n35 bias2.n34 1.375
R1933 bias2.n28 bias2.n27 0.293
R1934 bias2.n15 bias2.n14 0.203
R1935 bias2.n16 bias2.n15 0.203
R1936 bias2.n17 bias2.n16 0.203
R1937 bias2.n18 bias2.n17 0.203
R1938 bias2.n19 bias2.n18 0.203
R1939 bias2.n20 bias2.n19 0.203
R1940 bias2.n21 bias2.n20 0.203
R1941 bias2.n22 bias2.n21 0.203
R1942 bias2.n23 bias2.n22 0.203
R1943 bias2.n24 bias2.n23 0.203
R1944 bias2.n25 bias2.n24 0.203
R1945 bias2.n26 bias2.n25 0.203
R1946 bias2.n27 bias2.n26 0.203
R1947 bias2.n1 bias2.n0 0.203
R1948 bias2.n2 bias2.n1 0.203
R1949 bias2.n3 bias2.n2 0.203
R1950 bias2.n4 bias2.n3 0.203
R1951 bias2.n5 bias2.n4 0.203
R1952 bias2.n6 bias2.n5 0.203
R1953 bias2.n7 bias2.n6 0.203
R1954 bias2.n8 bias2.n7 0.203
R1955 bias2.n9 bias2.n8 0.203
R1956 bias2.n10 bias2.n9 0.203
R1957 bias2.n11 bias2.n10 0.203
R1958 bias2.n12 bias2.n11 0.203
R1959 bias2.n13 bias2.n12 0.203
R1960 bias2.n34 bias2.n13 0.191
R1961 bias2 bias2.n61 0.095
R1962 bias2.n60 bias2.n59 0.086
R1963 bias2.n30 bias2.n29 0.067
R1964 bias2.n31 bias2.n30 0.067
R1965 bias2.n32 bias2.n31 0.067
R1966 bias2.n33 bias2.n32 0.067
R1967 bias2.n46 bias2.n45 0.027
R1968 bias2.n60 bias2.n58 0.027
R1969 bias2.n45 bias2.n44 0.025
R1970 bias2.n43 bias2.n42 0.025
R1971 bias2.n42 bias2.n41 0.025
R1972 bias2.n41 bias2.n40 0.025
R1973 bias2.n40 bias2.n39 0.025
R1974 bias2.n39 bias2.n38 0.025
R1975 bias2.n38 bias2.n37 0.025
R1976 bias2.n37 bias2.n36 0.025
R1977 bias2.n36 bias2.n35 0.025
R1978 bias2.n46 bias2.n43 0.024
R1979 bias2.n61 bias2.n60 0.018
R1980 bias2.n58 bias2.n57 0.006
R1981 bias2.n57 bias2.n56 0.006
R1982 bias2.n55 bias2.n54 0.006
R1983 bias2.n54 bias2.n53 0.006
R1984 bias2.n53 bias2.n52 0.006
R1985 bias2.n52 bias2.n51 0.006
R1986 bias2.n51 bias2.n50 0.006
R1987 bias2.n50 bias2.n49 0.006
R1988 bias2.n49 bias2.n48 0.006
R1989 bias2.n48 bias2.n47 0.006
R1990 bias2.n56 bias2.n55 0.005
R1991 bias2.n29 bias2.n28 0.004
R1992 bias2.n34 bias2.n33 0.004
R1993 bias2.n56 bias2.n46 0.001
R1994 tank_out.n445 tank_out.t15 19.8
R1995 tank_out.n415 tank_out.t12 19.8
R1996 tank_out.n415 tank_out.t18 19.8
R1997 tank_out.n385 tank_out.t19 19.8
R1998 tank_out.n385 tank_out.t16 19.8
R1999 tank_out.n355 tank_out.t17 19.8
R2000 tank_out.n355 tank_out.t13 19.8
R2001 tank_out.n325 tank_out.t14 19.8
R2002 tank_out.n325 tank_out.t11 19.8
R2003 tank_out.n295 tank_out.t8 19.8
R2004 tank_out.n295 tank_out.t10 19.8
R2005 tank_out.n265 tank_out.t23 19.8
R2006 tank_out.n265 tank_out.t9 19.8
R2007 tank_out.n235 tank_out.t27 19.8
R2008 tank_out.n235 tank_out.t24 19.8
R2009 tank_out.n19 tank_out.t25 19.8
R2010 tank_out.n19 tank_out.t21 19.8
R2011 tank_out.n49 tank_out.t22 19.8
R2012 tank_out.n49 tank_out.t20 19.8
R2013 tank_out.n79 tank_out.t5 19.8
R2014 tank_out.n79 tank_out.t26 19.8
R2015 tank_out.n109 tank_out.t1 19.8
R2016 tank_out.n109 tank_out.t6 19.8
R2017 tank_out.n139 tank_out.t7 19.8
R2018 tank_out.n139 tank_out.t3 19.8
R2019 tank_out.n169 tank_out.t4 19.8
R2020 tank_out.n169 tank_out.t2 19.8
R2021 tank_out.n199 tank_out.t0 19.8
R2022 tank_out.n416 tank_out.n415 8.5
R2023 tank_out.n386 tank_out.n385 8.5
R2024 tank_out.n356 tank_out.n355 8.5
R2025 tank_out.n326 tank_out.n325 8.5
R2026 tank_out.n296 tank_out.n295 8.5
R2027 tank_out.n266 tank_out.n265 8.5
R2028 tank_out.n236 tank_out.n235 8.5
R2029 tank_out.n20 tank_out.n19 8.5
R2030 tank_out.n50 tank_out.n49 8.5
R2031 tank_out.n80 tank_out.n79 8.5
R2032 tank_out.n110 tank_out.n109 8.5
R2033 tank_out.n140 tank_out.n139 8.5
R2034 tank_out.n170 tank_out.n169 8.5
R2035 tank_out.n200 tank_out.n199 8.5
R2036 tank_out.n446 tank_out.n445 8.5
R2037 tank_out.n435 tank_out.n434 7.529
R2038 tank_out.n405 tank_out.n404 7.529
R2039 tank_out.n375 tank_out.n374 7.529
R2040 tank_out.n345 tank_out.n344 7.529
R2041 tank_out.n315 tank_out.n314 7.529
R2042 tank_out.n285 tank_out.n284 7.529
R2043 tank_out.n255 tank_out.n254 7.529
R2044 tank_out.n225 tank_out.n224 7.529
R2045 tank_out.n9 tank_out.n8 7.529
R2046 tank_out.n39 tank_out.n38 7.529
R2047 tank_out.n69 tank_out.n68 7.529
R2048 tank_out.n99 tank_out.n98 7.529
R2049 tank_out.n129 tank_out.n128 7.529
R2050 tank_out.n159 tank_out.n158 7.529
R2051 tank_out.n189 tank_out.n188 7.529
R2052 tank_out.n448 tank_out.n447 4.5
R2053 tank_out.n442 tank_out.n441 4.5
R2054 tank_out.n436 tank_out.n435 4.5
R2055 tank_out.n430 tank_out.n429 4.5
R2056 tank_out.n418 tank_out.n417 4.5
R2057 tank_out.n412 tank_out.n411 4.5
R2058 tank_out.n406 tank_out.n405 4.5
R2059 tank_out.n400 tank_out.n399 4.5
R2060 tank_out.n388 tank_out.n387 4.5
R2061 tank_out.n382 tank_out.n381 4.5
R2062 tank_out.n376 tank_out.n375 4.5
R2063 tank_out.n370 tank_out.n369 4.5
R2064 tank_out.n358 tank_out.n357 4.5
R2065 tank_out.n352 tank_out.n351 4.5
R2066 tank_out.n346 tank_out.n345 4.5
R2067 tank_out.n340 tank_out.n339 4.5
R2068 tank_out.n328 tank_out.n327 4.5
R2069 tank_out.n322 tank_out.n321 4.5
R2070 tank_out.n316 tank_out.n315 4.5
R2071 tank_out.n310 tank_out.n309 4.5
R2072 tank_out.n298 tank_out.n297 4.5
R2073 tank_out.n292 tank_out.n291 4.5
R2074 tank_out.n286 tank_out.n285 4.5
R2075 tank_out.n280 tank_out.n279 4.5
R2076 tank_out.n268 tank_out.n267 4.5
R2077 tank_out.n262 tank_out.n261 4.5
R2078 tank_out.n256 tank_out.n255 4.5
R2079 tank_out.n250 tank_out.n249 4.5
R2080 tank_out.n238 tank_out.n237 4.5
R2081 tank_out.n232 tank_out.n231 4.5
R2082 tank_out.n226 tank_out.n225 4.5
R2083 tank_out.n220 tank_out.n219 4.5
R2084 tank_out.n22 tank_out.n21 4.5
R2085 tank_out.n16 tank_out.n15 4.5
R2086 tank_out.n10 tank_out.n9 4.5
R2087 tank_out.n4 tank_out.n3 4.5
R2088 tank_out.n52 tank_out.n51 4.5
R2089 tank_out.n46 tank_out.n45 4.5
R2090 tank_out.n40 tank_out.n39 4.5
R2091 tank_out.n34 tank_out.n33 4.5
R2092 tank_out.n82 tank_out.n81 4.5
R2093 tank_out.n76 tank_out.n75 4.5
R2094 tank_out.n70 tank_out.n69 4.5
R2095 tank_out.n64 tank_out.n63 4.5
R2096 tank_out.n112 tank_out.n111 4.5
R2097 tank_out.n106 tank_out.n105 4.5
R2098 tank_out.n100 tank_out.n99 4.5
R2099 tank_out.n94 tank_out.n93 4.5
R2100 tank_out.n142 tank_out.n141 4.5
R2101 tank_out.n136 tank_out.n135 4.5
R2102 tank_out.n130 tank_out.n129 4.5
R2103 tank_out.n124 tank_out.n123 4.5
R2104 tank_out.n172 tank_out.n171 4.5
R2105 tank_out.n166 tank_out.n165 4.5
R2106 tank_out.n160 tank_out.n159 4.5
R2107 tank_out.n154 tank_out.n153 4.5
R2108 tank_out.n202 tank_out.n201 4.5
R2109 tank_out.n196 tank_out.n195 4.5
R2110 tank_out.n190 tank_out.n189 4.5
R2111 tank_out.n184 tank_out.n183 4.5
R2112 tank_out.n441 tank_out.n440 3.764
R2113 tank_out.n411 tank_out.n410 3.764
R2114 tank_out.n381 tank_out.n380 3.764
R2115 tank_out.n351 tank_out.n350 3.764
R2116 tank_out.n321 tank_out.n320 3.764
R2117 tank_out.n291 tank_out.n290 3.764
R2118 tank_out.n261 tank_out.n260 3.764
R2119 tank_out.n231 tank_out.n230 3.764
R2120 tank_out.n15 tank_out.n14 3.764
R2121 tank_out.n45 tank_out.n44 3.764
R2122 tank_out.n75 tank_out.n74 3.764
R2123 tank_out.n105 tank_out.n104 3.764
R2124 tank_out.n135 tank_out.n134 3.764
R2125 tank_out.n165 tank_out.n164 3.764
R2126 tank_out.n195 tank_out.n194 3.764
R2127 tank_out.n429 tank_out.n427 3.388
R2128 tank_out.n399 tank_out.n397 3.388
R2129 tank_out.n369 tank_out.n367 3.388
R2130 tank_out.n339 tank_out.n337 3.388
R2131 tank_out.n309 tank_out.n307 3.388
R2132 tank_out.n279 tank_out.n277 3.388
R2133 tank_out.n249 tank_out.n247 3.388
R2134 tank_out.n219 tank_out.n217 3.388
R2135 tank_out.n3 tank_out.n1 3.388
R2136 tank_out.n33 tank_out.n31 3.388
R2137 tank_out.n63 tank_out.n61 3.388
R2138 tank_out.n93 tank_out.n91 3.388
R2139 tank_out.n123 tank_out.n121 3.388
R2140 tank_out.n153 tank_out.n151 3.388
R2141 tank_out.n183 tank_out.n181 3.388
R2142 tank_out.n429 tank_out.n428 3.011
R2143 tank_out.n435 tank_out.n433 3.011
R2144 tank_out.n399 tank_out.n398 3.011
R2145 tank_out.n405 tank_out.n403 3.011
R2146 tank_out.n369 tank_out.n368 3.011
R2147 tank_out.n375 tank_out.n373 3.011
R2148 tank_out.n339 tank_out.n338 3.011
R2149 tank_out.n345 tank_out.n343 3.011
R2150 tank_out.n309 tank_out.n308 3.011
R2151 tank_out.n315 tank_out.n313 3.011
R2152 tank_out.n279 tank_out.n278 3.011
R2153 tank_out.n285 tank_out.n283 3.011
R2154 tank_out.n249 tank_out.n248 3.011
R2155 tank_out.n255 tank_out.n253 3.011
R2156 tank_out.n219 tank_out.n218 3.011
R2157 tank_out.n225 tank_out.n223 3.011
R2158 tank_out.n3 tank_out.n2 3.011
R2159 tank_out.n9 tank_out.n7 3.011
R2160 tank_out.n33 tank_out.n32 3.011
R2161 tank_out.n39 tank_out.n37 3.011
R2162 tank_out.n63 tank_out.n62 3.011
R2163 tank_out.n69 tank_out.n67 3.011
R2164 tank_out.n93 tank_out.n92 3.011
R2165 tank_out.n99 tank_out.n97 3.011
R2166 tank_out.n123 tank_out.n122 3.011
R2167 tank_out.n129 tank_out.n127 3.011
R2168 tank_out.n153 tank_out.n152 3.011
R2169 tank_out.n159 tank_out.n157 3.011
R2170 tank_out.n183 tank_out.n182 3.011
R2171 tank_out.n189 tank_out.n187 3.011
R2172 tank_out.n447 tank_out.n446 1.505
R2173 tank_out.n417 tank_out.n416 1.505
R2174 tank_out.n387 tank_out.n386 1.505
R2175 tank_out.n357 tank_out.n356 1.505
R2176 tank_out.n327 tank_out.n326 1.505
R2177 tank_out.n297 tank_out.n296 1.505
R2178 tank_out.n267 tank_out.n266 1.505
R2179 tank_out.n237 tank_out.n236 1.505
R2180 tank_out.n21 tank_out.n20 1.505
R2181 tank_out.n51 tank_out.n50 1.505
R2182 tank_out.n81 tank_out.n80 1.505
R2183 tank_out.n111 tank_out.n110 1.505
R2184 tank_out.n141 tank_out.n140 1.505
R2185 tank_out.n171 tank_out.n170 1.505
R2186 tank_out.n201 tank_out.n200 1.505
R2187 tank_out.n450 tank_out.n449 0.955
R2188 tank_out.n420 tank_out.n419 0.955
R2189 tank_out.n390 tank_out.n389 0.955
R2190 tank_out.n360 tank_out.n359 0.955
R2191 tank_out.n330 tank_out.n329 0.955
R2192 tank_out.n300 tank_out.n299 0.955
R2193 tank_out.n270 tank_out.n269 0.955
R2194 tank_out.n240 tank_out.n239 0.955
R2195 tank_out.n24 tank_out.n23 0.955
R2196 tank_out.n54 tank_out.n53 0.955
R2197 tank_out.n84 tank_out.n83 0.955
R2198 tank_out.n114 tank_out.n113 0.955
R2199 tank_out.n144 tank_out.n143 0.955
R2200 tank_out.n174 tank_out.n173 0.955
R2201 tank_out.n204 tank_out.n203 0.955
R2202 tank_out.n440 tank_out.n439 0.376
R2203 tank_out.n410 tank_out.n409 0.376
R2204 tank_out.n380 tank_out.n379 0.376
R2205 tank_out.n350 tank_out.n349 0.376
R2206 tank_out.n320 tank_out.n319 0.376
R2207 tank_out.n290 tank_out.n289 0.376
R2208 tank_out.n260 tank_out.n259 0.376
R2209 tank_out.n230 tank_out.n229 0.376
R2210 tank_out.n14 tank_out.n13 0.376
R2211 tank_out.n44 tank_out.n43 0.376
R2212 tank_out.n74 tank_out.n73 0.376
R2213 tank_out.n104 tank_out.n103 0.376
R2214 tank_out.n134 tank_out.n133 0.376
R2215 tank_out.n164 tank_out.n163 0.376
R2216 tank_out.n194 tank_out.n193 0.376
R2217 tank_out.n456 tank_out.n455 0.242
R2218 tank_out.n210 tank_out.n209 0.242
R2219 tank_out.n456 tank_out.n425 0.216
R2220 tank_out.n457 tank_out.n395 0.216
R2221 tank_out.n458 tank_out.n365 0.216
R2222 tank_out.n459 tank_out.n335 0.216
R2223 tank_out.n460 tank_out.n305 0.216
R2224 tank_out.n461 tank_out.n275 0.216
R2225 tank_out.n462 tank_out.n245 0.216
R2226 tank_out.n215 tank_out.n29 0.216
R2227 tank_out.n214 tank_out.n59 0.216
R2228 tank_out.n213 tank_out.n89 0.216
R2229 tank_out.n212 tank_out.n119 0.216
R2230 tank_out.n211 tank_out.n149 0.216
R2231 tank_out.n210 tank_out.n179 0.216
R2232 tank_out.n454 tank_out.n453 0.044
R2233 tank_out.n424 tank_out.n423 0.044
R2234 tank_out.n394 tank_out.n393 0.044
R2235 tank_out.n364 tank_out.n363 0.044
R2236 tank_out.n334 tank_out.n333 0.044
R2237 tank_out.n304 tank_out.n303 0.044
R2238 tank_out.n274 tank_out.n273 0.044
R2239 tank_out.n244 tank_out.n243 0.044
R2240 tank_out.n28 tank_out.n27 0.044
R2241 tank_out.n58 tank_out.n57 0.044
R2242 tank_out.n88 tank_out.n87 0.044
R2243 tank_out.n118 tank_out.n117 0.044
R2244 tank_out.n148 tank_out.n147 0.044
R2245 tank_out.n178 tank_out.n177 0.044
R2246 tank_out.n208 tank_out.n207 0.044
R2247 tank_out.n455 tank_out.n454 0.042
R2248 tank_out.n425 tank_out.n424 0.042
R2249 tank_out.n395 tank_out.n394 0.042
R2250 tank_out.n365 tank_out.n364 0.042
R2251 tank_out.n335 tank_out.n334 0.042
R2252 tank_out.n305 tank_out.n304 0.042
R2253 tank_out.n275 tank_out.n274 0.042
R2254 tank_out.n245 tank_out.n244 0.042
R2255 tank_out.n29 tank_out.n28 0.042
R2256 tank_out.n59 tank_out.n58 0.042
R2257 tank_out.n89 tank_out.n88 0.042
R2258 tank_out.n119 tank_out.n118 0.042
R2259 tank_out.n149 tank_out.n148 0.042
R2260 tank_out.n179 tank_out.n178 0.042
R2261 tank_out.n209 tank_out.n208 0.042
R2262 tank_out.n442 tank_out.n438 0.041
R2263 tank_out.n451 tank_out.n450 0.041
R2264 tank_out.n412 tank_out.n408 0.041
R2265 tank_out.n421 tank_out.n420 0.041
R2266 tank_out.n382 tank_out.n378 0.041
R2267 tank_out.n391 tank_out.n390 0.041
R2268 tank_out.n352 tank_out.n348 0.041
R2269 tank_out.n361 tank_out.n360 0.041
R2270 tank_out.n322 tank_out.n318 0.041
R2271 tank_out.n331 tank_out.n330 0.041
R2272 tank_out.n292 tank_out.n288 0.041
R2273 tank_out.n301 tank_out.n300 0.041
R2274 tank_out.n262 tank_out.n258 0.041
R2275 tank_out.n271 tank_out.n270 0.041
R2276 tank_out.n232 tank_out.n228 0.041
R2277 tank_out.n241 tank_out.n240 0.041
R2278 tank_out.n16 tank_out.n12 0.041
R2279 tank_out.n25 tank_out.n24 0.041
R2280 tank_out.n46 tank_out.n42 0.041
R2281 tank_out.n55 tank_out.n54 0.041
R2282 tank_out.n76 tank_out.n72 0.041
R2283 tank_out.n85 tank_out.n84 0.041
R2284 tank_out.n106 tank_out.n102 0.041
R2285 tank_out.n115 tank_out.n114 0.041
R2286 tank_out.n136 tank_out.n132 0.041
R2287 tank_out.n145 tank_out.n144 0.041
R2288 tank_out.n166 tank_out.n162 0.041
R2289 tank_out.n175 tank_out.n174 0.041
R2290 tank_out.n196 tank_out.n192 0.041
R2291 tank_out.n205 tank_out.n204 0.041
R2292 tank_out.n437 tank_out.n436 0.039
R2293 tank_out.n453 tank_out.n452 0.039
R2294 tank_out.n407 tank_out.n406 0.039
R2295 tank_out.n423 tank_out.n422 0.039
R2296 tank_out.n377 tank_out.n376 0.039
R2297 tank_out.n393 tank_out.n392 0.039
R2298 tank_out.n347 tank_out.n346 0.039
R2299 tank_out.n363 tank_out.n362 0.039
R2300 tank_out.n317 tank_out.n316 0.039
R2301 tank_out.n333 tank_out.n332 0.039
R2302 tank_out.n287 tank_out.n286 0.039
R2303 tank_out.n303 tank_out.n302 0.039
R2304 tank_out.n257 tank_out.n256 0.039
R2305 tank_out.n273 tank_out.n272 0.039
R2306 tank_out.n227 tank_out.n226 0.039
R2307 tank_out.n243 tank_out.n242 0.039
R2308 tank_out.n11 tank_out.n10 0.039
R2309 tank_out.n27 tank_out.n26 0.039
R2310 tank_out.n41 tank_out.n40 0.039
R2311 tank_out.n57 tank_out.n56 0.039
R2312 tank_out.n71 tank_out.n70 0.039
R2313 tank_out.n87 tank_out.n86 0.039
R2314 tank_out.n101 tank_out.n100 0.039
R2315 tank_out.n117 tank_out.n116 0.039
R2316 tank_out.n131 tank_out.n130 0.039
R2317 tank_out.n147 tank_out.n146 0.039
R2318 tank_out.n161 tank_out.n160 0.039
R2319 tank_out.n177 tank_out.n176 0.039
R2320 tank_out.n191 tank_out.n190 0.039
R2321 tank_out.n207 tank_out.n206 0.039
R2322 tank_out.n211 tank_out.n210 0.026
R2323 tank_out.n212 tank_out.n211 0.026
R2324 tank_out.n213 tank_out.n212 0.026
R2325 tank_out.n214 tank_out.n213 0.026
R2326 tank_out.n215 tank_out.n214 0.026
R2327 tank_out.n462 tank_out.n215 0.026
R2328 tank_out.n462 tank_out.n461 0.026
R2329 tank_out.n461 tank_out.n460 0.026
R2330 tank_out.n460 tank_out.n459 0.026
R2331 tank_out.n459 tank_out.n458 0.026
R2332 tank_out.n458 tank_out.n457 0.026
R2333 tank_out.n457 tank_out.n456 0.026
R2334 tank_out.n448 tank_out.n444 0.023
R2335 tank_out.n418 tank_out.n414 0.023
R2336 tank_out.n388 tank_out.n384 0.023
R2337 tank_out.n358 tank_out.n354 0.023
R2338 tank_out.n328 tank_out.n324 0.023
R2339 tank_out.n298 tank_out.n294 0.023
R2340 tank_out.n268 tank_out.n264 0.023
R2341 tank_out.n238 tank_out.n234 0.023
R2342 tank_out.n22 tank_out.n18 0.023
R2343 tank_out.n52 tank_out.n48 0.023
R2344 tank_out.n82 tank_out.n78 0.023
R2345 tank_out.n112 tank_out.n108 0.023
R2346 tank_out.n142 tank_out.n138 0.023
R2347 tank_out.n172 tank_out.n168 0.023
R2348 tank_out.n202 tank_out.n198 0.023
R2349 tank_out.n443 tank_out.n442 0.019
R2350 tank_out.n413 tank_out.n412 0.019
R2351 tank_out.n383 tank_out.n382 0.019
R2352 tank_out.n353 tank_out.n352 0.019
R2353 tank_out.n323 tank_out.n322 0.019
R2354 tank_out.n293 tank_out.n292 0.019
R2355 tank_out.n263 tank_out.n262 0.019
R2356 tank_out.n233 tank_out.n232 0.019
R2357 tank_out.n17 tank_out.n16 0.019
R2358 tank_out.n47 tank_out.n46 0.019
R2359 tank_out.n77 tank_out.n76 0.019
R2360 tank_out.n107 tank_out.n106 0.019
R2361 tank_out.n137 tank_out.n136 0.019
R2362 tank_out.n167 tank_out.n166 0.019
R2363 tank_out.n197 tank_out.n196 0.019
R2364 tank_out.n430 tank_out.n426 0.017
R2365 tank_out.n400 tank_out.n396 0.017
R2366 tank_out.n370 tank_out.n366 0.017
R2367 tank_out.n340 tank_out.n336 0.017
R2368 tank_out.n310 tank_out.n306 0.017
R2369 tank_out.n280 tank_out.n276 0.017
R2370 tank_out.n250 tank_out.n246 0.017
R2371 tank_out.n220 tank_out.n216 0.017
R2372 tank_out.n4 tank_out.n0 0.017
R2373 tank_out.n34 tank_out.n30 0.017
R2374 tank_out.n64 tank_out.n60 0.017
R2375 tank_out.n94 tank_out.n90 0.017
R2376 tank_out.n124 tank_out.n120 0.017
R2377 tank_out.n154 tank_out.n150 0.017
R2378 tank_out.n184 tank_out.n180 0.017
R2379 tank_out.n431 tank_out.n430 0.015
R2380 tank_out.n436 tank_out.n432 0.015
R2381 tank_out.n401 tank_out.n400 0.015
R2382 tank_out.n406 tank_out.n402 0.015
R2383 tank_out.n371 tank_out.n370 0.015
R2384 tank_out.n376 tank_out.n372 0.015
R2385 tank_out.n341 tank_out.n340 0.015
R2386 tank_out.n346 tank_out.n342 0.015
R2387 tank_out.n311 tank_out.n310 0.015
R2388 tank_out.n316 tank_out.n312 0.015
R2389 tank_out.n281 tank_out.n280 0.015
R2390 tank_out.n286 tank_out.n282 0.015
R2391 tank_out.n251 tank_out.n250 0.015
R2392 tank_out.n256 tank_out.n252 0.015
R2393 tank_out.n221 tank_out.n220 0.015
R2394 tank_out.n226 tank_out.n222 0.015
R2395 tank_out.n5 tank_out.n4 0.015
R2396 tank_out.n10 tank_out.n6 0.015
R2397 tank_out.n35 tank_out.n34 0.015
R2398 tank_out.n40 tank_out.n36 0.015
R2399 tank_out.n65 tank_out.n64 0.015
R2400 tank_out.n70 tank_out.n66 0.015
R2401 tank_out.n95 tank_out.n94 0.015
R2402 tank_out.n100 tank_out.n96 0.015
R2403 tank_out.n125 tank_out.n124 0.015
R2404 tank_out.n130 tank_out.n126 0.015
R2405 tank_out.n155 tank_out.n154 0.015
R2406 tank_out.n160 tank_out.n156 0.015
R2407 tank_out.n185 tank_out.n184 0.015
R2408 tank_out.n190 tank_out.n186 0.015
R2409 tank_out.n432 tank_out.n431 0.013
R2410 tank_out.n402 tank_out.n401 0.013
R2411 tank_out.n372 tank_out.n371 0.013
R2412 tank_out.n342 tank_out.n341 0.013
R2413 tank_out.n312 tank_out.n311 0.013
R2414 tank_out.n282 tank_out.n281 0.013
R2415 tank_out.n252 tank_out.n251 0.013
R2416 tank_out.n222 tank_out.n221 0.013
R2417 tank_out.n6 tank_out.n5 0.013
R2418 tank_out.n36 tank_out.n35 0.013
R2419 tank_out.n66 tank_out.n65 0.013
R2420 tank_out.n96 tank_out.n95 0.013
R2421 tank_out.n126 tank_out.n125 0.013
R2422 tank_out.n156 tank_out.n155 0.013
R2423 tank_out.n186 tank_out.n185 0.013
R2424 tank_out.n438 tank_out.n437 0.007
R2425 tank_out.n452 tank_out.n451 0.007
R2426 tank_out.n408 tank_out.n407 0.007
R2427 tank_out.n422 tank_out.n421 0.007
R2428 tank_out.n378 tank_out.n377 0.007
R2429 tank_out.n392 tank_out.n391 0.007
R2430 tank_out.n348 tank_out.n347 0.007
R2431 tank_out.n362 tank_out.n361 0.007
R2432 tank_out.n318 tank_out.n317 0.007
R2433 tank_out.n332 tank_out.n331 0.007
R2434 tank_out.n288 tank_out.n287 0.007
R2435 tank_out.n302 tank_out.n301 0.007
R2436 tank_out.n258 tank_out.n257 0.007
R2437 tank_out.n272 tank_out.n271 0.007
R2438 tank_out.n228 tank_out.n227 0.007
R2439 tank_out.n242 tank_out.n241 0.007
R2440 tank_out.n12 tank_out.n11 0.007
R2441 tank_out.n26 tank_out.n25 0.007
R2442 tank_out.n42 tank_out.n41 0.007
R2443 tank_out.n56 tank_out.n55 0.007
R2444 tank_out.n72 tank_out.n71 0.007
R2445 tank_out.n86 tank_out.n85 0.007
R2446 tank_out.n102 tank_out.n101 0.007
R2447 tank_out.n116 tank_out.n115 0.007
R2448 tank_out.n132 tank_out.n131 0.007
R2449 tank_out.n146 tank_out.n145 0.007
R2450 tank_out.n162 tank_out.n161 0.007
R2451 tank_out.n176 tank_out.n175 0.007
R2452 tank_out.n192 tank_out.n191 0.007
R2453 tank_out.n206 tank_out.n205 0.007
R2454 tank_out.n449 tank_out.n448 0.003
R2455 tank_out.n419 tank_out.n418 0.003
R2456 tank_out.n389 tank_out.n388 0.003
R2457 tank_out.n359 tank_out.n358 0.003
R2458 tank_out.n329 tank_out.n328 0.003
R2459 tank_out.n299 tank_out.n298 0.003
R2460 tank_out.n269 tank_out.n268 0.003
R2461 tank_out.n239 tank_out.n238 0.003
R2462 tank_out.n23 tank_out.n22 0.003
R2463 tank_out.n53 tank_out.n52 0.003
R2464 tank_out.n83 tank_out.n82 0.003
R2465 tank_out.n113 tank_out.n112 0.003
R2466 tank_out.n143 tank_out.n142 0.003
R2467 tank_out.n173 tank_out.n172 0.003
R2468 tank_out.n203 tank_out.n202 0.003
R2469 tank_out tank_out.n462 0.002
R2470 tank_out.n444 tank_out.n443 0.001
R2471 tank_out.n414 tank_out.n413 0.001
R2472 tank_out.n384 tank_out.n383 0.001
R2473 tank_out.n354 tank_out.n353 0.001
R2474 tank_out.n324 tank_out.n323 0.001
R2475 tank_out.n294 tank_out.n293 0.001
R2476 tank_out.n264 tank_out.n263 0.001
R2477 tank_out.n234 tank_out.n233 0.001
R2478 tank_out.n18 tank_out.n17 0.001
R2479 tank_out.n48 tank_out.n47 0.001
R2480 tank_out.n78 tank_out.n77 0.001
R2481 tank_out.n108 tank_out.n107 0.001
R2482 tank_out.n138 tank_out.n137 0.001
R2483 tank_out.n168 tank_out.n167 0.001
R2484 tank_out.n198 tank_out.n197 0.001
C6 source bulk 12.96185fF
C7 bias1_input bulk 15.02466fF
C8 tank_out bulk 11.96716fF
C9 bias2 bulk 8.51594fF
C10 tank_out.n0 bulk 0.01068fF
C11 tank_out.n1 bulk 0.00586fF
C12 tank_out.n2 bulk 0.00082fF
C13 tank_out.n3 bulk 0.00093fF
C14 tank_out.n4 bulk 0.00174fF
C15 tank_out.n5 bulk 0.00154fF
C16 tank_out.n6 bulk 0.00154fF
C17 tank_out.n7 bulk 0.00082fF
C18 tank_out.n8 bulk 0.00245fF
C19 tank_out.n9 bulk 0.00153fF
C20 tank_out.n10 bulk 0.00287fF
C21 tank_out.n11 bulk 0.00246fF
C22 tank_out.n12 bulk 0.00256fF
C23 tank_out.n13 bulk 0.00071fF
C24 tank_out.n14 bulk 0.00060fF
C25 tank_out.n15 bulk 0.00191fF
C26 tank_out.n16 bulk 0.00318fF
C27 tank_out.n17 bulk 0.00113fF
C28 tank_out.n18 bulk 0.00133fF
C29 tank_out.t25 bulk 0.01058fF 
C30 tank_out.t21 bulk 0.01058fF 
C31 tank_out.n19 bulk 0.02175fF
C32 tank_out.n20 bulk 0.00559fF
C33 tank_out.n21 bulk 0.00087fF
C34 tank_out.n22 bulk 0.00164fF
C35 tank_out.n23 bulk 0.01088fF
C36 tank_out.n24 bulk 0.01690fF
C37 tank_out.n25 bulk 0.00256fF
C38 tank_out.n26 bulk 0.00246fF
C39 tank_out.n27 bulk 0.00441fF
C40 tank_out.n28 bulk 0.00467fF
C41 tank_out.n29 bulk 0.01349fF
C42 tank_out.n30 bulk 0.01068fF
C43 tank_out.n31 bulk 0.00586fF
C44 tank_out.n32 bulk 0.00082fF
C45 tank_out.n33 bulk 0.00093fF
C46 tank_out.n34 bulk 0.00174fF
C47 tank_out.n35 bulk 0.00154fF
C48 tank_out.n36 bulk 0.00154fF
C49 tank_out.n37 bulk 0.00082fF
C50 tank_out.n38 bulk 0.00245fF
C51 tank_out.n39 bulk 0.00153fF
C52 tank_out.n40 bulk 0.00287fF
C53 tank_out.n41 bulk 0.00246fF
C54 tank_out.n42 bulk 0.00256fF
C55 tank_out.n43 bulk 0.00071fF
C56 tank_out.n44 bulk 0.00060fF
C57 tank_out.n45 bulk 0.00191fF
C58 tank_out.n46 bulk 0.00318fF
C59 tank_out.n47 bulk 0.00113fF
C60 tank_out.n48 bulk 0.00133fF
C61 tank_out.t22 bulk 0.01058fF 
C62 tank_out.t20 bulk 0.01058fF 
C63 tank_out.n49 bulk 0.02175fF
C64 tank_out.n50 bulk 0.00559fF
C65 tank_out.n51 bulk 0.00087fF
C66 tank_out.n52 bulk 0.00164fF
C67 tank_out.n53 bulk 0.01088fF
C68 tank_out.n54 bulk 0.01690fF
C69 tank_out.n55 bulk 0.00256fF
C70 tank_out.n56 bulk 0.00246fF
C71 tank_out.n57 bulk 0.00441fF
C72 tank_out.n58 bulk 0.00467fF
C73 tank_out.n59 bulk 0.01349fF
C74 tank_out.n60 bulk 0.01068fF
C75 tank_out.n61 bulk 0.00586fF
C76 tank_out.n62 bulk 0.00082fF
C77 tank_out.n63 bulk 0.00093fF
C78 tank_out.n64 bulk 0.00174fF
C79 tank_out.n65 bulk 0.00154fF
C80 tank_out.n66 bulk 0.00154fF
C81 tank_out.n67 bulk 0.00082fF
C82 tank_out.n68 bulk 0.00245fF
C83 tank_out.n69 bulk 0.00153fF
C84 tank_out.n70 bulk 0.00287fF
C85 tank_out.n71 bulk 0.00246fF
C86 tank_out.n72 bulk 0.00256fF
C87 tank_out.n73 bulk 0.00071fF
C88 tank_out.n74 bulk 0.00060fF
C89 tank_out.n75 bulk 0.00191fF
C90 tank_out.n76 bulk 0.00318fF
C91 tank_out.n77 bulk 0.00113fF
C92 tank_out.n78 bulk 0.00133fF
C93 tank_out.t5 bulk 0.01058fF 
C94 tank_out.t26 bulk 0.01058fF 
C95 tank_out.n79 bulk 0.02175fF
C96 tank_out.n80 bulk 0.00559fF
C97 tank_out.n81 bulk 0.00087fF
C98 tank_out.n82 bulk 0.00164fF
C99 tank_out.n83 bulk 0.01088fF
C100 tank_out.n84 bulk 0.01690fF
C101 tank_out.n85 bulk 0.00256fF
C102 tank_out.n86 bulk 0.00246fF
C103 tank_out.n87 bulk 0.00441fF
C104 tank_out.n88 bulk 0.00467fF
C105 tank_out.n89 bulk 0.01349fF
C106 tank_out.n90 bulk 0.01068fF
C107 tank_out.n91 bulk 0.00586fF
C108 tank_out.n92 bulk 0.00082fF
C109 tank_out.n93 bulk 0.00093fF
C110 tank_out.n94 bulk 0.00174fF
C111 tank_out.n95 bulk 0.00154fF
C112 tank_out.n96 bulk 0.00154fF
C113 tank_out.n97 bulk 0.00082fF
C114 tank_out.n98 bulk 0.00245fF
C115 tank_out.n99 bulk 0.00153fF
C116 tank_out.n100 bulk 0.00287fF
C117 tank_out.n101 bulk 0.00246fF
C118 tank_out.n102 bulk 0.00256fF
C119 tank_out.n103 bulk 0.00071fF
C120 tank_out.n104 bulk 0.00060fF
C121 tank_out.n105 bulk 0.00191fF
C122 tank_out.n106 bulk 0.00318fF
C123 tank_out.n107 bulk 0.00113fF
C124 tank_out.n108 bulk 0.00133fF
C125 tank_out.t1 bulk 0.01058fF 
C126 tank_out.t6 bulk 0.01058fF 
C127 tank_out.n109 bulk 0.02175fF
C128 tank_out.n110 bulk 0.00559fF
C129 tank_out.n111 bulk 0.00087fF
C130 tank_out.n112 bulk 0.00164fF
C131 tank_out.n113 bulk 0.01088fF
C132 tank_out.n114 bulk 0.01690fF
C133 tank_out.n115 bulk 0.00256fF
C134 tank_out.n116 bulk 0.00246fF
C135 tank_out.n117 bulk 0.00441fF
C136 tank_out.n118 bulk 0.00467fF
C137 tank_out.n119 bulk 0.01349fF
C138 tank_out.n120 bulk 0.01068fF
C139 tank_out.n121 bulk 0.00586fF
C140 tank_out.n122 bulk 0.00082fF
C141 tank_out.n123 bulk 0.00093fF
C142 tank_out.n124 bulk 0.00174fF
C143 tank_out.n125 bulk 0.00154fF
C144 tank_out.n126 bulk 0.00154fF
C145 tank_out.n127 bulk 0.00082fF
C146 tank_out.n128 bulk 0.00245fF
C147 tank_out.n129 bulk 0.00153fF
C148 tank_out.n130 bulk 0.00287fF
C149 tank_out.n131 bulk 0.00246fF
C150 tank_out.n132 bulk 0.00256fF
C151 tank_out.n133 bulk 0.00071fF
C152 tank_out.n134 bulk 0.00060fF
C153 tank_out.n135 bulk 0.00191fF
C154 tank_out.n136 bulk 0.00318fF
C155 tank_out.n137 bulk 0.00113fF
C156 tank_out.n138 bulk 0.00133fF
C157 tank_out.t7 bulk 0.01058fF 
C158 tank_out.t3 bulk 0.01058fF 
C159 tank_out.n139 bulk 0.02175fF
C160 tank_out.n140 bulk 0.00559fF
C161 tank_out.n141 bulk 0.00087fF
C162 tank_out.n142 bulk 0.00164fF
C163 tank_out.n143 bulk 0.01088fF
C164 tank_out.n144 bulk 0.01690fF
C165 tank_out.n145 bulk 0.00256fF
C166 tank_out.n146 bulk 0.00246fF
C167 tank_out.n147 bulk 0.00441fF
C168 tank_out.n148 bulk 0.00467fF
C169 tank_out.n149 bulk 0.01349fF
C170 tank_out.n150 bulk 0.01068fF
C171 tank_out.n151 bulk 0.00586fF
C172 tank_out.n152 bulk 0.00082fF
C173 tank_out.n153 bulk 0.00093fF
C174 tank_out.n154 bulk 0.00174fF
C175 tank_out.n155 bulk 0.00154fF
C176 tank_out.n156 bulk 0.00154fF
C177 tank_out.n157 bulk 0.00082fF
C178 tank_out.n158 bulk 0.00245fF
C179 tank_out.n159 bulk 0.00153fF
C180 tank_out.n160 bulk 0.00287fF
C181 tank_out.n161 bulk 0.00246fF
C182 tank_out.n162 bulk 0.00256fF
C183 tank_out.n163 bulk 0.00071fF
C184 tank_out.n164 bulk 0.00060fF
C185 tank_out.n165 bulk 0.00191fF
C186 tank_out.n166 bulk 0.00318fF
C187 tank_out.n167 bulk 0.00113fF
C188 tank_out.n168 bulk 0.00133fF
C189 tank_out.t4 bulk 0.01058fF 
C190 tank_out.t2 bulk 0.01058fF 
C191 tank_out.n169 bulk 0.02175fF
C192 tank_out.n170 bulk 0.00559fF
C193 tank_out.n171 bulk 0.00087fF
C194 tank_out.n172 bulk 0.00164fF
C195 tank_out.n173 bulk 0.01088fF
C196 tank_out.n174 bulk 0.01690fF
C197 tank_out.n175 bulk 0.00256fF
C198 tank_out.n176 bulk 0.00246fF
C199 tank_out.n177 bulk 0.00441fF
C200 tank_out.n178 bulk 0.00467fF
C201 tank_out.n179 bulk 0.01349fF
C202 tank_out.n180 bulk 0.01068fF
C203 tank_out.n181 bulk 0.00586fF
C204 tank_out.n182 bulk 0.00082fF
C205 tank_out.n183 bulk 0.00093fF
C206 tank_out.n184 bulk 0.00174fF
C207 tank_out.n185 bulk 0.00154fF
C208 tank_out.n186 bulk 0.00154fF
C209 tank_out.n187 bulk 0.00082fF
C210 tank_out.n188 bulk 0.00245fF
C211 tank_out.n189 bulk 0.00153fF
C212 tank_out.n190 bulk 0.00287fF
C213 tank_out.n191 bulk 0.00246fF
C214 tank_out.n192 bulk 0.00256fF
C215 tank_out.n193 bulk 0.00071fF
C216 tank_out.n194 bulk 0.00060fF
C217 tank_out.n195 bulk 0.00191fF
C218 tank_out.n196 bulk 0.00318fF
C219 tank_out.n197 bulk 0.00113fF
C220 tank_out.n198 bulk 0.00133fF
C221 tank_out.t0 bulk 0.01058fF 
C222 tank_out.n199 bulk 0.02977fF
C223 tank_out.n200 bulk 0.00559fF
C224 tank_out.n201 bulk 0.00087fF
C225 tank_out.n202 bulk 0.00164fF
C226 tank_out.n203 bulk 0.01088fF
C227 tank_out.n204 bulk 0.01690fF
C228 tank_out.n205 bulk 0.00256fF
C229 tank_out.n206 bulk 0.00246fF
C230 tank_out.n207 bulk 0.00441fF
C231 tank_out.n208 bulk 0.00467fF
C232 tank_out.n209 bulk 0.05393fF
C233 tank_out.n210 bulk 0.89506fF
C234 tank_out.n211 bulk 0.55903fF
C235 tank_out.n212 bulk 0.55903fF
C236 tank_out.n213 bulk 0.55903fF
C237 tank_out.n214 bulk 0.55903fF
C238 tank_out.n215 bulk 0.55476fF
C239 tank_out.n216 bulk 0.01068fF
C240 tank_out.n217 bulk 0.00586fF
C241 tank_out.n218 bulk 0.00082fF
C242 tank_out.n219 bulk 0.00093fF
C243 tank_out.n220 bulk 0.00174fF
C244 tank_out.n221 bulk 0.00154fF
C245 tank_out.n222 bulk 0.00154fF
C246 tank_out.n223 bulk 0.00082fF
C247 tank_out.n224 bulk 0.00245fF
C248 tank_out.n225 bulk 0.00153fF
C249 tank_out.n226 bulk 0.00287fF
C250 tank_out.n227 bulk 0.00246fF
C251 tank_out.n228 bulk 0.00256fF
C252 tank_out.n229 bulk 0.00071fF
C253 tank_out.n230 bulk 0.00060fF
C254 tank_out.n231 bulk 0.00191fF
C255 tank_out.n232 bulk 0.00318fF
C256 tank_out.n233 bulk 0.00113fF
C257 tank_out.n234 bulk 0.00133fF
C258 tank_out.t27 bulk 0.01058fF 
C259 tank_out.t24 bulk 0.01058fF 
C260 tank_out.n235 bulk 0.02175fF
C261 tank_out.n236 bulk 0.00559fF
C262 tank_out.n237 bulk 0.00087fF
C263 tank_out.n238 bulk 0.00164fF
C264 tank_out.n239 bulk 0.01088fF
C265 tank_out.n240 bulk 0.01690fF
C266 tank_out.n241 bulk 0.00256fF
C267 tank_out.n242 bulk 0.00246fF
C268 tank_out.n243 bulk 0.00441fF
C269 tank_out.n244 bulk 0.00467fF
C270 tank_out.n245 bulk 0.01349fF
C271 tank_out.n246 bulk 0.01068fF
C272 tank_out.n247 bulk 0.00586fF
C273 tank_out.n248 bulk 0.00082fF
C274 tank_out.n249 bulk 0.00093fF
C275 tank_out.n250 bulk 0.00174fF
C276 tank_out.n251 bulk 0.00154fF
C277 tank_out.n252 bulk 0.00154fF
C278 tank_out.n253 bulk 0.00082fF
C279 tank_out.n254 bulk 0.00245fF
C280 tank_out.n255 bulk 0.00153fF
C281 tank_out.n256 bulk 0.00287fF
C282 tank_out.n257 bulk 0.00246fF
C283 tank_out.n258 bulk 0.00256fF
C284 tank_out.n259 bulk 0.00071fF
C285 tank_out.n260 bulk 0.00060fF
C286 tank_out.n261 bulk 0.00191fF
C287 tank_out.n262 bulk 0.00318fF
C288 tank_out.n263 bulk 0.00113fF
C289 tank_out.n264 bulk 0.00133fF
C290 tank_out.t23 bulk 0.01058fF 
C291 tank_out.t9 bulk 0.01058fF 
C292 tank_out.n265 bulk 0.02175fF
C293 tank_out.n266 bulk 0.00559fF
C294 tank_out.n267 bulk 0.00087fF
C295 tank_out.n268 bulk 0.00164fF
C296 tank_out.n269 bulk 0.01088fF
C297 tank_out.n270 bulk 0.01690fF
C298 tank_out.n271 bulk 0.00256fF
C299 tank_out.n272 bulk 0.00246fF
C300 tank_out.n273 bulk 0.00441fF
C301 tank_out.n274 bulk 0.00467fF
C302 tank_out.n275 bulk 0.01349fF
C303 tank_out.n276 bulk 0.01068fF
C304 tank_out.n277 bulk 0.00586fF
C305 tank_out.n278 bulk 0.00082fF
C306 tank_out.n279 bulk 0.00093fF
C307 tank_out.n280 bulk 0.00174fF
C308 tank_out.n281 bulk 0.00154fF
C309 tank_out.n282 bulk 0.00154fF
C310 tank_out.n283 bulk 0.00082fF
C311 tank_out.n284 bulk 0.00245fF
C312 tank_out.n285 bulk 0.00153fF
C313 tank_out.n286 bulk 0.00287fF
C314 tank_out.n287 bulk 0.00246fF
C315 tank_out.n288 bulk 0.00256fF
C316 tank_out.n289 bulk 0.00071fF
C317 tank_out.n290 bulk 0.00060fF
C318 tank_out.n291 bulk 0.00191fF
C319 tank_out.n292 bulk 0.00318fF
C320 tank_out.n293 bulk 0.00113fF
C321 tank_out.n294 bulk 0.00133fF
C322 tank_out.t8 bulk 0.01058fF 
C323 tank_out.t10 bulk 0.01058fF 
C324 tank_out.n295 bulk 0.02175fF
C325 tank_out.n296 bulk 0.00559fF
C326 tank_out.n297 bulk 0.00087fF
C327 tank_out.n298 bulk 0.00164fF
C328 tank_out.n299 bulk 0.01088fF
C329 tank_out.n300 bulk 0.01690fF
C330 tank_out.n301 bulk 0.00256fF
C331 tank_out.n302 bulk 0.00246fF
C332 tank_out.n303 bulk 0.00441fF
C333 tank_out.n304 bulk 0.00467fF
C334 tank_out.n305 bulk 0.01349fF
C335 tank_out.n306 bulk 0.01068fF
C336 tank_out.n307 bulk 0.00586fF
C337 tank_out.n308 bulk 0.00082fF
C338 tank_out.n309 bulk 0.00093fF
C339 tank_out.n310 bulk 0.00174fF
C340 tank_out.n311 bulk 0.00154fF
C341 tank_out.n312 bulk 0.00154fF
C342 tank_out.n313 bulk 0.00082fF
C343 tank_out.n314 bulk 0.00245fF
C344 tank_out.n315 bulk 0.00153fF
C345 tank_out.n316 bulk 0.00287fF
C346 tank_out.n317 bulk 0.00246fF
C347 tank_out.n318 bulk 0.00256fF
C348 tank_out.n319 bulk 0.00071fF
C349 tank_out.n320 bulk 0.00060fF
C350 tank_out.n321 bulk 0.00191fF
C351 tank_out.n322 bulk 0.00318fF
C352 tank_out.n323 bulk 0.00113fF
C353 tank_out.n324 bulk 0.00133fF
C354 tank_out.t14 bulk 0.01058fF 
C355 tank_out.t11 bulk 0.01058fF 
C356 tank_out.n325 bulk 0.02175fF
C357 tank_out.n326 bulk 0.00559fF
C358 tank_out.n327 bulk 0.00087fF
C359 tank_out.n328 bulk 0.00164fF
C360 tank_out.n329 bulk 0.01088fF
C361 tank_out.n330 bulk 0.01690fF
C362 tank_out.n331 bulk 0.00256fF
C363 tank_out.n332 bulk 0.00246fF
C364 tank_out.n333 bulk 0.00441fF
C365 tank_out.n334 bulk 0.00467fF
C366 tank_out.n335 bulk 0.01349fF
C367 tank_out.n336 bulk 0.01068fF
C368 tank_out.n337 bulk 0.00586fF
C369 tank_out.n338 bulk 0.00082fF
C370 tank_out.n339 bulk 0.00093fF
C371 tank_out.n340 bulk 0.00174fF
C372 tank_out.n341 bulk 0.00154fF
C373 tank_out.n342 bulk 0.00154fF
C374 tank_out.n343 bulk 0.00082fF
C375 tank_out.n344 bulk 0.00245fF
C376 tank_out.n345 bulk 0.00153fF
C377 tank_out.n346 bulk 0.00287fF
C378 tank_out.n347 bulk 0.00246fF
C379 tank_out.n348 bulk 0.00256fF
C380 tank_out.n349 bulk 0.00071fF
C381 tank_out.n350 bulk 0.00060fF
C382 tank_out.n351 bulk 0.00191fF
C383 tank_out.n352 bulk 0.00318fF
C384 tank_out.n353 bulk 0.00113fF
C385 tank_out.n354 bulk 0.00133fF
C386 tank_out.t17 bulk 0.01058fF 
C387 tank_out.t13 bulk 0.01058fF 
C388 tank_out.n355 bulk 0.02175fF
C389 tank_out.n356 bulk 0.00559fF
C390 tank_out.n357 bulk 0.00087fF
C391 tank_out.n358 bulk 0.00164fF
C392 tank_out.n359 bulk 0.01088fF
C393 tank_out.n360 bulk 0.01690fF
C394 tank_out.n361 bulk 0.00256fF
C395 tank_out.n362 bulk 0.00246fF
C396 tank_out.n363 bulk 0.00441fF
C397 tank_out.n364 bulk 0.00467fF
C398 tank_out.n365 bulk 0.01349fF
C399 tank_out.n366 bulk 0.01068fF
C400 tank_out.n367 bulk 0.00586fF
C401 tank_out.n368 bulk 0.00082fF
C402 tank_out.n369 bulk 0.00093fF
C403 tank_out.n370 bulk 0.00174fF
C404 tank_out.n371 bulk 0.00154fF
C405 tank_out.n372 bulk 0.00154fF
C406 tank_out.n373 bulk 0.00082fF
C407 tank_out.n374 bulk 0.00245fF
C408 tank_out.n375 bulk 0.00153fF
C409 tank_out.n376 bulk 0.00287fF
C410 tank_out.n377 bulk 0.00246fF
C411 tank_out.n378 bulk 0.00256fF
C412 tank_out.n379 bulk 0.00071fF
C413 tank_out.n380 bulk 0.00060fF
C414 tank_out.n381 bulk 0.00191fF
C415 tank_out.n382 bulk 0.00318fF
C416 tank_out.n383 bulk 0.00113fF
C417 tank_out.n384 bulk 0.00133fF
C418 tank_out.t19 bulk 0.01058fF 
C419 tank_out.t16 bulk 0.01058fF 
C420 tank_out.n385 bulk 0.02175fF
C421 tank_out.n386 bulk 0.00559fF
C422 tank_out.n387 bulk 0.00087fF
C423 tank_out.n388 bulk 0.00164fF
C424 tank_out.n389 bulk 0.01088fF
C425 tank_out.n390 bulk 0.01690fF
C426 tank_out.n391 bulk 0.00256fF
C427 tank_out.n392 bulk 0.00246fF
C428 tank_out.n393 bulk 0.00441fF
C429 tank_out.n394 bulk 0.00467fF
C430 tank_out.n395 bulk 0.01349fF
C431 tank_out.n396 bulk 0.01068fF
C432 tank_out.n397 bulk 0.00586fF
C433 tank_out.n398 bulk 0.00082fF
C434 tank_out.n399 bulk 0.00093fF
C435 tank_out.n400 bulk 0.00174fF
C436 tank_out.n401 bulk 0.00154fF
C437 tank_out.n402 bulk 0.00154fF
C438 tank_out.n403 bulk 0.00082fF
C439 tank_out.n404 bulk 0.00245fF
C440 tank_out.n405 bulk 0.00153fF
C441 tank_out.n406 bulk 0.00287fF
C442 tank_out.n407 bulk 0.00246fF
C443 tank_out.n408 bulk 0.00256fF
C444 tank_out.n409 bulk 0.00071fF
C445 tank_out.n410 bulk 0.00060fF
C446 tank_out.n411 bulk 0.00191fF
C447 tank_out.n412 bulk 0.00318fF
C448 tank_out.n413 bulk 0.00113fF
C449 tank_out.n414 bulk 0.00133fF
C450 tank_out.t12 bulk 0.01058fF 
C451 tank_out.t18 bulk 0.01058fF 
C452 tank_out.n415 bulk 0.02175fF
C453 tank_out.n416 bulk 0.00559fF
C454 tank_out.n417 bulk 0.00087fF
C455 tank_out.n418 bulk 0.00164fF
C456 tank_out.n419 bulk 0.01088fF
C457 tank_out.n420 bulk 0.01690fF
C458 tank_out.n421 bulk 0.00256fF
C459 tank_out.n422 bulk 0.00246fF
C460 tank_out.n423 bulk 0.00441fF
C461 tank_out.n424 bulk 0.00467fF
C462 tank_out.n425 bulk 0.01349fF
C463 tank_out.n426 bulk 0.01068fF
C464 tank_out.n427 bulk 0.00586fF
C465 tank_out.n428 bulk 0.00082fF
C466 tank_out.n429 bulk 0.00093fF
C467 tank_out.n430 bulk 0.00174fF
C468 tank_out.n431 bulk 0.00154fF
C469 tank_out.n432 bulk 0.00154fF
C470 tank_out.n433 bulk 0.00082fF
C471 tank_out.n434 bulk 0.00245fF
C472 tank_out.n435 bulk 0.00153fF
C473 tank_out.n436 bulk 0.00287fF
C474 tank_out.n437 bulk 0.00246fF
C475 tank_out.n438 bulk 0.00256fF
C476 tank_out.n439 bulk 0.00071fF
C477 tank_out.n440 bulk 0.00060fF
C478 tank_out.n441 bulk 0.00191fF
C479 tank_out.n442 bulk 0.00318fF
C480 tank_out.n443 bulk 0.00113fF
C481 tank_out.n444 bulk 0.00133fF
C482 tank_out.t15 bulk 0.01058fF 
C483 tank_out.n445 bulk 0.02977fF
C484 tank_out.n446 bulk 0.00559fF
C485 tank_out.n447 bulk 0.00087fF
C486 tank_out.n448 bulk 0.00164fF
C487 tank_out.n449 bulk 0.01088fF
C488 tank_out.n450 bulk 0.01690fF
C489 tank_out.n451 bulk 0.00256fF
C490 tank_out.n452 bulk 0.00246fF
C491 tank_out.n453 bulk 0.00441fF
C492 tank_out.n454 bulk 0.00467fF
C493 tank_out.n455 bulk 0.05393fF
C494 tank_out.n456 bulk 0.89506fF
C495 tank_out.n457 bulk 0.55903fF
C496 tank_out.n458 bulk 0.55903fF
C497 tank_out.n459 bulk 0.55903fF
C498 tank_out.n460 bulk 0.55903fF
C499 tank_out.n461 bulk 0.55903fF
C500 tank_out.n462 bulk 17.33180fF
C501 bias2.t23 bulk 0.04736fF 
C502 bias2.n0 bulk 0.57751fF
C503 bias2.t20 bulk 0.04736fF 
C504 bias2.n1 bulk 0.28416fF
C505 bias2.t26 bulk 0.04736fF 
C506 bias2.n2 bulk 0.28416fF
C507 bias2.t22 bulk 0.04736fF 
C508 bias2.n3 bulk 0.28416fF
C509 bias2.t5 bulk 0.04736fF 
C510 bias2.n4 bulk 0.28416fF
C511 bias2.t2 bulk 0.04736fF 
C512 bias2.n5 bulk 0.28416fF
C513 bias2.t0 bulk 0.04736fF 
C514 bias2.n6 bulk 0.28416fF
C515 bias2.t4 bulk 0.04736fF 
C516 bias2.n7 bulk 0.28416fF
C517 bias2.t19 bulk 0.04736fF 
C518 bias2.n8 bulk 0.28416fF
C519 bias2.t13 bulk 0.04736fF 
C520 bias2.n9 bulk 0.28416fF
C521 bias2.t10 bulk 0.04736fF 
C522 bias2.n10 bulk 0.28416fF
C523 bias2.t8 bulk 0.04736fF 
C524 bias2.n11 bulk 0.28416fF
C525 bias2.t15 bulk 0.04736fF 
C526 bias2.n12 bulk 0.28416fF
C527 bias2.t12 bulk 0.04736fF 
C528 bias2.n13 bulk 0.27906fF
C529 bias2.t27 bulk 0.03953fF 
C530 bias2.n14 bulk 0.60030fF
C531 bias2.t25 bulk 0.03953fF 
C532 bias2.n15 bulk 0.29199fF
C533 bias2.t24 bulk 0.03953fF 
C534 bias2.n16 bulk 0.29199fF
C535 bias2.t21 bulk 0.03953fF 
C536 bias2.n17 bulk 0.29199fF
C537 bias2.t1 bulk 0.03953fF 
C538 bias2.n18 bulk 0.29199fF
C539 bias2.t7 bulk 0.03953fF 
C540 bias2.n19 bulk 0.29199fF
C541 bias2.t6 bulk 0.03953fF 
C542 bias2.n20 bulk 0.29199fF
C543 bias2.t3 bulk 0.03953fF 
C544 bias2.n21 bulk 0.29199fF
C545 bias2.t18 bulk 0.03953fF 
C546 bias2.n22 bulk 0.29199fF
C547 bias2.t17 bulk 0.03953fF 
C548 bias2.n23 bulk 0.29199fF
C549 bias2.t16 bulk 0.03953fF 
C550 bias2.n24 bulk 0.29199fF
C551 bias2.t14 bulk 0.03953fF 
C552 bias2.n25 bulk 0.29199fF
C553 bias2.t11 bulk 0.03953fF 
C554 bias2.n26 bulk 0.29199fF
C555 bias2.t9 bulk 0.03953fF 
C556 bias2.n27 bulk 0.33145fF
C557 bias2.n28 bulk 0.18480fF
C558 bias2.n29 bulk 0.03157fF
C559 bias2.n30 bulk 0.05942fF
C560 bias2.n31 bulk 0.05942fF
C561 bias2.n32 bulk 0.05942fF
C562 bias2.n33 bulk 0.03157fF
C563 bias2.n34 bulk 0.14016fF
C564 bias2.n35 bulk 0.05928fF
C565 bias2.n36 bulk 0.03817fF
C566 bias2.n37 bulk 0.03878fF
C567 bias2.n38 bulk 0.03878fF
C568 bias2.n39 bulk 0.03878fF
C569 bias2.n40 bulk 0.03878fF
C570 bias2.n41 bulk 0.03878fF
C571 bias2.n42 bulk 0.03878fF
C572 bias2.n43 bulk 0.03737fF
C573 bias2.n44 bulk 0.03878fF
C574 bias2.n45 bulk 0.04070fF
C575 bias2.n46 bulk 0.03825fF
C576 bias2.n47 bulk 0.14252fF
C577 bias2.n48 bulk 0.05849fF
C578 bias2.n49 bulk 0.05942fF
C579 bias2.n50 bulk 0.05942fF
C580 bias2.n51 bulk 0.05942fF
C581 bias2.n52 bulk 0.05942fF
C582 bias2.n53 bulk 0.05942fF
C583 bias2.n54 bulk 0.05942fF
C584 bias2.n55 bulk 0.05664fF
C585 bias2.n56 bulk 0.97100fF
C586 bias2.n57 bulk 0.05942fF
C587 bias2.n58 bulk 0.16742fF
C588 bias2.n59 bulk 0.09071fF
C589 bias2.n60 bulk 0.36985fF
C590 bias2.n61 bulk 1.94864fF
C591 source.n0 bulk 0.00595fF
C592 source.n1 bulk 0.00083fF
C593 source.n2 bulk 0.00094fF
C594 source.n3 bulk 0.00072fF
C595 source.n4 bulk 0.00061fF
C596 source.n5 bulk 0.00193fF
C597 source.t25 bulk 0.01072fF 
C598 source.t16 bulk 0.01072fF 
C599 source.n6 bulk 0.02204fF
C600 source.n7 bulk 0.00566fF
C601 source.n8 bulk 0.00088fF
C602 source.n9 bulk 0.01027fF
C603 source.n10 bulk 0.00166fF
C604 source.n11 bulk 0.00135fF
C605 source.n12 bulk 0.00114fF
C606 source.n13 bulk 0.00322fF
C607 source.n14 bulk 0.00260fF
C608 source.n15 bulk 0.00249fF
C609 source.n16 bulk 0.00083fF
C610 source.n17 bulk 0.00248fF
C611 source.n18 bulk 0.00155fF
C612 source.n19 bulk 0.00291fF
C613 source.n20 bulk 0.00156fF
C614 source.n21 bulk 0.00156fF
C615 source.n22 bulk 0.00177fF
C616 source.n23 bulk 0.01154fF
C617 source.n24 bulk 0.01641fF
C618 source.n25 bulk 0.00249fF
C619 source.n26 bulk 0.00260fF
C620 source.n27 bulk 0.00457fF
C621 source.n28 bulk 0.00483fF
C622 source.n29 bulk 0.02210fF
C623 source.n30 bulk 0.00595fF
C624 source.n31 bulk 0.00083fF
C625 source.n32 bulk 0.00094fF
C626 source.n33 bulk 0.00072fF
C627 source.n34 bulk 0.00061fF
C628 source.n35 bulk 0.00193fF
C629 source.t8 bulk 0.01072fF 
C630 source.t5 bulk 0.01072fF 
C631 source.n36 bulk 0.02204fF
C632 source.n37 bulk 0.00566fF
C633 source.n38 bulk 0.00088fF
C634 source.n39 bulk 0.01027fF
C635 source.n40 bulk 0.00166fF
C636 source.n41 bulk 0.00135fF
C637 source.n42 bulk 0.00114fF
C638 source.n43 bulk 0.00322fF
C639 source.n44 bulk 0.00260fF
C640 source.n45 bulk 0.00249fF
C641 source.n46 bulk 0.00083fF
C642 source.n47 bulk 0.00248fF
C643 source.n48 bulk 0.00155fF
C644 source.n49 bulk 0.00291fF
C645 source.n50 bulk 0.00156fF
C646 source.n51 bulk 0.00156fF
C647 source.n52 bulk 0.00177fF
C648 source.n53 bulk 0.01154fF
C649 source.n54 bulk 0.01641fF
C650 source.n55 bulk 0.00249fF
C651 source.n56 bulk 0.00260fF
C652 source.n57 bulk 0.00457fF
C653 source.n58 bulk 0.00483fF
C654 source.n59 bulk 0.02210fF
C655 source.n60 bulk 0.00595fF
C656 source.n61 bulk 0.00083fF
C657 source.n62 bulk 0.00094fF
C658 source.n63 bulk 0.00072fF
C659 source.n64 bulk 0.00061fF
C660 source.n65 bulk 0.00193fF
C661 source.t19 bulk 0.01072fF 
C662 source.t10 bulk 0.01072fF 
C663 source.n66 bulk 0.02204fF
C664 source.n67 bulk 0.00566fF
C665 source.n68 bulk 0.00088fF
C666 source.n69 bulk 0.01027fF
C667 source.n70 bulk 0.00166fF
C668 source.n71 bulk 0.00135fF
C669 source.n72 bulk 0.00114fF
C670 source.n73 bulk 0.00322fF
C671 source.n74 bulk 0.00260fF
C672 source.n75 bulk 0.00249fF
C673 source.n76 bulk 0.00083fF
C674 source.n77 bulk 0.00248fF
C675 source.n78 bulk 0.00155fF
C676 source.n79 bulk 0.00291fF
C677 source.n80 bulk 0.00156fF
C678 source.n81 bulk 0.00156fF
C679 source.n82 bulk 0.00177fF
C680 source.n83 bulk 0.01154fF
C681 source.n84 bulk 0.01641fF
C682 source.n85 bulk 0.00249fF
C683 source.n86 bulk 0.00260fF
C684 source.n87 bulk 0.00457fF
C685 source.n88 bulk 0.00483fF
C686 source.n89 bulk 0.02210fF
C687 source.n90 bulk 0.00595fF
C688 source.n91 bulk 0.00083fF
C689 source.n92 bulk 0.00094fF
C690 source.n93 bulk 0.00072fF
C691 source.n94 bulk 0.00061fF
C692 source.n95 bulk 0.00193fF
C693 source.t6 bulk 0.01072fF 
C694 source.t21 bulk 0.01072fF 
C695 source.n96 bulk 0.02204fF
C696 source.n97 bulk 0.00566fF
C697 source.n98 bulk 0.00088fF
C698 source.n99 bulk 0.01027fF
C699 source.n100 bulk 0.00166fF
C700 source.n101 bulk 0.00135fF
C701 source.n102 bulk 0.00114fF
C702 source.n103 bulk 0.00322fF
C703 source.n104 bulk 0.00260fF
C704 source.n105 bulk 0.00249fF
C705 source.n106 bulk 0.00083fF
C706 source.n107 bulk 0.00248fF
C707 source.n108 bulk 0.00155fF
C708 source.n109 bulk 0.00291fF
C709 source.n110 bulk 0.00156fF
C710 source.n111 bulk 0.00156fF
C711 source.n112 bulk 0.00177fF
C712 source.n113 bulk 0.01154fF
C713 source.n114 bulk 0.01641fF
C714 source.n115 bulk 0.00249fF
C715 source.n116 bulk 0.00260fF
C716 source.n117 bulk 0.00457fF
C717 source.n118 bulk 0.00483fF
C718 source.n119 bulk 0.02210fF
C719 source.n120 bulk 0.00595fF
C720 source.n121 bulk 0.00083fF
C721 source.n122 bulk 0.00094fF
C722 source.n123 bulk 0.00072fF
C723 source.n124 bulk 0.00061fF
C724 source.n125 bulk 0.00193fF
C725 source.t13 bulk 0.01072fF 
C726 source.t1 bulk 0.01072fF 
C727 source.n126 bulk 0.02204fF
C728 source.n127 bulk 0.00566fF
C729 source.n128 bulk 0.00088fF
C730 source.n129 bulk 0.01027fF
C731 source.n130 bulk 0.00166fF
C732 source.n131 bulk 0.00135fF
C733 source.n132 bulk 0.00114fF
C734 source.n133 bulk 0.00322fF
C735 source.n134 bulk 0.00260fF
C736 source.n135 bulk 0.00249fF
C737 source.n136 bulk 0.00083fF
C738 source.n137 bulk 0.00248fF
C739 source.n138 bulk 0.00155fF
C740 source.n139 bulk 0.00291fF
C741 source.n140 bulk 0.00156fF
C742 source.n141 bulk 0.00156fF
C743 source.n142 bulk 0.00177fF
C744 source.n143 bulk 0.01154fF
C745 source.n144 bulk 0.01641fF
C746 source.n145 bulk 0.00249fF
C747 source.n146 bulk 0.00260fF
C748 source.n147 bulk 0.00457fF
C749 source.n148 bulk 0.00483fF
C750 source.n149 bulk 0.02210fF
C751 source.n150 bulk 0.00595fF
C752 source.n151 bulk 0.00083fF
C753 source.n152 bulk 0.00094fF
C754 source.n153 bulk 0.00072fF
C755 source.n154 bulk 0.00061fF
C756 source.n155 bulk 0.00193fF
C757 source.t24 bulk 0.01072fF 
C758 source.t15 bulk 0.01072fF 
C759 source.n156 bulk 0.02204fF
C760 source.n157 bulk 0.00566fF
C761 source.n158 bulk 0.00088fF
C762 source.n159 bulk 0.01027fF
C763 source.n160 bulk 0.00166fF
C764 source.n161 bulk 0.00135fF
C765 source.n162 bulk 0.00114fF
C766 source.n163 bulk 0.00322fF
C767 source.n164 bulk 0.00260fF
C768 source.n165 bulk 0.00249fF
C769 source.n166 bulk 0.00083fF
C770 source.n167 bulk 0.00248fF
C771 source.n168 bulk 0.00155fF
C772 source.n169 bulk 0.00291fF
C773 source.n170 bulk 0.00156fF
C774 source.n171 bulk 0.00156fF
C775 source.n172 bulk 0.00177fF
C776 source.n173 bulk 0.01154fF
C777 source.n174 bulk 0.01641fF
C778 source.n175 bulk 0.00249fF
C779 source.n176 bulk 0.00260fF
C780 source.n177 bulk 0.00457fF
C781 source.n178 bulk 0.00483fF
C782 source.n179 bulk 0.02210fF
C783 source.n180 bulk 0.00072fF
C784 source.n181 bulk 0.00061fF
C785 source.n182 bulk 0.00193fF
C786 source.t3 bulk 0.01072fF 
C787 source.t26 bulk 0.01072fF 
C788 source.n183 bulk 0.02204fF
C789 source.n184 bulk 0.00566fF
C790 source.n185 bulk 0.00088fF
C791 source.n186 bulk 0.01027fF
C792 source.n187 bulk 0.00166fF
C793 source.n188 bulk 0.00135fF
C794 source.n189 bulk 0.00114fF
C795 source.n190 bulk 0.00322fF
C796 source.n191 bulk 0.00260fF
C797 source.n192 bulk 0.00249fF
C798 source.n193 bulk 0.00083fF
C799 source.n194 bulk 0.00248fF
C800 source.n195 bulk 0.00155fF
C801 source.n196 bulk 0.00291fF
C802 source.n197 bulk 0.00156fF
C803 source.n198 bulk 0.00156fF
C804 source.n199 bulk 0.00595fF
C805 source.n200 bulk 0.00083fF
C806 source.n201 bulk 0.00094fF
C807 source.n202 bulk 0.00177fF
C808 source.n203 bulk 0.01153fF
C809 source.n204 bulk 0.01641fF
C810 source.n205 bulk 0.00249fF
C811 source.n206 bulk 0.00260fF
C812 source.n207 bulk 0.00457fF
C813 source.n208 bulk 0.00483fF
C814 source.n209 bulk 0.05190fF
C815 source.n210 bulk 0.88512fF
C816 source.n211 bulk 0.51852fF
C817 source.n212 bulk 0.51852fF
C818 source.n213 bulk 0.51852fF
C819 source.n214 bulk 0.51852fF
C820 source.n215 bulk 0.39770fF
C821 source.n216 bulk 0.00595fF
C822 source.n217 bulk 0.00083fF
C823 source.n218 bulk 0.00094fF
C824 source.n219 bulk 0.00072fF
C825 source.n220 bulk 0.00061fF
C826 source.n221 bulk 0.00193fF
C827 source.t14 bulk 0.01072fF 
C828 source.t2 bulk 0.01072fF 
C829 source.n222 bulk 0.02204fF
C830 source.n223 bulk 0.00566fF
C831 source.n224 bulk 0.00088fF
C832 source.n225 bulk 0.01027fF
C833 source.n226 bulk 0.00166fF
C834 source.n227 bulk 0.00135fF
C835 source.n228 bulk 0.00114fF
C836 source.n229 bulk 0.00322fF
C837 source.n230 bulk 0.00260fF
C838 source.n231 bulk 0.00249fF
C839 source.n232 bulk 0.00083fF
C840 source.n233 bulk 0.00248fF
C841 source.n234 bulk 0.00155fF
C842 source.n235 bulk 0.00291fF
C843 source.n236 bulk 0.00156fF
C844 source.n237 bulk 0.00156fF
C845 source.n238 bulk 0.00177fF
C846 source.n239 bulk 0.01154fF
C847 source.n240 bulk 0.01641fF
C848 source.n241 bulk 0.00249fF
C849 source.n242 bulk 0.00260fF
C850 source.n243 bulk 0.00457fF
C851 source.n244 bulk 0.00483fF
C852 source.n245 bulk 0.02210fF
C853 source.n246 bulk 0.00595fF
C854 source.n247 bulk 0.00083fF
C855 source.n248 bulk 0.00094fF
C856 source.n249 bulk 0.00072fF
C857 source.n250 bulk 0.00061fF
C858 source.n251 bulk 0.00193fF
C859 source.t7 bulk 0.01072fF 
C860 source.t22 bulk 0.01072fF 
C861 source.n252 bulk 0.02204fF
C862 source.n253 bulk 0.00566fF
C863 source.n254 bulk 0.00088fF
C864 source.n255 bulk 0.01027fF
C865 source.n256 bulk 0.00166fF
C866 source.n257 bulk 0.00135fF
C867 source.n258 bulk 0.00114fF
C868 source.n259 bulk 0.00322fF
C869 source.n260 bulk 0.00260fF
C870 source.n261 bulk 0.00249fF
C871 source.n262 bulk 0.00083fF
C872 source.n263 bulk 0.00248fF
C873 source.n264 bulk 0.00155fF
C874 source.n265 bulk 0.00291fF
C875 source.n266 bulk 0.00156fF
C876 source.n267 bulk 0.00156fF
C877 source.n268 bulk 0.00177fF
C878 source.n269 bulk 0.01154fF
C879 source.n270 bulk 0.01641fF
C880 source.n271 bulk 0.00249fF
C881 source.n272 bulk 0.00260fF
C882 source.n273 bulk 0.00457fF
C883 source.n274 bulk 0.00483fF
C884 source.n275 bulk 0.02210fF
C885 source.n276 bulk 0.00595fF
C886 source.n277 bulk 0.00083fF
C887 source.n278 bulk 0.00094fF
C888 source.n279 bulk 0.00072fF
C889 source.n280 bulk 0.00061fF
C890 source.n281 bulk 0.00193fF
C891 source.t18 bulk 0.01072fF 
C892 source.t11 bulk 0.01072fF 
C893 source.n282 bulk 0.02204fF
C894 source.n283 bulk 0.00566fF
C895 source.n284 bulk 0.00088fF
C896 source.n285 bulk 0.01027fF
C897 source.n286 bulk 0.00166fF
C898 source.n287 bulk 0.00135fF
C899 source.n288 bulk 0.00114fF
C900 source.n289 bulk 0.00322fF
C901 source.n290 bulk 0.00260fF
C902 source.n291 bulk 0.00249fF
C903 source.n292 bulk 0.00083fF
C904 source.n293 bulk 0.00248fF
C905 source.n294 bulk 0.00155fF
C906 source.n295 bulk 0.00291fF
C907 source.n296 bulk 0.00156fF
C908 source.n297 bulk 0.00156fF
C909 source.n298 bulk 0.00177fF
C910 source.n299 bulk 0.01154fF
C911 source.n300 bulk 0.01641fF
C912 source.n301 bulk 0.00249fF
C913 source.n302 bulk 0.00260fF
C914 source.n303 bulk 0.00457fF
C915 source.n304 bulk 0.00483fF
C916 source.n305 bulk 0.02210fF
C917 source.n306 bulk 0.00595fF
C918 source.n307 bulk 0.00083fF
C919 source.n308 bulk 0.00094fF
C920 source.n309 bulk 0.00072fF
C921 source.n310 bulk 0.00061fF
C922 source.n311 bulk 0.00193fF
C923 source.t0 bulk 0.01072fF 
C924 source.t23 bulk 0.01072fF 
C925 source.n312 bulk 0.02204fF
C926 source.n313 bulk 0.00566fF
C927 source.n314 bulk 0.00088fF
C928 source.n315 bulk 0.01027fF
C929 source.n316 bulk 0.00166fF
C930 source.n317 bulk 0.00135fF
C931 source.n318 bulk 0.00114fF
C932 source.n319 bulk 0.00322fF
C933 source.n320 bulk 0.00260fF
C934 source.n321 bulk 0.00249fF
C935 source.n322 bulk 0.00083fF
C936 source.n323 bulk 0.00248fF
C937 source.n324 bulk 0.00155fF
C938 source.n325 bulk 0.00291fF
C939 source.n326 bulk 0.00156fF
C940 source.n327 bulk 0.00156fF
C941 source.n328 bulk 0.00177fF
C942 source.n329 bulk 0.01154fF
C943 source.n330 bulk 0.01641fF
C944 source.n331 bulk 0.00249fF
C945 source.n332 bulk 0.00260fF
C946 source.n333 bulk 0.00457fF
C947 source.n334 bulk 0.00483fF
C948 source.n335 bulk 0.02210fF
C949 source.n336 bulk 0.00595fF
C950 source.n337 bulk 0.00083fF
C951 source.n338 bulk 0.00094fF
C952 source.n339 bulk 0.00072fF
C953 source.n340 bulk 0.00061fF
C954 source.n341 bulk 0.00193fF
C955 source.t20 bulk 0.01072fF 
C956 source.t12 bulk 0.01072fF 
C957 source.n342 bulk 0.02204fF
C958 source.n343 bulk 0.00566fF
C959 source.n344 bulk 0.00088fF
C960 source.n345 bulk 0.01027fF
C961 source.n346 bulk 0.00166fF
C962 source.n347 bulk 0.00135fF
C963 source.n348 bulk 0.00114fF
C964 source.n349 bulk 0.00322fF
C965 source.n350 bulk 0.00260fF
C966 source.n351 bulk 0.00249fF
C967 source.n352 bulk 0.00083fF
C968 source.n353 bulk 0.00248fF
C969 source.n354 bulk 0.00155fF
C970 source.n355 bulk 0.00291fF
C971 source.n356 bulk 0.00156fF
C972 source.n357 bulk 0.00156fF
C973 source.n358 bulk 0.00177fF
C974 source.n359 bulk 0.01154fF
C975 source.n360 bulk 0.01641fF
C976 source.n361 bulk 0.00249fF
C977 source.n362 bulk 0.00260fF
C978 source.n363 bulk 0.00457fF
C979 source.n364 bulk 0.00483fF
C980 source.n365 bulk 0.02210fF
C981 source.n366 bulk 0.00595fF
C982 source.n367 bulk 0.00083fF
C983 source.n368 bulk 0.00094fF
C984 source.n369 bulk 0.00072fF
C985 source.n370 bulk 0.00061fF
C986 source.n371 bulk 0.00193fF
C987 source.t9 bulk 0.01072fF 
C988 source.t27 bulk 0.01072fF 
C989 source.n372 bulk 0.02204fF
C990 source.n373 bulk 0.00566fF
C991 source.n374 bulk 0.00088fF
C992 source.n375 bulk 0.01027fF
C993 source.n376 bulk 0.00166fF
C994 source.n377 bulk 0.00135fF
C995 source.n378 bulk 0.00114fF
C996 source.n379 bulk 0.00322fF
C997 source.n380 bulk 0.00260fF
C998 source.n381 bulk 0.00249fF
C999 source.n382 bulk 0.00083fF
C1000 source.n383 bulk 0.00248fF
C1001 source.n384 bulk 0.00155fF
C1002 source.n385 bulk 0.00291fF
C1003 source.n386 bulk 0.00156fF
C1004 source.n387 bulk 0.00156fF
C1005 source.n388 bulk 0.00177fF
C1006 source.n389 bulk 0.01154fF
C1007 source.n390 bulk 0.01641fF
C1008 source.n391 bulk 0.00249fF
C1009 source.n392 bulk 0.00260fF
C1010 source.n393 bulk 0.00457fF
C1011 source.n394 bulk 0.00483fF
C1012 source.n395 bulk 0.02210fF
C1013 source.n396 bulk 0.00595fF
C1014 source.n397 bulk 0.00083fF
C1015 source.n398 bulk 0.00094fF
C1016 source.n399 bulk 0.00072fF
C1017 source.n400 bulk 0.00061fF
C1018 source.n401 bulk 0.00193fF
C1019 source.t4 bulk 0.01072fF 
C1020 source.t17 bulk 0.01072fF 
C1021 source.n402 bulk 0.02204fF
C1022 source.n403 bulk 0.00566fF
C1023 source.n404 bulk 0.00088fF
C1024 source.n405 bulk 0.01027fF
C1025 source.n406 bulk 0.00166fF
C1026 source.n407 bulk 0.00135fF
C1027 source.n408 bulk 0.00114fF
C1028 source.n409 bulk 0.00322fF
C1029 source.n410 bulk 0.00260fF
C1030 source.n411 bulk 0.00249fF
C1031 source.n412 bulk 0.00083fF
C1032 source.n413 bulk 0.00248fF
C1033 source.n414 bulk 0.00155fF
C1034 source.n415 bulk 0.00291fF
C1035 source.n416 bulk 0.00156fF
C1036 source.n417 bulk 0.00156fF
C1037 source.n418 bulk 0.00177fF
C1038 source.n419 bulk 0.01154fF
C1039 source.n420 bulk 0.01641fF
C1040 source.n421 bulk 0.00249fF
C1041 source.n422 bulk 0.00260fF
C1042 source.n423 bulk 0.00457fF
C1043 source.n424 bulk 0.00483fF
C1044 source.n425 bulk 0.05308fF
C1045 source.n426 bulk 0.89954fF
C1046 source.n427 bulk 0.51852fF
C1047 source.n428 bulk 0.51852fF
C1048 source.n429 bulk 0.51852fF
C1049 source.n430 bulk 0.51852fF
C1050 source.n431 bulk 0.38991fF
C1051 source.n432 bulk 17.24210fF
C1052 a_85_n463.n0 bulk 0.37931fF
C1053 a_85_n463.n1 bulk 0.37942fF
C1054 a_85_n463.n2 bulk 0.37942fF
C1055 a_85_n463.n3 bulk 0.37942fF
C1056 a_85_n463.n4 bulk 0.37942fF
C1057 a_85_n463.n5 bulk 0.37942fF
C1058 a_85_n463.n6 bulk 0.37942fF
C1059 a_85_n463.n7 bulk 0.37942fF
C1060 a_85_n463.n8 bulk 0.37942fF
C1061 a_85_n463.n9 bulk 0.37942fF
C1062 a_85_n463.n10 bulk 0.37942fF
C1063 a_85_n463.n11 bulk 0.37942fF
C1064 a_85_n463.n12 bulk 0.37942fF
C1065 a_85_n463.n13 bulk 0.03885fF
C1066 a_85_n463.n14 bulk 0.00541fF
C1067 a_85_n463.n15 bulk 0.00613fF
C1068 a_85_n463.n16 bulk 0.82648fF
C1069 a_85_n463.n17 bulk 0.00469fF
C1070 a_85_n463.n18 bulk 0.00397fF
C1071 a_85_n463.n19 bulk 0.01262fF
C1072 a_85_n463.t1 bulk 0.07001fF 
C1073 a_85_n463.t10 bulk 0.07001fF 
C1074 a_85_n463.n20 bulk 0.14401fF
C1075 a_85_n463.n21 bulk 0.03696fF
C1076 a_85_n463.n22 bulk 0.00658fF
C1077 a_85_n463.n23 bulk 0.00541fF
C1078 a_85_n463.n24 bulk 0.01623fF
C1079 a_85_n463.n25 bulk 0.01010fF
C1080 a_85_n463.n26 bulk 0.03885fF
C1081 a_85_n463.n27 bulk 0.00541fF
C1082 a_85_n463.n28 bulk 0.00613fF
C1083 a_85_n463.n29 bulk 0.55932fF
C1084 a_85_n463.n30 bulk 0.00469fF
C1085 a_85_n463.n31 bulk 0.00397fF
C1086 a_85_n463.n32 bulk 0.01262fF
C1087 a_85_n463.t49 bulk 0.07001fF 
C1088 a_85_n463.t2 bulk 0.07001fF 
C1089 a_85_n463.n33 bulk 0.14401fF
C1090 a_85_n463.n34 bulk 0.03696fF
C1091 a_85_n463.n35 bulk 0.00658fF
C1092 a_85_n463.n36 bulk 0.00541fF
C1093 a_85_n463.n37 bulk 0.01623fF
C1094 a_85_n463.n38 bulk 0.01010fF
C1095 a_85_n463.n39 bulk 0.03885fF
C1096 a_85_n463.n40 bulk 0.00541fF
C1097 a_85_n463.n41 bulk 0.00613fF
C1098 a_85_n463.n42 bulk 0.55932fF
C1099 a_85_n463.n43 bulk 0.00469fF
C1100 a_85_n463.n44 bulk 0.00397fF
C1101 a_85_n463.n45 bulk 0.01262fF
C1102 a_85_n463.t4 bulk 0.07001fF 
C1103 a_85_n463.t39 bulk 0.07001fF 
C1104 a_85_n463.n46 bulk 0.14401fF
C1105 a_85_n463.n47 bulk 0.03696fF
C1106 a_85_n463.n48 bulk 0.00658fF
C1107 a_85_n463.n49 bulk 0.00541fF
C1108 a_85_n463.n50 bulk 0.01623fF
C1109 a_85_n463.n51 bulk 0.01010fF
C1110 a_85_n463.n52 bulk 0.03885fF
C1111 a_85_n463.n53 bulk 0.00541fF
C1112 a_85_n463.n54 bulk 0.00613fF
C1113 a_85_n463.n55 bulk 0.55932fF
C1114 a_85_n463.n56 bulk 0.00469fF
C1115 a_85_n463.n57 bulk 0.00397fF
C1116 a_85_n463.n58 bulk 0.01262fF
C1117 a_85_n463.t5 bulk 0.07001fF 
C1118 a_85_n463.t46 bulk 0.07001fF 
C1119 a_85_n463.n59 bulk 0.14401fF
C1120 a_85_n463.n60 bulk 0.03696fF
C1121 a_85_n463.n61 bulk 0.00658fF
C1122 a_85_n463.n62 bulk 0.00541fF
C1123 a_85_n463.n63 bulk 0.01623fF
C1124 a_85_n463.n64 bulk 0.01010fF
C1125 a_85_n463.n65 bulk 0.03885fF
C1126 a_85_n463.n66 bulk 0.00541fF
C1127 a_85_n463.n67 bulk 0.00613fF
C1128 a_85_n463.n68 bulk 0.55932fF
C1129 a_85_n463.n69 bulk 0.00469fF
C1130 a_85_n463.n70 bulk 0.00397fF
C1131 a_85_n463.n71 bulk 0.01262fF
C1132 a_85_n463.t50 bulk 0.07001fF 
C1133 a_85_n463.t9 bulk 0.07001fF 
C1134 a_85_n463.n72 bulk 0.14401fF
C1135 a_85_n463.n73 bulk 0.03696fF
C1136 a_85_n463.n74 bulk 0.00658fF
C1137 a_85_n463.n75 bulk 0.00541fF
C1138 a_85_n463.n76 bulk 0.01623fF
C1139 a_85_n463.n77 bulk 0.01010fF
C1140 a_85_n463.n78 bulk 0.03885fF
C1141 a_85_n463.n79 bulk 0.00541fF
C1142 a_85_n463.n80 bulk 0.00613fF
C1143 a_85_n463.n81 bulk 0.55932fF
C1144 a_85_n463.n82 bulk 0.00469fF
C1145 a_85_n463.n83 bulk 0.00397fF
C1146 a_85_n463.n84 bulk 0.01262fF
C1147 a_85_n463.t41 bulk 0.07001fF 
C1148 a_85_n463.t6 bulk 0.07001fF 
C1149 a_85_n463.n85 bulk 0.14401fF
C1150 a_85_n463.n86 bulk 0.03696fF
C1151 a_85_n463.n87 bulk 0.00658fF
C1152 a_85_n463.n88 bulk 0.00541fF
C1153 a_85_n463.n89 bulk 0.01623fF
C1154 a_85_n463.n90 bulk 0.01010fF
C1155 a_85_n463.n91 bulk 0.03885fF
C1156 a_85_n463.n92 bulk 0.00541fF
C1157 a_85_n463.n93 bulk 0.00613fF
C1158 a_85_n463.n94 bulk 0.55932fF
C1159 a_85_n463.n95 bulk 0.00469fF
C1160 a_85_n463.n96 bulk 0.00397fF
C1161 a_85_n463.n97 bulk 0.01262fF
C1162 a_85_n463.t44 bulk 0.07001fF 
C1163 a_85_n463.t40 bulk 0.07001fF 
C1164 a_85_n463.n98 bulk 0.14401fF
C1165 a_85_n463.n99 bulk 0.03696fF
C1166 a_85_n463.n100 bulk 0.00658fF
C1167 a_85_n463.n101 bulk 0.00541fF
C1168 a_85_n463.n102 bulk 0.01623fF
C1169 a_85_n463.n103 bulk 0.01010fF
C1170 a_85_n463.n104 bulk 0.03885fF
C1171 a_85_n463.n105 bulk 0.00541fF
C1172 a_85_n463.n106 bulk 0.00613fF
C1173 a_85_n463.n107 bulk 0.55932fF
C1174 a_85_n463.n108 bulk 0.00469fF
C1175 a_85_n463.n109 bulk 0.00397fF
C1176 a_85_n463.n110 bulk 0.01262fF
C1177 a_85_n463.t45 bulk 0.07001fF 
C1178 a_85_n463.t43 bulk 0.07001fF 
C1179 a_85_n463.n111 bulk 0.14401fF
C1180 a_85_n463.n112 bulk 0.03696fF
C1181 a_85_n463.n113 bulk 0.00658fF
C1182 a_85_n463.n114 bulk 0.00541fF
C1183 a_85_n463.n115 bulk 0.01623fF
C1184 a_85_n463.n116 bulk 0.01010fF
C1185 a_85_n463.n117 bulk 0.03885fF
C1186 a_85_n463.n118 bulk 0.00541fF
C1187 a_85_n463.n119 bulk 0.00613fF
C1188 a_85_n463.n120 bulk 0.55932fF
C1189 a_85_n463.n121 bulk 0.00469fF
C1190 a_85_n463.n122 bulk 0.00397fF
C1191 a_85_n463.n123 bulk 0.01262fF
C1192 a_85_n463.t42 bulk 0.07001fF 
C1193 a_85_n463.t53 bulk 0.07001fF 
C1194 a_85_n463.n124 bulk 0.14401fF
C1195 a_85_n463.n125 bulk 0.03696fF
C1196 a_85_n463.n126 bulk 0.00658fF
C1197 a_85_n463.n127 bulk 0.00541fF
C1198 a_85_n463.n128 bulk 0.01623fF
C1199 a_85_n463.n129 bulk 0.01010fF
C1200 a_85_n463.n130 bulk 0.03885fF
C1201 a_85_n463.n131 bulk 0.00541fF
C1202 a_85_n463.n132 bulk 0.00613fF
C1203 a_85_n463.n133 bulk 0.55932fF
C1204 a_85_n463.n134 bulk 0.00469fF
C1205 a_85_n463.n135 bulk 0.00397fF
C1206 a_85_n463.n136 bulk 0.01262fF
C1207 a_85_n463.t51 bulk 0.07001fF 
C1208 a_85_n463.t55 bulk 0.07001fF 
C1209 a_85_n463.n137 bulk 0.14401fF
C1210 a_85_n463.n138 bulk 0.03696fF
C1211 a_85_n463.n139 bulk 0.00658fF
C1212 a_85_n463.n140 bulk 0.00541fF
C1213 a_85_n463.n141 bulk 0.01623fF
C1214 a_85_n463.n142 bulk 0.01010fF
C1215 a_85_n463.n143 bulk 0.03885fF
C1216 a_85_n463.n144 bulk 0.00541fF
C1217 a_85_n463.n145 bulk 0.00613fF
C1218 a_85_n463.n146 bulk 0.55932fF
C1219 a_85_n463.n147 bulk 0.00469fF
C1220 a_85_n463.n148 bulk 0.00397fF
C1221 a_85_n463.n149 bulk 0.01262fF
C1222 a_85_n463.t48 bulk 0.07001fF 
C1223 a_85_n463.t47 bulk 0.07001fF 
C1224 a_85_n463.n150 bulk 0.14401fF
C1225 a_85_n463.n151 bulk 0.03696fF
C1226 a_85_n463.n152 bulk 0.00658fF
C1227 a_85_n463.n153 bulk 0.00541fF
C1228 a_85_n463.n154 bulk 0.01623fF
C1229 a_85_n463.n155 bulk 0.01010fF
C1230 a_85_n463.n156 bulk 0.03885fF
C1231 a_85_n463.n157 bulk 0.00541fF
C1232 a_85_n463.n158 bulk 0.00613fF
C1233 a_85_n463.n159 bulk 0.55932fF
C1234 a_85_n463.n160 bulk 0.00469fF
C1235 a_85_n463.n161 bulk 0.00397fF
C1236 a_85_n463.n162 bulk 0.01262fF
C1237 a_85_n463.t3 bulk 0.07001fF 
C1238 a_85_n463.t52 bulk 0.07001fF 
C1239 a_85_n463.n163 bulk 0.14401fF
C1240 a_85_n463.n164 bulk 0.03696fF
C1241 a_85_n463.n165 bulk 0.00658fF
C1242 a_85_n463.n166 bulk 0.00541fF
C1243 a_85_n463.n167 bulk 0.01623fF
C1244 a_85_n463.n168 bulk 0.01010fF
C1245 a_85_n463.n169 bulk 0.03886fF
C1246 a_85_n463.n170 bulk 0.00541fF
C1247 a_85_n463.n171 bulk 0.00613fF
C1248 a_85_n463.n172 bulk 0.82658fF
C1249 a_85_n463.n173 bulk 0.00469fF
C1250 a_85_n463.n174 bulk 0.00397fF
C1251 a_85_n463.n175 bulk 0.01262fF
C1252 a_85_n463.t8 bulk 0.07001fF 
C1253 a_85_n463.t54 bulk 0.07001fF 
C1254 a_85_n463.n176 bulk 0.14401fF
C1255 a_85_n463.n177 bulk 0.03696fF
C1256 a_85_n463.n178 bulk 0.00658fF
C1257 a_85_n463.n179 bulk 0.00541fF
C1258 a_85_n463.n180 bulk 0.01623fF
C1259 a_85_n463.n181 bulk 0.01010fF
C1260 a_85_n463.n182 bulk 0.04621fF
C1261 a_85_n463.n183 bulk 0.09032fF
C1262 a_85_n463.n184 bulk 0.04621fF
C1263 a_85_n463.n185 bulk 0.09032fF
C1264 a_85_n463.n186 bulk 0.04621fF
C1265 a_85_n463.n187 bulk 0.09032fF
C1266 a_85_n463.n188 bulk 0.04621fF
C1267 a_85_n463.n189 bulk 0.09032fF
C1268 a_85_n463.n190 bulk 0.04621fF
C1269 a_85_n463.n191 bulk 0.09032fF
C1270 a_85_n463.n192 bulk 0.04621fF
C1271 a_85_n463.n193 bulk 0.09032fF
C1272 a_85_n463.n194 bulk 0.04621fF
C1273 a_85_n463.n195 bulk 0.09032fF
C1274 a_85_n463.n196 bulk 0.04621fF
C1275 a_85_n463.n197 bulk 0.09032fF
C1276 a_85_n463.n198 bulk 0.04621fF
C1277 a_85_n463.n199 bulk 0.09032fF
C1278 a_85_n463.n200 bulk 0.04621fF
C1279 a_85_n463.n201 bulk 0.09032fF
C1280 a_85_n463.n202 bulk 0.04621fF
C1281 a_85_n463.n203 bulk 0.09032fF
C1282 a_85_n463.n204 bulk 0.04621fF
C1283 a_85_n463.n205 bulk 0.09032fF
C1284 a_85_n463.n206 bulk 0.04621fF
C1285 a_85_n463.n207 bulk 0.09032fF
C1286 a_85_n463.n208 bulk 0.04621fF
C1287 a_85_n463.n209 bulk 0.09032fF
C1288 a_85_n463.n210 bulk 0.04621fF
C1289 a_85_n463.n211 bulk 0.09032fF
C1290 a_85_n463.t7 bulk 0.07001fF 
C1291 a_85_n463.n212 bulk 0.00541fF
C1292 a_85_n463.n213 bulk 0.00541fF
C1293 a_85_n463.n214 bulk 0.00613fF
C1294 a_85_n463.n215 bulk 0.03885fF
C1295 a_85_n463.n216 bulk 0.01262fF
C1296 a_85_n463.n217 bulk 0.00397fF
C1297 a_85_n463.n218 bulk 0.00469fF
C1298 a_85_n463.n219 bulk 0.03877fF
C1299 a_85_n463.n220 bulk 0.00541fF
C1300 a_85_n463.n221 bulk 0.00701fF
C1301 a_85_n463.n222 bulk 0.13774fF
C1302 a_85_n463.n223 bulk 0.00541fF
C1303 a_85_n463.n224 bulk 0.01623fF
C1304 a_85_n463.n225 bulk 0.01010fF
C1305 a_85_n463.n226 bulk 0.00469fF
C1306 a_85_n463.n227 bulk 0.00397fF
C1307 a_85_n463.n228 bulk 0.01262fF
C1308 a_85_n463.t27 bulk 0.07001fF 
C1309 a_85_n463.t37 bulk 0.07001fF 
C1310 a_85_n463.n229 bulk 0.14401fF
C1311 a_85_n463.n230 bulk 0.03700fF
C1312 a_85_n463.n231 bulk 0.00577fF
C1313 a_85_n463.n232 bulk 0.11190fF
C1314 a_85_n463.n233 bulk 0.19775fF
C1315 a_85_n463.n234 bulk 0.03877fF
C1316 a_85_n463.n235 bulk 0.00541fF
C1317 a_85_n463.n236 bulk 0.00701fF
C1318 a_85_n463.n237 bulk 0.13774fF
C1319 a_85_n463.n238 bulk 0.00541fF
C1320 a_85_n463.n239 bulk 0.01623fF
C1321 a_85_n463.n240 bulk 0.01010fF
C1322 a_85_n463.n241 bulk 0.00469fF
C1323 a_85_n463.n242 bulk 0.00397fF
C1324 a_85_n463.n243 bulk 0.01262fF
C1325 a_85_n463.t30 bulk 0.07001fF 
C1326 a_85_n463.t32 bulk 0.07001fF 
C1327 a_85_n463.n244 bulk 0.14401fF
C1328 a_85_n463.n245 bulk 0.03700fF
C1329 a_85_n463.n246 bulk 0.00577fF
C1330 a_85_n463.n247 bulk 0.11190fF
C1331 a_85_n463.n248 bulk 0.19775fF
C1332 a_85_n463.n249 bulk 0.03877fF
C1333 a_85_n463.n250 bulk 0.00541fF
C1334 a_85_n463.n251 bulk 0.00701fF
C1335 a_85_n463.n252 bulk 0.13774fF
C1336 a_85_n463.n253 bulk 0.00541fF
C1337 a_85_n463.n254 bulk 0.01623fF
C1338 a_85_n463.n255 bulk 0.01010fF
C1339 a_85_n463.n256 bulk 0.00469fF
C1340 a_85_n463.n257 bulk 0.00397fF
C1341 a_85_n463.n258 bulk 0.01262fF
C1342 a_85_n463.t19 bulk 0.07001fF 
C1343 a_85_n463.n259 bulk 0.19704fF
C1344 a_85_n463.n260 bulk 0.03700fF
C1345 a_85_n463.n261 bulk 0.00577fF
C1346 a_85_n463.n262 bulk 0.11190fF
C1347 a_85_n463.n263 bulk 0.26569fF
C1348 a_85_n463.n264 bulk 0.36565fF
C1349 a_85_n463.n265 bulk 0.36565fF
C1350 a_85_n463.n266 bulk 0.03877fF
C1351 a_85_n463.n267 bulk 0.00541fF
C1352 a_85_n463.n268 bulk 0.00701fF
C1353 a_85_n463.n269 bulk 0.13774fF
C1354 a_85_n463.n270 bulk 0.00541fF
C1355 a_85_n463.n271 bulk 0.01623fF
C1356 a_85_n463.n272 bulk 0.01010fF
C1357 a_85_n463.n273 bulk 0.00469fF
C1358 a_85_n463.n274 bulk 0.00397fF
C1359 a_85_n463.n275 bulk 0.01262fF
C1360 a_85_n463.t17 bulk 0.07001fF 
C1361 a_85_n463.t24 bulk 0.07001fF 
C1362 a_85_n463.n276 bulk 0.14401fF
C1363 a_85_n463.n277 bulk 0.03700fF
C1364 a_85_n463.n278 bulk 0.00577fF
C1365 a_85_n463.n279 bulk 0.11190fF
C1366 a_85_n463.n280 bulk 0.19775fF
C1367 a_85_n463.n281 bulk 0.03877fF
C1368 a_85_n463.n282 bulk 0.00541fF
C1369 a_85_n463.n283 bulk 0.00701fF
C1370 a_85_n463.n284 bulk 0.13774fF
C1371 a_85_n463.n285 bulk 0.00541fF
C1372 a_85_n463.n286 bulk 0.01623fF
C1373 a_85_n463.n287 bulk 0.01010fF
C1374 a_85_n463.n288 bulk 0.00469fF
C1375 a_85_n463.n289 bulk 0.00397fF
C1376 a_85_n463.n290 bulk 0.01262fF
C1377 a_85_n463.t12 bulk 0.07001fF 
C1378 a_85_n463.t21 bulk 0.07001fF 
C1379 a_85_n463.n291 bulk 0.14401fF
C1380 a_85_n463.n292 bulk 0.03700fF
C1381 a_85_n463.n293 bulk 0.00577fF
C1382 a_85_n463.n294 bulk 0.11190fF
C1383 a_85_n463.n295 bulk 0.19775fF
C1384 a_85_n463.n296 bulk 0.03877fF
C1385 a_85_n463.n297 bulk 0.00541fF
C1386 a_85_n463.n298 bulk 0.00701fF
C1387 a_85_n463.n299 bulk 0.13774fF
C1388 a_85_n463.n300 bulk 0.00541fF
C1389 a_85_n463.n301 bulk 0.01623fF
C1390 a_85_n463.n302 bulk 0.01010fF
C1391 a_85_n463.n303 bulk 0.00469fF
C1392 a_85_n463.n304 bulk 0.00397fF
C1393 a_85_n463.n305 bulk 0.01262fF
C1394 a_85_n463.t22 bulk 0.07001fF 
C1395 a_85_n463.t11 bulk 0.07001fF 
C1396 a_85_n463.n306 bulk 0.14401fF
C1397 a_85_n463.n307 bulk 0.03700fF
C1398 a_85_n463.n308 bulk 0.00577fF
C1399 a_85_n463.n309 bulk 0.11190fF
C1400 a_85_n463.n310 bulk 0.19775fF
C1401 a_85_n463.n311 bulk 0.03877fF
C1402 a_85_n463.n312 bulk 0.00541fF
C1403 a_85_n463.n313 bulk 0.00701fF
C1404 a_85_n463.n314 bulk 0.13774fF
C1405 a_85_n463.n315 bulk 0.00541fF
C1406 a_85_n463.n316 bulk 0.01623fF
C1407 a_85_n463.n317 bulk 0.01010fF
C1408 a_85_n463.n318 bulk 0.00469fF
C1409 a_85_n463.n319 bulk 0.00397fF
C1410 a_85_n463.n320 bulk 0.01262fF
C1411 a_85_n463.t36 bulk 0.07001fF 
C1412 a_85_n463.t31 bulk 0.07001fF 
C1413 a_85_n463.n321 bulk 0.14401fF
C1414 a_85_n463.n322 bulk 0.03700fF
C1415 a_85_n463.n323 bulk 0.00577fF
C1416 a_85_n463.n324 bulk 0.11190fF
C1417 a_85_n463.n325 bulk 0.19775fF
C1418 a_85_n463.n326 bulk 0.03877fF
C1419 a_85_n463.n327 bulk 0.00541fF
C1420 a_85_n463.n328 bulk 0.00701fF
C1421 a_85_n463.n329 bulk 0.13774fF
C1422 a_85_n463.n330 bulk 0.00541fF
C1423 a_85_n463.n331 bulk 0.01623fF
C1424 a_85_n463.n332 bulk 0.01010fF
C1425 a_85_n463.n333 bulk 0.00469fF
C1426 a_85_n463.n334 bulk 0.00397fF
C1427 a_85_n463.n335 bulk 0.01262fF
C1428 a_85_n463.t16 bulk 0.07001fF 
C1429 a_85_n463.t18 bulk 0.07001fF 
C1430 a_85_n463.n336 bulk 0.14401fF
C1431 a_85_n463.n337 bulk 0.03700fF
C1432 a_85_n463.n338 bulk 0.00577fF
C1433 a_85_n463.n339 bulk 0.11190fF
C1434 a_85_n463.n340 bulk 0.19775fF
C1435 a_85_n463.n341 bulk 0.03877fF
C1436 a_85_n463.n342 bulk 0.00541fF
C1437 a_85_n463.n343 bulk 0.00701fF
C1438 a_85_n463.n344 bulk 0.13774fF
C1439 a_85_n463.n345 bulk 0.00541fF
C1440 a_85_n463.n346 bulk 0.01623fF
C1441 a_85_n463.n347 bulk 0.01010fF
C1442 a_85_n463.n348 bulk 0.00469fF
C1443 a_85_n463.n349 bulk 0.00397fF
C1444 a_85_n463.n350 bulk 0.01262fF
C1445 a_85_n463.t14 bulk 0.07001fF 
C1446 a_85_n463.t29 bulk 0.07001fF 
C1447 a_85_n463.n351 bulk 0.14401fF
C1448 a_85_n463.n352 bulk 0.03700fF
C1449 a_85_n463.n353 bulk 0.00577fF
C1450 a_85_n463.n354 bulk 0.11190fF
C1451 a_85_n463.n355 bulk 0.19775fF
C1452 a_85_n463.n356 bulk 0.03877fF
C1453 a_85_n463.n357 bulk 0.00541fF
C1454 a_85_n463.n358 bulk 0.00701fF
C1455 a_85_n463.n359 bulk 0.13774fF
C1456 a_85_n463.n360 bulk 0.00541fF
C1457 a_85_n463.n361 bulk 0.01623fF
C1458 a_85_n463.n362 bulk 0.01010fF
C1459 a_85_n463.n363 bulk 0.00469fF
C1460 a_85_n463.n364 bulk 0.00397fF
C1461 a_85_n463.n365 bulk 0.01262fF
C1462 a_85_n463.t13 bulk 0.07001fF 
C1463 a_85_n463.t23 bulk 0.07001fF 
C1464 a_85_n463.n366 bulk 0.14401fF
C1465 a_85_n463.n367 bulk 0.03700fF
C1466 a_85_n463.n368 bulk 0.00577fF
C1467 a_85_n463.n369 bulk 0.11190fF
C1468 a_85_n463.n370 bulk 0.19775fF
C1469 a_85_n463.n371 bulk 0.03877fF
C1470 a_85_n463.n372 bulk 0.00541fF
C1471 a_85_n463.n373 bulk 0.00701fF
C1472 a_85_n463.n374 bulk 0.13774fF
C1473 a_85_n463.n375 bulk 0.00541fF
C1474 a_85_n463.n376 bulk 0.01623fF
C1475 a_85_n463.n377 bulk 0.01010fF
C1476 a_85_n463.n378 bulk 0.00469fF
C1477 a_85_n463.n379 bulk 0.00397fF
C1478 a_85_n463.n380 bulk 0.01262fF
C1479 a_85_n463.t25 bulk 0.07001fF 
C1480 a_85_n463.t26 bulk 0.07001fF 
C1481 a_85_n463.n381 bulk 0.14401fF
C1482 a_85_n463.n382 bulk 0.03700fF
C1483 a_85_n463.n383 bulk 0.00577fF
C1484 a_85_n463.n384 bulk 0.11190fF
C1485 a_85_n463.n385 bulk 0.19775fF
C1486 a_85_n463.n386 bulk 0.03877fF
C1487 a_85_n463.n387 bulk 0.00541fF
C1488 a_85_n463.n388 bulk 0.00701fF
C1489 a_85_n463.n389 bulk 0.13774fF
C1490 a_85_n463.n390 bulk 0.00541fF
C1491 a_85_n463.n391 bulk 0.01623fF
C1492 a_85_n463.n392 bulk 0.01010fF
C1493 a_85_n463.n393 bulk 0.00469fF
C1494 a_85_n463.n394 bulk 0.00397fF
C1495 a_85_n463.n395 bulk 0.01262fF
C1496 a_85_n463.t34 bulk 0.07001fF 
C1497 a_85_n463.t38 bulk 0.07001fF 
C1498 a_85_n463.n396 bulk 0.14401fF
C1499 a_85_n463.n397 bulk 0.03700fF
C1500 a_85_n463.n398 bulk 0.00577fF
C1501 a_85_n463.n399 bulk 0.11190fF
C1502 a_85_n463.n400 bulk 0.19775fF
C1503 a_85_n463.n401 bulk 0.03877fF
C1504 a_85_n463.n402 bulk 0.00541fF
C1505 a_85_n463.n403 bulk 0.00701fF
C1506 a_85_n463.n404 bulk 0.13774fF
C1507 a_85_n463.n405 bulk 0.00541fF
C1508 a_85_n463.n406 bulk 0.01623fF
C1509 a_85_n463.n407 bulk 0.01010fF
C1510 a_85_n463.n408 bulk 0.00469fF
C1511 a_85_n463.n409 bulk 0.00397fF
C1512 a_85_n463.n410 bulk 0.01262fF
C1513 a_85_n463.t35 bulk 0.07001fF 
C1514 a_85_n463.t15 bulk 0.07001fF 
C1515 a_85_n463.n411 bulk 0.14401fF
C1516 a_85_n463.n412 bulk 0.03700fF
C1517 a_85_n463.n413 bulk 0.00577fF
C1518 a_85_n463.n414 bulk 0.11190fF
C1519 a_85_n463.n415 bulk 0.19775fF
C1520 a_85_n463.n416 bulk 0.03877fF
C1521 a_85_n463.n417 bulk 0.00541fF
C1522 a_85_n463.n418 bulk 0.00701fF
C1523 a_85_n463.n419 bulk 0.13774fF
C1524 a_85_n463.n420 bulk 0.00541fF
C1525 a_85_n463.n421 bulk 0.01623fF
C1526 a_85_n463.n422 bulk 0.01010fF
C1527 a_85_n463.n423 bulk 0.00469fF
C1528 a_85_n463.n424 bulk 0.00397fF
C1529 a_85_n463.n425 bulk 0.01262fF
C1530 a_85_n463.t33 bulk 0.07001fF 
C1531 a_85_n463.t20 bulk 0.07001fF 
C1532 a_85_n463.n426 bulk 0.14401fF
C1533 a_85_n463.n427 bulk 0.03700fF
C1534 a_85_n463.n428 bulk 0.00577fF
C1535 a_85_n463.n429 bulk 0.11190fF
C1536 a_85_n463.n430 bulk 0.19775fF
C1537 a_85_n463.n431 bulk 0.03877fF
C1538 a_85_n463.n432 bulk 0.00541fF
C1539 a_85_n463.n433 bulk 0.00701fF
C1540 a_85_n463.n434 bulk 0.13774fF
C1541 a_85_n463.n435 bulk 0.00541fF
C1542 a_85_n463.n436 bulk 0.01623fF
C1543 a_85_n463.n437 bulk 0.01010fF
C1544 a_85_n463.n438 bulk 0.00469fF
C1545 a_85_n463.n439 bulk 0.00397fF
C1546 a_85_n463.n440 bulk 0.01262fF
C1547 a_85_n463.t28 bulk 0.07001fF 
C1548 a_85_n463.n441 bulk 0.19704fF
C1549 a_85_n463.n442 bulk 0.03700fF
C1550 a_85_n463.n443 bulk 0.00577fF
C1551 a_85_n463.n444 bulk 0.11190fF
C1552 a_85_n463.n445 bulk 0.26569fF
C1553 a_85_n463.n446 bulk 0.36565fF
C1554 a_85_n463.n447 bulk 0.36565fF
C1555 a_85_n463.n448 bulk 0.36565fF
C1556 a_85_n463.n449 bulk 0.36565fF
C1557 a_85_n463.n450 bulk 0.36565fF
C1558 a_85_n463.n451 bulk 0.36565fF
C1559 a_85_n463.n452 bulk 0.36565fF
C1560 a_85_n463.n453 bulk 0.36565fF
C1561 a_85_n463.n454 bulk 0.36565fF
C1562 a_85_n463.n455 bulk 0.36565fF
C1563 a_85_n463.n456 bulk 0.36565fF
C1564 a_85_n463.n457 bulk 0.31510fF
C1565 a_85_n463.n458 bulk 0.14776fF
C1566 a_85_n463.n459 bulk 0.18986fF
C1567 a_85_n463.n460 bulk 0.28355fF
C1568 a_85_n463.n461 bulk 0.01623fF
C1569 a_85_n463.n462 bulk 0.01010fF
C1570 a_85_n463.n463 bulk 0.00904fF
C1571 a_85_n463.n464 bulk 0.03697fF
C1572 a_85_n463.n465 bulk 0.14400fF
C1573 a_85_n463.t0 bulk 0.07001fF 
C1574 bias1_input.n0 bulk 0.01551fF
C1575 bias1_input.n1 bulk 0.00965fF
C1576 bias1_input.n2 bulk 0.01413fF
C1577 bias1_input.n3 bulk 0.00896fF
C1578 bias1_input.n4 bulk 0.00276fF
C1579 bias1_input.n5 bulk 0.01034fF
C1580 bias1_input.n6 bulk 0.00965fF
C1581 bias1_input.n7 bulk 0.01034fF
C1582 bias1_input.n8 bulk 0.00930fF
C1583 bias1_input.n9 bulk 0.01275fF
C1584 bias1_input.n10 bulk 0.01413fF
C1585 bias1_input.n11 bulk 0.01137fF
C1586 bias1_input.n12 bulk 0.00896fF
C1587 bias1_input.n13 bulk 0.00827fF
C1588 bias1_input.n14 bulk 0.01034fF
C1589 bias1_input.n15 bulk 0.00724fF
C1590 bias1_input.n16 bulk 0.00724fF
C1591 bias1_input.n17 bulk 0.00724fF
C1592 bias1_input.n18 bulk 0.00724fF
C1593 bias1_input.n19 bulk 0.01476fF
C1594 bias1_input.n20 bulk 0.00758fF
C1595 bias1_input.n21 bulk 0.00999fF
C1596 bias1_input.n22 bulk 0.00999fF
C1597 bias1_input.n23 bulk 0.00724fF
C1598 bias1_input.n24 bulk 0.01413fF
C1599 bias1_input.n25 bulk 0.00896fF
C1600 bias1_input.n26 bulk 0.01689fF
C1601 bias1_input.n27 bulk 0.02102fF
C1602 bias1_input.n28 bulk 0.00896fF
C1603 bias1_input.n29 bulk 0.01241fF
C1604 bias1_input.t23 bulk 0.02935fF 
C1605 bias1_input.n30 bulk 0.44560fF
C1606 bias1_input.t18 bulk 0.02935fF 
C1607 bias1_input.n31 bulk 0.21674fF
C1608 bias1_input.t7 bulk 0.02935fF 
C1609 bias1_input.n32 bulk 0.21674fF
C1610 bias1_input.t27 bulk 0.02935fF 
C1611 bias1_input.n33 bulk 0.21674fF
C1612 bias1_input.t9 bulk 0.02935fF 
C1613 bias1_input.n34 bulk 0.21674fF
C1614 bias1_input.t20 bulk 0.02935fF 
C1615 bias1_input.n35 bulk 0.21674fF
C1616 bias1_input.t13 bulk 0.02935fF 
C1617 bias1_input.n36 bulk 0.21674fF
C1618 bias1_input.t2 bulk 0.02935fF 
C1619 bias1_input.n37 bulk 0.21674fF
C1620 bias1_input.t19 bulk 0.02935fF 
C1621 bias1_input.n38 bulk 0.21674fF
C1622 bias1_input.t8 bulk 0.02935fF 
C1623 bias1_input.n39 bulk 0.21674fF
C1624 bias1_input.t21 bulk 0.02935fF 
C1625 bias1_input.n40 bulk 0.21674fF
C1626 bias1_input.t14 bulk 0.02935fF 
C1627 bias1_input.n41 bulk 0.21674fF
C1628 bias1_input.t3 bulk 0.02935fF 
C1629 bias1_input.n42 bulk 0.21674fF
C1630 bias1_input.t24 bulk 0.02935fF 
C1631 bias1_input.n43 bulk 0.24603fF
C1632 bias1_input.n44 bulk 0.14489fF
C1633 bias1_input.n45 bulk 0.00548fF
C1634 bias1_input.n46 bulk 0.01491fF
C1635 bias1_input.n47 bulk 0.00758fF
C1636 bias1_input.n48 bulk 0.00724fF
C1637 bias1_input.n49 bulk 0.00724fF
C1638 bias1_input.n50 bulk 0.00724fF
C1639 bias1_input.n51 bulk 0.03000fF
C1640 bias1_input.n52 bulk 0.03063fF
C1641 bias1_input.n53 bulk 0.14689fF
C1642 bias1_input.n54 bulk 0.04103fF
C1643 bias1_input.n55 bulk 0.04924fF
C1644 bias1_input.n56 bulk 0.04103fF
C1645 bias1_input.n57 bulk 0.04103fF
C1646 bias1_input.n58 bulk 0.04924fF
C1647 bias1_input.n59 bulk 0.03283fF
C1648 bias1_input.n60 bulk 0.01551fF
C1649 bias1_input.n61 bulk 0.01413fF
C1650 bias1_input.n62 bulk 0.00896fF
C1651 bias1_input.n63 bulk 0.00965fF
C1652 bias1_input.n64 bulk 0.00276fF
C1653 bias1_input.n65 bulk 0.01034fF
C1654 bias1_input.n66 bulk 0.00965fF
C1655 bias1_input.n67 bulk 0.01034fF
C1656 bias1_input.n68 bulk 0.00930fF
C1657 bias1_input.n69 bulk 0.01275fF
C1658 bias1_input.n70 bulk 0.01413fF
C1659 bias1_input.n71 bulk 0.01137fF
C1660 bias1_input.n72 bulk 0.00896fF
C1661 bias1_input.n73 bulk 0.00827fF
C1662 bias1_input.n74 bulk 0.01034fF
C1663 bias1_input.n75 bulk 0.00724fF
C1664 bias1_input.n76 bulk 0.00724fF
C1665 bias1_input.n77 bulk 0.00724fF
C1666 bias1_input.n78 bulk 0.00724fF
C1667 bias1_input.n79 bulk 0.01476fF
C1668 bias1_input.n80 bulk 0.00758fF
C1669 bias1_input.n81 bulk 0.00999fF
C1670 bias1_input.n82 bulk 0.00999fF
C1671 bias1_input.n83 bulk 0.01413fF
C1672 bias1_input.n84 bulk 0.00896fF
C1673 bias1_input.n85 bulk 0.01689fF
C1674 bias1_input.n86 bulk 0.02102fF
C1675 bias1_input.n87 bulk 0.00896fF
C1676 bias1_input.n88 bulk 0.01241fF
C1677 bias1_input.t10 bulk 0.03515fF 
C1678 bias1_input.n89 bulk 0.42868fF
C1679 bias1_input.t0 bulk 0.03515fF 
C1680 bias1_input.n90 bulk 0.21093fF
C1681 bias1_input.t15 bulk 0.03515fF 
C1682 bias1_input.n91 bulk 0.21093fF
C1683 bias1_input.t4 bulk 0.03515fF 
C1684 bias1_input.n92 bulk 0.21093fF
C1685 bias1_input.t16 bulk 0.03515fF 
C1686 bias1_input.n93 bulk 0.21093fF
C1687 bias1_input.t5 bulk 0.03515fF 
C1688 bias1_input.n94 bulk 0.21093fF
C1689 bias1_input.t25 bulk 0.03515fF 
C1690 bias1_input.n95 bulk 0.21093fF
C1691 bias1_input.t11 bulk 0.03515fF 
C1692 bias1_input.n96 bulk 0.21093fF
C1693 bias1_input.t22 bulk 0.03515fF 
C1694 bias1_input.n97 bulk 0.21093fF
C1695 bias1_input.t17 bulk 0.03515fF 
C1696 bias1_input.n98 bulk 0.21093fF
C1697 bias1_input.t6 bulk 0.03515fF 
C1698 bias1_input.n99 bulk 0.21093fF
C1699 bias1_input.t26 bulk 0.03515fF 
C1700 bias1_input.n100 bulk 0.21093fF
C1701 bias1_input.t12 bulk 0.03515fF 
C1702 bias1_input.n101 bulk 0.21093fF
C1703 bias1_input.t1 bulk 0.03515fF 
C1704 bias1_input.n102 bulk 0.20714fF
C1705 bias1_input.n103 bulk 0.11180fF
C1706 bias1_input.n104 bulk 0.00548fF
C1707 bias1_input.n105 bulk 0.00724fF
C1708 bias1_input.n106 bulk 0.01491fF
C1709 bias1_input.n107 bulk 0.00758fF
C1710 bias1_input.n108 bulk 0.00724fF
C1711 bias1_input.n109 bulk 0.00724fF
C1712 bias1_input.n110 bulk 0.00724fF
C1713 bias1_input.n111 bulk 0.03001fF
C1714 bias1_input.n112 bulk 0.03063fF
C1715 bias1_input.n113 bulk 0.14689fF
C1716 bias1_input.n114 bulk 0.04103fF
C1717 bias1_input.n115 bulk 0.04924fF
C1718 bias1_input.n116 bulk 0.04103fF
C1719 bias1_input.n117 bulk 0.04103fF
C1720 bias1_input.n118 bulk 0.04924fF
C1721 bias1_input.n119 bulk 0.03283fF
C1722 bias1_input.n120 bulk 4.64110fF
