* NGSPICE file created from VGA_final.ext - technology: sky130A

.subckt VGA_final RF_in RF_out Vctrl Vgg_1v2 Vdd_1v8 Gnd
XMOM_capacitor_0 Vdd_1v8 RF_out Gnd MOM_capacitor
X0 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X2 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D0 Gnd Vdd_1v8 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X8 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X11 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X21 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X23 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X24 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X28 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X30 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X32 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X33 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X34 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X35 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X36 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 a_47_7088# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X43 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X44 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X45 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X46 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X47 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X48 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X49 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X50 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X51 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X52 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X53 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X54 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X55 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X56 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X57 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X58 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X60 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X61 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X62 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X63 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X64 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X65 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X66 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X67 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X68 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X69 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X70 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X71 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X72 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X73 Vdd_1v8 Gnd sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X74 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X75 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 Vctrl a_n45858_n64215# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X76 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X78 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X79 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X80 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X82 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X83 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X84 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X85 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X86 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X87 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X88 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X92 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X93 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X94 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X95 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X96 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X98 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X99 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X100 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X101 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X102 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X103 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X104 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X105 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X106 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X107 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X108 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X109 Gnd Gnd a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X110 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X111 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X112 a_n45858_n24875# RF_in sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X113 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X114 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X115 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X116 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X117 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X118 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X120 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X122 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X123 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X124 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X126 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X127 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X128 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X129 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X130 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X131 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X132 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X133 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X134 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X135 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X136 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X138 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X139 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X141 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X142 a_n45858_n64215# Gnd sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X143 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X144 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X145 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X146 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X147 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X149 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X150 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X151 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X152 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X153 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X155 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X156 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X157 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X158 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X161 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X162 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X163 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X164 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X165 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X166 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X167 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X169 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X171 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X172 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X173 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X174 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X175 a_47_7088# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X176 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X177 Gnd Gnd a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X178 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X179 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X180 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X181 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X182 Gnd a_n45858_n24875# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X183 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X185 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X186 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X188 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X189 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D1 Gnd a_n45858_n24875# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X190 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X191 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X192 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X193 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X195 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X196 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X197 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X198 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X199 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X201 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X202 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X203 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X206 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X207 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X208 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X209 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D2 Gnd a_n45858_n64215# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X213 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X214 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X215 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X216 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X217 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X218 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X219 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X220 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X221 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X222 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X223 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X224 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X225 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X226 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X227 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X228 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X229 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X230 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X231 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X232 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X233 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X234 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X235 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X236 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X237 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X238 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X239 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X241 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X242 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X243 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X245 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X246 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X247 Gnd a_n45858_n24875# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X248 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X249 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X250 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X251 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X252 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X253 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X254 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X255 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X256 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X257 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X258 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X259 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X260 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X261 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X262 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X263 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X265 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X266 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X267 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R1 Vgg_1v2 a_n45858_n24875# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X268 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X269 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X270 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X271 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X272 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X273 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X274 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X275 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X276 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X277 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X278 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X279 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X280 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X281 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X282 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X283 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X284 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X285 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X286 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X287 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X288 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X289 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X290 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X291 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X292 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X293 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X294 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X295 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X296 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X297 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X298 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X299 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X300 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X301 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X302 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X303 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X304 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X305 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X306 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt MOM_capacitor in out gnd
.ends

