**.subckt MOM_capacitor in in_dummy out out_dummy
*.iopin in
*.iopin in_dummy
*.iopin out
*.iopin out_dummy
XR1 in in_dummy sky130_fd_pr__res_generic_m5 W=1.145 L=7.82 mult=1 m=1
XR2 out out_dummy sky130_fd_pr__res_generic_m5 W=1.145 L=7.82 mult=1 m=1
**.ends
** flattened .save nodes
.end
