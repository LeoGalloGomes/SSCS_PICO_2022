magic
tech sky130A
magscale 1 2
timestamp 1668378167
<< nwell >>
rect -50534 32812 -48746 33609
rect 2813 32812 4601 33609
<< pwell >>
rect -50485 32399 -48795 32681
rect -50499 32193 -48781 32399
rect 1997 32349 2343 32695
rect 2862 32399 4552 32681
rect 2848 32193 4566 32399
rect -50925 31845 -50579 32191
rect -42562 4611 -40628 5463
rect 66 4599 2000 5451
rect -42563 -5563 -40629 -4711
rect 78 -5589 2012 -4737
<< pmoslvt >>
rect -50401 32912 -50301 33312
rect -50243 32912 -50143 33312
rect -50085 32912 -49985 33312
rect -49927 32912 -49827 33312
rect -49769 32912 -49669 33312
rect -49611 32912 -49511 33312
rect -49453 32912 -49353 33312
rect -49295 32912 -49195 33312
rect -49137 32912 -49037 33312
rect -48979 32912 -48879 33312
rect 2946 32912 3046 33312
rect 3104 32912 3204 33312
rect 3262 32912 3362 33312
rect 3420 32912 3520 33312
rect 3578 32912 3678 33312
rect 3736 32912 3836 33312
rect 3894 32912 3994 33312
rect 4052 32912 4152 33312
rect 4210 32912 4310 33312
rect 4368 32912 4468 33312
<< nmoslvt >>
rect -50401 32455 -50301 32655
rect -50243 32455 -50143 32655
rect -50085 32455 -49985 32655
rect -49927 32455 -49827 32655
rect -49769 32455 -49669 32655
rect -49611 32455 -49511 32655
rect -49453 32455 -49353 32655
rect -49295 32455 -49195 32655
rect -49137 32455 -49037 32655
rect -48979 32455 -48879 32655
rect 2946 32455 3046 32655
rect 3104 32455 3204 32655
rect 3262 32455 3362 32655
rect 3420 32455 3520 32655
rect 3578 32455 3678 32655
rect 3736 32455 3836 32655
rect 3894 32455 3994 32655
rect 4052 32455 4152 32655
rect 4210 32455 4310 32655
rect 4368 32455 4468 32655
rect -42474 4637 -42444 5437
rect -42378 4637 -42348 5437
rect -42282 4637 -42252 5437
rect -42186 4637 -42156 5437
rect -42090 4637 -42060 5437
rect -41994 4637 -41964 5437
rect -41898 4637 -41868 5437
rect -41802 4637 -41772 5437
rect -41706 4637 -41676 5437
rect -41610 4637 -41580 5437
rect -41514 4637 -41484 5437
rect -41418 4637 -41388 5437
rect -41322 4637 -41292 5437
rect -41226 4637 -41196 5437
rect -41130 4637 -41100 5437
rect -41034 4637 -41004 5437
rect -40938 4637 -40908 5437
rect -40842 4637 -40812 5437
rect -40746 4637 -40716 5437
rect 154 4625 184 5425
rect 250 4625 280 5425
rect 346 4625 376 5425
rect 442 4625 472 5425
rect 538 4625 568 5425
rect 634 4625 664 5425
rect 730 4625 760 5425
rect 826 4625 856 5425
rect 922 4625 952 5425
rect 1018 4625 1048 5425
rect 1114 4625 1144 5425
rect 1210 4625 1240 5425
rect 1306 4625 1336 5425
rect 1402 4625 1432 5425
rect 1498 4625 1528 5425
rect 1594 4625 1624 5425
rect 1690 4625 1720 5425
rect 1786 4625 1816 5425
rect 1882 4625 1912 5425
rect -42475 -5537 -42445 -4737
rect -42379 -5537 -42349 -4737
rect -42283 -5537 -42253 -4737
rect -42187 -5537 -42157 -4737
rect -42091 -5537 -42061 -4737
rect -41995 -5537 -41965 -4737
rect -41899 -5537 -41869 -4737
rect -41803 -5537 -41773 -4737
rect -41707 -5537 -41677 -4737
rect -41611 -5537 -41581 -4737
rect -41515 -5537 -41485 -4737
rect -41419 -5537 -41389 -4737
rect -41323 -5537 -41293 -4737
rect -41227 -5537 -41197 -4737
rect -41131 -5537 -41101 -4737
rect -41035 -5537 -41005 -4737
rect -40939 -5537 -40909 -4737
rect -40843 -5537 -40813 -4737
rect -40747 -5537 -40717 -4737
rect 166 -5563 196 -4763
rect 262 -5563 292 -4763
rect 358 -5563 388 -4763
rect 454 -5563 484 -4763
rect 550 -5563 580 -4763
rect 646 -5563 676 -4763
rect 742 -5563 772 -4763
rect 838 -5563 868 -4763
rect 934 -5563 964 -4763
rect 1030 -5563 1060 -4763
rect 1126 -5563 1156 -4763
rect 1222 -5563 1252 -4763
rect 1318 -5563 1348 -4763
rect 1414 -5563 1444 -4763
rect 1510 -5563 1540 -4763
rect 1606 -5563 1636 -4763
rect 1702 -5563 1732 -4763
rect 1798 -5563 1828 -4763
rect 1894 -5563 1924 -4763
<< ndiff >>
rect -50459 32640 -50401 32655
rect -50459 32606 -50447 32640
rect -50413 32606 -50401 32640
rect -50459 32572 -50401 32606
rect -50459 32538 -50447 32572
rect -50413 32538 -50401 32572
rect -50459 32504 -50401 32538
rect -50459 32470 -50447 32504
rect -50413 32470 -50401 32504
rect -50459 32455 -50401 32470
rect -50301 32640 -50243 32655
rect -50301 32606 -50289 32640
rect -50255 32606 -50243 32640
rect -50301 32572 -50243 32606
rect -50301 32538 -50289 32572
rect -50255 32538 -50243 32572
rect -50301 32504 -50243 32538
rect -50301 32470 -50289 32504
rect -50255 32470 -50243 32504
rect -50301 32455 -50243 32470
rect -50143 32640 -50085 32655
rect -50143 32606 -50131 32640
rect -50097 32606 -50085 32640
rect -50143 32572 -50085 32606
rect -50143 32538 -50131 32572
rect -50097 32538 -50085 32572
rect -50143 32504 -50085 32538
rect -50143 32470 -50131 32504
rect -50097 32470 -50085 32504
rect -50143 32455 -50085 32470
rect -49985 32640 -49927 32655
rect -49985 32606 -49973 32640
rect -49939 32606 -49927 32640
rect -49985 32572 -49927 32606
rect -49985 32538 -49973 32572
rect -49939 32538 -49927 32572
rect -49985 32504 -49927 32538
rect -49985 32470 -49973 32504
rect -49939 32470 -49927 32504
rect -49985 32455 -49927 32470
rect -49827 32640 -49769 32655
rect -49827 32606 -49815 32640
rect -49781 32606 -49769 32640
rect -49827 32572 -49769 32606
rect -49827 32538 -49815 32572
rect -49781 32538 -49769 32572
rect -49827 32504 -49769 32538
rect -49827 32470 -49815 32504
rect -49781 32470 -49769 32504
rect -49827 32455 -49769 32470
rect -49669 32640 -49611 32655
rect -49669 32606 -49657 32640
rect -49623 32606 -49611 32640
rect -49669 32572 -49611 32606
rect -49669 32538 -49657 32572
rect -49623 32538 -49611 32572
rect -49669 32504 -49611 32538
rect -49669 32470 -49657 32504
rect -49623 32470 -49611 32504
rect -49669 32455 -49611 32470
rect -49511 32640 -49453 32655
rect -49511 32606 -49499 32640
rect -49465 32606 -49453 32640
rect -49511 32572 -49453 32606
rect -49511 32538 -49499 32572
rect -49465 32538 -49453 32572
rect -49511 32504 -49453 32538
rect -49511 32470 -49499 32504
rect -49465 32470 -49453 32504
rect -49511 32455 -49453 32470
rect -49353 32640 -49295 32655
rect -49353 32606 -49341 32640
rect -49307 32606 -49295 32640
rect -49353 32572 -49295 32606
rect -49353 32538 -49341 32572
rect -49307 32538 -49295 32572
rect -49353 32504 -49295 32538
rect -49353 32470 -49341 32504
rect -49307 32470 -49295 32504
rect -49353 32455 -49295 32470
rect -49195 32640 -49137 32655
rect -49195 32606 -49183 32640
rect -49149 32606 -49137 32640
rect -49195 32572 -49137 32606
rect -49195 32538 -49183 32572
rect -49149 32538 -49137 32572
rect -49195 32504 -49137 32538
rect -49195 32470 -49183 32504
rect -49149 32470 -49137 32504
rect -49195 32455 -49137 32470
rect -49037 32640 -48979 32655
rect -49037 32606 -49025 32640
rect -48991 32606 -48979 32640
rect -49037 32572 -48979 32606
rect -49037 32538 -49025 32572
rect -48991 32538 -48979 32572
rect -49037 32504 -48979 32538
rect -49037 32470 -49025 32504
rect -48991 32470 -48979 32504
rect -49037 32455 -48979 32470
rect -48879 32640 -48821 32655
rect -48879 32606 -48867 32640
rect -48833 32606 -48821 32640
rect -48879 32572 -48821 32606
rect -48879 32538 -48867 32572
rect -48833 32538 -48821 32572
rect -48879 32504 -48821 32538
rect -48879 32470 -48867 32504
rect -48833 32470 -48821 32504
rect -48879 32455 -48821 32470
rect 2888 32640 2946 32655
rect 2888 32606 2900 32640
rect 2934 32606 2946 32640
rect 2888 32572 2946 32606
rect 2888 32538 2900 32572
rect 2934 32538 2946 32572
rect 2888 32504 2946 32538
rect 2888 32470 2900 32504
rect 2934 32470 2946 32504
rect 2888 32455 2946 32470
rect 3046 32640 3104 32655
rect 3046 32606 3058 32640
rect 3092 32606 3104 32640
rect 3046 32572 3104 32606
rect 3046 32538 3058 32572
rect 3092 32538 3104 32572
rect 3046 32504 3104 32538
rect 3046 32470 3058 32504
rect 3092 32470 3104 32504
rect 3046 32455 3104 32470
rect 3204 32640 3262 32655
rect 3204 32606 3216 32640
rect 3250 32606 3262 32640
rect 3204 32572 3262 32606
rect 3204 32538 3216 32572
rect 3250 32538 3262 32572
rect 3204 32504 3262 32538
rect 3204 32470 3216 32504
rect 3250 32470 3262 32504
rect 3204 32455 3262 32470
rect 3362 32640 3420 32655
rect 3362 32606 3374 32640
rect 3408 32606 3420 32640
rect 3362 32572 3420 32606
rect 3362 32538 3374 32572
rect 3408 32538 3420 32572
rect 3362 32504 3420 32538
rect 3362 32470 3374 32504
rect 3408 32470 3420 32504
rect 3362 32455 3420 32470
rect 3520 32640 3578 32655
rect 3520 32606 3532 32640
rect 3566 32606 3578 32640
rect 3520 32572 3578 32606
rect 3520 32538 3532 32572
rect 3566 32538 3578 32572
rect 3520 32504 3578 32538
rect 3520 32470 3532 32504
rect 3566 32470 3578 32504
rect 3520 32455 3578 32470
rect 3678 32640 3736 32655
rect 3678 32606 3690 32640
rect 3724 32606 3736 32640
rect 3678 32572 3736 32606
rect 3678 32538 3690 32572
rect 3724 32538 3736 32572
rect 3678 32504 3736 32538
rect 3678 32470 3690 32504
rect 3724 32470 3736 32504
rect 3678 32455 3736 32470
rect 3836 32640 3894 32655
rect 3836 32606 3848 32640
rect 3882 32606 3894 32640
rect 3836 32572 3894 32606
rect 3836 32538 3848 32572
rect 3882 32538 3894 32572
rect 3836 32504 3894 32538
rect 3836 32470 3848 32504
rect 3882 32470 3894 32504
rect 3836 32455 3894 32470
rect 3994 32640 4052 32655
rect 3994 32606 4006 32640
rect 4040 32606 4052 32640
rect 3994 32572 4052 32606
rect 3994 32538 4006 32572
rect 4040 32538 4052 32572
rect 3994 32504 4052 32538
rect 3994 32470 4006 32504
rect 4040 32470 4052 32504
rect 3994 32455 4052 32470
rect 4152 32640 4210 32655
rect 4152 32606 4164 32640
rect 4198 32606 4210 32640
rect 4152 32572 4210 32606
rect 4152 32538 4164 32572
rect 4198 32538 4210 32572
rect 4152 32504 4210 32538
rect 4152 32470 4164 32504
rect 4198 32470 4210 32504
rect 4152 32455 4210 32470
rect 4310 32640 4368 32655
rect 4310 32606 4322 32640
rect 4356 32606 4368 32640
rect 4310 32572 4368 32606
rect 4310 32538 4322 32572
rect 4356 32538 4368 32572
rect 4310 32504 4368 32538
rect 4310 32470 4322 32504
rect 4356 32470 4368 32504
rect 4310 32455 4368 32470
rect 4468 32640 4526 32655
rect 4468 32606 4480 32640
rect 4514 32606 4526 32640
rect 4468 32572 4526 32606
rect 4468 32538 4480 32572
rect 4514 32538 4526 32572
rect 4468 32504 4526 32538
rect 4468 32470 4480 32504
rect 4514 32470 4526 32504
rect 4468 32455 4526 32470
rect -42536 5394 -42474 5437
rect -42536 5360 -42524 5394
rect -42490 5360 -42474 5394
rect -42536 5326 -42474 5360
rect -42536 5292 -42524 5326
rect -42490 5292 -42474 5326
rect -42536 5258 -42474 5292
rect -42536 5224 -42524 5258
rect -42490 5224 -42474 5258
rect -42536 5190 -42474 5224
rect -42536 5156 -42524 5190
rect -42490 5156 -42474 5190
rect -42536 5122 -42474 5156
rect -42536 5088 -42524 5122
rect -42490 5088 -42474 5122
rect -42536 5054 -42474 5088
rect -42536 5020 -42524 5054
rect -42490 5020 -42474 5054
rect -42536 4986 -42474 5020
rect -42536 4952 -42524 4986
rect -42490 4952 -42474 4986
rect -42536 4918 -42474 4952
rect -42536 4884 -42524 4918
rect -42490 4884 -42474 4918
rect -42536 4850 -42474 4884
rect -42536 4816 -42524 4850
rect -42490 4816 -42474 4850
rect -42536 4782 -42474 4816
rect -42536 4748 -42524 4782
rect -42490 4748 -42474 4782
rect -42536 4714 -42474 4748
rect -42536 4680 -42524 4714
rect -42490 4680 -42474 4714
rect -42536 4637 -42474 4680
rect -42444 5394 -42378 5437
rect -42444 5360 -42428 5394
rect -42394 5360 -42378 5394
rect -42444 5326 -42378 5360
rect -42444 5292 -42428 5326
rect -42394 5292 -42378 5326
rect -42444 5258 -42378 5292
rect -42444 5224 -42428 5258
rect -42394 5224 -42378 5258
rect -42444 5190 -42378 5224
rect -42444 5156 -42428 5190
rect -42394 5156 -42378 5190
rect -42444 5122 -42378 5156
rect -42444 5088 -42428 5122
rect -42394 5088 -42378 5122
rect -42444 5054 -42378 5088
rect -42444 5020 -42428 5054
rect -42394 5020 -42378 5054
rect -42444 4986 -42378 5020
rect -42444 4952 -42428 4986
rect -42394 4952 -42378 4986
rect -42444 4918 -42378 4952
rect -42444 4884 -42428 4918
rect -42394 4884 -42378 4918
rect -42444 4850 -42378 4884
rect -42444 4816 -42428 4850
rect -42394 4816 -42378 4850
rect -42444 4782 -42378 4816
rect -42444 4748 -42428 4782
rect -42394 4748 -42378 4782
rect -42444 4714 -42378 4748
rect -42444 4680 -42428 4714
rect -42394 4680 -42378 4714
rect -42444 4637 -42378 4680
rect -42348 5394 -42282 5437
rect -42348 5360 -42332 5394
rect -42298 5360 -42282 5394
rect -42348 5326 -42282 5360
rect -42348 5292 -42332 5326
rect -42298 5292 -42282 5326
rect -42348 5258 -42282 5292
rect -42348 5224 -42332 5258
rect -42298 5224 -42282 5258
rect -42348 5190 -42282 5224
rect -42348 5156 -42332 5190
rect -42298 5156 -42282 5190
rect -42348 5122 -42282 5156
rect -42348 5088 -42332 5122
rect -42298 5088 -42282 5122
rect -42348 5054 -42282 5088
rect -42348 5020 -42332 5054
rect -42298 5020 -42282 5054
rect -42348 4986 -42282 5020
rect -42348 4952 -42332 4986
rect -42298 4952 -42282 4986
rect -42348 4918 -42282 4952
rect -42348 4884 -42332 4918
rect -42298 4884 -42282 4918
rect -42348 4850 -42282 4884
rect -42348 4816 -42332 4850
rect -42298 4816 -42282 4850
rect -42348 4782 -42282 4816
rect -42348 4748 -42332 4782
rect -42298 4748 -42282 4782
rect -42348 4714 -42282 4748
rect -42348 4680 -42332 4714
rect -42298 4680 -42282 4714
rect -42348 4637 -42282 4680
rect -42252 5394 -42186 5437
rect -42252 5360 -42236 5394
rect -42202 5360 -42186 5394
rect -42252 5326 -42186 5360
rect -42252 5292 -42236 5326
rect -42202 5292 -42186 5326
rect -42252 5258 -42186 5292
rect -42252 5224 -42236 5258
rect -42202 5224 -42186 5258
rect -42252 5190 -42186 5224
rect -42252 5156 -42236 5190
rect -42202 5156 -42186 5190
rect -42252 5122 -42186 5156
rect -42252 5088 -42236 5122
rect -42202 5088 -42186 5122
rect -42252 5054 -42186 5088
rect -42252 5020 -42236 5054
rect -42202 5020 -42186 5054
rect -42252 4986 -42186 5020
rect -42252 4952 -42236 4986
rect -42202 4952 -42186 4986
rect -42252 4918 -42186 4952
rect -42252 4884 -42236 4918
rect -42202 4884 -42186 4918
rect -42252 4850 -42186 4884
rect -42252 4816 -42236 4850
rect -42202 4816 -42186 4850
rect -42252 4782 -42186 4816
rect -42252 4748 -42236 4782
rect -42202 4748 -42186 4782
rect -42252 4714 -42186 4748
rect -42252 4680 -42236 4714
rect -42202 4680 -42186 4714
rect -42252 4637 -42186 4680
rect -42156 5394 -42090 5437
rect -42156 5360 -42140 5394
rect -42106 5360 -42090 5394
rect -42156 5326 -42090 5360
rect -42156 5292 -42140 5326
rect -42106 5292 -42090 5326
rect -42156 5258 -42090 5292
rect -42156 5224 -42140 5258
rect -42106 5224 -42090 5258
rect -42156 5190 -42090 5224
rect -42156 5156 -42140 5190
rect -42106 5156 -42090 5190
rect -42156 5122 -42090 5156
rect -42156 5088 -42140 5122
rect -42106 5088 -42090 5122
rect -42156 5054 -42090 5088
rect -42156 5020 -42140 5054
rect -42106 5020 -42090 5054
rect -42156 4986 -42090 5020
rect -42156 4952 -42140 4986
rect -42106 4952 -42090 4986
rect -42156 4918 -42090 4952
rect -42156 4884 -42140 4918
rect -42106 4884 -42090 4918
rect -42156 4850 -42090 4884
rect -42156 4816 -42140 4850
rect -42106 4816 -42090 4850
rect -42156 4782 -42090 4816
rect -42156 4748 -42140 4782
rect -42106 4748 -42090 4782
rect -42156 4714 -42090 4748
rect -42156 4680 -42140 4714
rect -42106 4680 -42090 4714
rect -42156 4637 -42090 4680
rect -42060 5394 -41994 5437
rect -42060 5360 -42044 5394
rect -42010 5360 -41994 5394
rect -42060 5326 -41994 5360
rect -42060 5292 -42044 5326
rect -42010 5292 -41994 5326
rect -42060 5258 -41994 5292
rect -42060 5224 -42044 5258
rect -42010 5224 -41994 5258
rect -42060 5190 -41994 5224
rect -42060 5156 -42044 5190
rect -42010 5156 -41994 5190
rect -42060 5122 -41994 5156
rect -42060 5088 -42044 5122
rect -42010 5088 -41994 5122
rect -42060 5054 -41994 5088
rect -42060 5020 -42044 5054
rect -42010 5020 -41994 5054
rect -42060 4986 -41994 5020
rect -42060 4952 -42044 4986
rect -42010 4952 -41994 4986
rect -42060 4918 -41994 4952
rect -42060 4884 -42044 4918
rect -42010 4884 -41994 4918
rect -42060 4850 -41994 4884
rect -42060 4816 -42044 4850
rect -42010 4816 -41994 4850
rect -42060 4782 -41994 4816
rect -42060 4748 -42044 4782
rect -42010 4748 -41994 4782
rect -42060 4714 -41994 4748
rect -42060 4680 -42044 4714
rect -42010 4680 -41994 4714
rect -42060 4637 -41994 4680
rect -41964 5394 -41898 5437
rect -41964 5360 -41948 5394
rect -41914 5360 -41898 5394
rect -41964 5326 -41898 5360
rect -41964 5292 -41948 5326
rect -41914 5292 -41898 5326
rect -41964 5258 -41898 5292
rect -41964 5224 -41948 5258
rect -41914 5224 -41898 5258
rect -41964 5190 -41898 5224
rect -41964 5156 -41948 5190
rect -41914 5156 -41898 5190
rect -41964 5122 -41898 5156
rect -41964 5088 -41948 5122
rect -41914 5088 -41898 5122
rect -41964 5054 -41898 5088
rect -41964 5020 -41948 5054
rect -41914 5020 -41898 5054
rect -41964 4986 -41898 5020
rect -41964 4952 -41948 4986
rect -41914 4952 -41898 4986
rect -41964 4918 -41898 4952
rect -41964 4884 -41948 4918
rect -41914 4884 -41898 4918
rect -41964 4850 -41898 4884
rect -41964 4816 -41948 4850
rect -41914 4816 -41898 4850
rect -41964 4782 -41898 4816
rect -41964 4748 -41948 4782
rect -41914 4748 -41898 4782
rect -41964 4714 -41898 4748
rect -41964 4680 -41948 4714
rect -41914 4680 -41898 4714
rect -41964 4637 -41898 4680
rect -41868 5394 -41802 5437
rect -41868 5360 -41852 5394
rect -41818 5360 -41802 5394
rect -41868 5326 -41802 5360
rect -41868 5292 -41852 5326
rect -41818 5292 -41802 5326
rect -41868 5258 -41802 5292
rect -41868 5224 -41852 5258
rect -41818 5224 -41802 5258
rect -41868 5190 -41802 5224
rect -41868 5156 -41852 5190
rect -41818 5156 -41802 5190
rect -41868 5122 -41802 5156
rect -41868 5088 -41852 5122
rect -41818 5088 -41802 5122
rect -41868 5054 -41802 5088
rect -41868 5020 -41852 5054
rect -41818 5020 -41802 5054
rect -41868 4986 -41802 5020
rect -41868 4952 -41852 4986
rect -41818 4952 -41802 4986
rect -41868 4918 -41802 4952
rect -41868 4884 -41852 4918
rect -41818 4884 -41802 4918
rect -41868 4850 -41802 4884
rect -41868 4816 -41852 4850
rect -41818 4816 -41802 4850
rect -41868 4782 -41802 4816
rect -41868 4748 -41852 4782
rect -41818 4748 -41802 4782
rect -41868 4714 -41802 4748
rect -41868 4680 -41852 4714
rect -41818 4680 -41802 4714
rect -41868 4637 -41802 4680
rect -41772 5394 -41706 5437
rect -41772 5360 -41756 5394
rect -41722 5360 -41706 5394
rect -41772 5326 -41706 5360
rect -41772 5292 -41756 5326
rect -41722 5292 -41706 5326
rect -41772 5258 -41706 5292
rect -41772 5224 -41756 5258
rect -41722 5224 -41706 5258
rect -41772 5190 -41706 5224
rect -41772 5156 -41756 5190
rect -41722 5156 -41706 5190
rect -41772 5122 -41706 5156
rect -41772 5088 -41756 5122
rect -41722 5088 -41706 5122
rect -41772 5054 -41706 5088
rect -41772 5020 -41756 5054
rect -41722 5020 -41706 5054
rect -41772 4986 -41706 5020
rect -41772 4952 -41756 4986
rect -41722 4952 -41706 4986
rect -41772 4918 -41706 4952
rect -41772 4884 -41756 4918
rect -41722 4884 -41706 4918
rect -41772 4850 -41706 4884
rect -41772 4816 -41756 4850
rect -41722 4816 -41706 4850
rect -41772 4782 -41706 4816
rect -41772 4748 -41756 4782
rect -41722 4748 -41706 4782
rect -41772 4714 -41706 4748
rect -41772 4680 -41756 4714
rect -41722 4680 -41706 4714
rect -41772 4637 -41706 4680
rect -41676 5394 -41610 5437
rect -41676 5360 -41660 5394
rect -41626 5360 -41610 5394
rect -41676 5326 -41610 5360
rect -41676 5292 -41660 5326
rect -41626 5292 -41610 5326
rect -41676 5258 -41610 5292
rect -41676 5224 -41660 5258
rect -41626 5224 -41610 5258
rect -41676 5190 -41610 5224
rect -41676 5156 -41660 5190
rect -41626 5156 -41610 5190
rect -41676 5122 -41610 5156
rect -41676 5088 -41660 5122
rect -41626 5088 -41610 5122
rect -41676 5054 -41610 5088
rect -41676 5020 -41660 5054
rect -41626 5020 -41610 5054
rect -41676 4986 -41610 5020
rect -41676 4952 -41660 4986
rect -41626 4952 -41610 4986
rect -41676 4918 -41610 4952
rect -41676 4884 -41660 4918
rect -41626 4884 -41610 4918
rect -41676 4850 -41610 4884
rect -41676 4816 -41660 4850
rect -41626 4816 -41610 4850
rect -41676 4782 -41610 4816
rect -41676 4748 -41660 4782
rect -41626 4748 -41610 4782
rect -41676 4714 -41610 4748
rect -41676 4680 -41660 4714
rect -41626 4680 -41610 4714
rect -41676 4637 -41610 4680
rect -41580 5394 -41514 5437
rect -41580 5360 -41564 5394
rect -41530 5360 -41514 5394
rect -41580 5326 -41514 5360
rect -41580 5292 -41564 5326
rect -41530 5292 -41514 5326
rect -41580 5258 -41514 5292
rect -41580 5224 -41564 5258
rect -41530 5224 -41514 5258
rect -41580 5190 -41514 5224
rect -41580 5156 -41564 5190
rect -41530 5156 -41514 5190
rect -41580 5122 -41514 5156
rect -41580 5088 -41564 5122
rect -41530 5088 -41514 5122
rect -41580 5054 -41514 5088
rect -41580 5020 -41564 5054
rect -41530 5020 -41514 5054
rect -41580 4986 -41514 5020
rect -41580 4952 -41564 4986
rect -41530 4952 -41514 4986
rect -41580 4918 -41514 4952
rect -41580 4884 -41564 4918
rect -41530 4884 -41514 4918
rect -41580 4850 -41514 4884
rect -41580 4816 -41564 4850
rect -41530 4816 -41514 4850
rect -41580 4782 -41514 4816
rect -41580 4748 -41564 4782
rect -41530 4748 -41514 4782
rect -41580 4714 -41514 4748
rect -41580 4680 -41564 4714
rect -41530 4680 -41514 4714
rect -41580 4637 -41514 4680
rect -41484 5394 -41418 5437
rect -41484 5360 -41468 5394
rect -41434 5360 -41418 5394
rect -41484 5326 -41418 5360
rect -41484 5292 -41468 5326
rect -41434 5292 -41418 5326
rect -41484 5258 -41418 5292
rect -41484 5224 -41468 5258
rect -41434 5224 -41418 5258
rect -41484 5190 -41418 5224
rect -41484 5156 -41468 5190
rect -41434 5156 -41418 5190
rect -41484 5122 -41418 5156
rect -41484 5088 -41468 5122
rect -41434 5088 -41418 5122
rect -41484 5054 -41418 5088
rect -41484 5020 -41468 5054
rect -41434 5020 -41418 5054
rect -41484 4986 -41418 5020
rect -41484 4952 -41468 4986
rect -41434 4952 -41418 4986
rect -41484 4918 -41418 4952
rect -41484 4884 -41468 4918
rect -41434 4884 -41418 4918
rect -41484 4850 -41418 4884
rect -41484 4816 -41468 4850
rect -41434 4816 -41418 4850
rect -41484 4782 -41418 4816
rect -41484 4748 -41468 4782
rect -41434 4748 -41418 4782
rect -41484 4714 -41418 4748
rect -41484 4680 -41468 4714
rect -41434 4680 -41418 4714
rect -41484 4637 -41418 4680
rect -41388 5394 -41322 5437
rect -41388 5360 -41372 5394
rect -41338 5360 -41322 5394
rect -41388 5326 -41322 5360
rect -41388 5292 -41372 5326
rect -41338 5292 -41322 5326
rect -41388 5258 -41322 5292
rect -41388 5224 -41372 5258
rect -41338 5224 -41322 5258
rect -41388 5190 -41322 5224
rect -41388 5156 -41372 5190
rect -41338 5156 -41322 5190
rect -41388 5122 -41322 5156
rect -41388 5088 -41372 5122
rect -41338 5088 -41322 5122
rect -41388 5054 -41322 5088
rect -41388 5020 -41372 5054
rect -41338 5020 -41322 5054
rect -41388 4986 -41322 5020
rect -41388 4952 -41372 4986
rect -41338 4952 -41322 4986
rect -41388 4918 -41322 4952
rect -41388 4884 -41372 4918
rect -41338 4884 -41322 4918
rect -41388 4850 -41322 4884
rect -41388 4816 -41372 4850
rect -41338 4816 -41322 4850
rect -41388 4782 -41322 4816
rect -41388 4748 -41372 4782
rect -41338 4748 -41322 4782
rect -41388 4714 -41322 4748
rect -41388 4680 -41372 4714
rect -41338 4680 -41322 4714
rect -41388 4637 -41322 4680
rect -41292 5394 -41226 5437
rect -41292 5360 -41276 5394
rect -41242 5360 -41226 5394
rect -41292 5326 -41226 5360
rect -41292 5292 -41276 5326
rect -41242 5292 -41226 5326
rect -41292 5258 -41226 5292
rect -41292 5224 -41276 5258
rect -41242 5224 -41226 5258
rect -41292 5190 -41226 5224
rect -41292 5156 -41276 5190
rect -41242 5156 -41226 5190
rect -41292 5122 -41226 5156
rect -41292 5088 -41276 5122
rect -41242 5088 -41226 5122
rect -41292 5054 -41226 5088
rect -41292 5020 -41276 5054
rect -41242 5020 -41226 5054
rect -41292 4986 -41226 5020
rect -41292 4952 -41276 4986
rect -41242 4952 -41226 4986
rect -41292 4918 -41226 4952
rect -41292 4884 -41276 4918
rect -41242 4884 -41226 4918
rect -41292 4850 -41226 4884
rect -41292 4816 -41276 4850
rect -41242 4816 -41226 4850
rect -41292 4782 -41226 4816
rect -41292 4748 -41276 4782
rect -41242 4748 -41226 4782
rect -41292 4714 -41226 4748
rect -41292 4680 -41276 4714
rect -41242 4680 -41226 4714
rect -41292 4637 -41226 4680
rect -41196 5394 -41130 5437
rect -41196 5360 -41180 5394
rect -41146 5360 -41130 5394
rect -41196 5326 -41130 5360
rect -41196 5292 -41180 5326
rect -41146 5292 -41130 5326
rect -41196 5258 -41130 5292
rect -41196 5224 -41180 5258
rect -41146 5224 -41130 5258
rect -41196 5190 -41130 5224
rect -41196 5156 -41180 5190
rect -41146 5156 -41130 5190
rect -41196 5122 -41130 5156
rect -41196 5088 -41180 5122
rect -41146 5088 -41130 5122
rect -41196 5054 -41130 5088
rect -41196 5020 -41180 5054
rect -41146 5020 -41130 5054
rect -41196 4986 -41130 5020
rect -41196 4952 -41180 4986
rect -41146 4952 -41130 4986
rect -41196 4918 -41130 4952
rect -41196 4884 -41180 4918
rect -41146 4884 -41130 4918
rect -41196 4850 -41130 4884
rect -41196 4816 -41180 4850
rect -41146 4816 -41130 4850
rect -41196 4782 -41130 4816
rect -41196 4748 -41180 4782
rect -41146 4748 -41130 4782
rect -41196 4714 -41130 4748
rect -41196 4680 -41180 4714
rect -41146 4680 -41130 4714
rect -41196 4637 -41130 4680
rect -41100 5394 -41034 5437
rect -41100 5360 -41084 5394
rect -41050 5360 -41034 5394
rect -41100 5326 -41034 5360
rect -41100 5292 -41084 5326
rect -41050 5292 -41034 5326
rect -41100 5258 -41034 5292
rect -41100 5224 -41084 5258
rect -41050 5224 -41034 5258
rect -41100 5190 -41034 5224
rect -41100 5156 -41084 5190
rect -41050 5156 -41034 5190
rect -41100 5122 -41034 5156
rect -41100 5088 -41084 5122
rect -41050 5088 -41034 5122
rect -41100 5054 -41034 5088
rect -41100 5020 -41084 5054
rect -41050 5020 -41034 5054
rect -41100 4986 -41034 5020
rect -41100 4952 -41084 4986
rect -41050 4952 -41034 4986
rect -41100 4918 -41034 4952
rect -41100 4884 -41084 4918
rect -41050 4884 -41034 4918
rect -41100 4850 -41034 4884
rect -41100 4816 -41084 4850
rect -41050 4816 -41034 4850
rect -41100 4782 -41034 4816
rect -41100 4748 -41084 4782
rect -41050 4748 -41034 4782
rect -41100 4714 -41034 4748
rect -41100 4680 -41084 4714
rect -41050 4680 -41034 4714
rect -41100 4637 -41034 4680
rect -41004 5394 -40938 5437
rect -41004 5360 -40988 5394
rect -40954 5360 -40938 5394
rect -41004 5326 -40938 5360
rect -41004 5292 -40988 5326
rect -40954 5292 -40938 5326
rect -41004 5258 -40938 5292
rect -41004 5224 -40988 5258
rect -40954 5224 -40938 5258
rect -41004 5190 -40938 5224
rect -41004 5156 -40988 5190
rect -40954 5156 -40938 5190
rect -41004 5122 -40938 5156
rect -41004 5088 -40988 5122
rect -40954 5088 -40938 5122
rect -41004 5054 -40938 5088
rect -41004 5020 -40988 5054
rect -40954 5020 -40938 5054
rect -41004 4986 -40938 5020
rect -41004 4952 -40988 4986
rect -40954 4952 -40938 4986
rect -41004 4918 -40938 4952
rect -41004 4884 -40988 4918
rect -40954 4884 -40938 4918
rect -41004 4850 -40938 4884
rect -41004 4816 -40988 4850
rect -40954 4816 -40938 4850
rect -41004 4782 -40938 4816
rect -41004 4748 -40988 4782
rect -40954 4748 -40938 4782
rect -41004 4714 -40938 4748
rect -41004 4680 -40988 4714
rect -40954 4680 -40938 4714
rect -41004 4637 -40938 4680
rect -40908 5394 -40842 5437
rect -40908 5360 -40892 5394
rect -40858 5360 -40842 5394
rect -40908 5326 -40842 5360
rect -40908 5292 -40892 5326
rect -40858 5292 -40842 5326
rect -40908 5258 -40842 5292
rect -40908 5224 -40892 5258
rect -40858 5224 -40842 5258
rect -40908 5190 -40842 5224
rect -40908 5156 -40892 5190
rect -40858 5156 -40842 5190
rect -40908 5122 -40842 5156
rect -40908 5088 -40892 5122
rect -40858 5088 -40842 5122
rect -40908 5054 -40842 5088
rect -40908 5020 -40892 5054
rect -40858 5020 -40842 5054
rect -40908 4986 -40842 5020
rect -40908 4952 -40892 4986
rect -40858 4952 -40842 4986
rect -40908 4918 -40842 4952
rect -40908 4884 -40892 4918
rect -40858 4884 -40842 4918
rect -40908 4850 -40842 4884
rect -40908 4816 -40892 4850
rect -40858 4816 -40842 4850
rect -40908 4782 -40842 4816
rect -40908 4748 -40892 4782
rect -40858 4748 -40842 4782
rect -40908 4714 -40842 4748
rect -40908 4680 -40892 4714
rect -40858 4680 -40842 4714
rect -40908 4637 -40842 4680
rect -40812 5394 -40746 5437
rect -40812 5360 -40796 5394
rect -40762 5360 -40746 5394
rect -40812 5326 -40746 5360
rect -40812 5292 -40796 5326
rect -40762 5292 -40746 5326
rect -40812 5258 -40746 5292
rect -40812 5224 -40796 5258
rect -40762 5224 -40746 5258
rect -40812 5190 -40746 5224
rect -40812 5156 -40796 5190
rect -40762 5156 -40746 5190
rect -40812 5122 -40746 5156
rect -40812 5088 -40796 5122
rect -40762 5088 -40746 5122
rect -40812 5054 -40746 5088
rect -40812 5020 -40796 5054
rect -40762 5020 -40746 5054
rect -40812 4986 -40746 5020
rect -40812 4952 -40796 4986
rect -40762 4952 -40746 4986
rect -40812 4918 -40746 4952
rect -40812 4884 -40796 4918
rect -40762 4884 -40746 4918
rect -40812 4850 -40746 4884
rect -40812 4816 -40796 4850
rect -40762 4816 -40746 4850
rect -40812 4782 -40746 4816
rect -40812 4748 -40796 4782
rect -40762 4748 -40746 4782
rect -40812 4714 -40746 4748
rect -40812 4680 -40796 4714
rect -40762 4680 -40746 4714
rect -40812 4637 -40746 4680
rect -40716 5394 -40654 5437
rect -40716 5360 -40700 5394
rect -40666 5360 -40654 5394
rect -40716 5326 -40654 5360
rect -40716 5292 -40700 5326
rect -40666 5292 -40654 5326
rect -40716 5258 -40654 5292
rect -40716 5224 -40700 5258
rect -40666 5224 -40654 5258
rect -40716 5190 -40654 5224
rect -40716 5156 -40700 5190
rect -40666 5156 -40654 5190
rect -40716 5122 -40654 5156
rect -40716 5088 -40700 5122
rect -40666 5088 -40654 5122
rect -40716 5054 -40654 5088
rect -40716 5020 -40700 5054
rect -40666 5020 -40654 5054
rect -40716 4986 -40654 5020
rect -40716 4952 -40700 4986
rect -40666 4952 -40654 4986
rect -40716 4918 -40654 4952
rect -40716 4884 -40700 4918
rect -40666 4884 -40654 4918
rect -40716 4850 -40654 4884
rect -40716 4816 -40700 4850
rect -40666 4816 -40654 4850
rect -40716 4782 -40654 4816
rect -40716 4748 -40700 4782
rect -40666 4748 -40654 4782
rect -40716 4714 -40654 4748
rect -40716 4680 -40700 4714
rect -40666 4680 -40654 4714
rect -40716 4637 -40654 4680
rect 92 5382 154 5425
rect 92 5348 104 5382
rect 138 5348 154 5382
rect 92 5314 154 5348
rect 92 5280 104 5314
rect 138 5280 154 5314
rect 92 5246 154 5280
rect 92 5212 104 5246
rect 138 5212 154 5246
rect 92 5178 154 5212
rect 92 5144 104 5178
rect 138 5144 154 5178
rect 92 5110 154 5144
rect 92 5076 104 5110
rect 138 5076 154 5110
rect 92 5042 154 5076
rect 92 5008 104 5042
rect 138 5008 154 5042
rect 92 4974 154 5008
rect 92 4940 104 4974
rect 138 4940 154 4974
rect 92 4906 154 4940
rect 92 4872 104 4906
rect 138 4872 154 4906
rect 92 4838 154 4872
rect 92 4804 104 4838
rect 138 4804 154 4838
rect 92 4770 154 4804
rect 92 4736 104 4770
rect 138 4736 154 4770
rect 92 4702 154 4736
rect 92 4668 104 4702
rect 138 4668 154 4702
rect 92 4625 154 4668
rect 184 5382 250 5425
rect 184 5348 200 5382
rect 234 5348 250 5382
rect 184 5314 250 5348
rect 184 5280 200 5314
rect 234 5280 250 5314
rect 184 5246 250 5280
rect 184 5212 200 5246
rect 234 5212 250 5246
rect 184 5178 250 5212
rect 184 5144 200 5178
rect 234 5144 250 5178
rect 184 5110 250 5144
rect 184 5076 200 5110
rect 234 5076 250 5110
rect 184 5042 250 5076
rect 184 5008 200 5042
rect 234 5008 250 5042
rect 184 4974 250 5008
rect 184 4940 200 4974
rect 234 4940 250 4974
rect 184 4906 250 4940
rect 184 4872 200 4906
rect 234 4872 250 4906
rect 184 4838 250 4872
rect 184 4804 200 4838
rect 234 4804 250 4838
rect 184 4770 250 4804
rect 184 4736 200 4770
rect 234 4736 250 4770
rect 184 4702 250 4736
rect 184 4668 200 4702
rect 234 4668 250 4702
rect 184 4625 250 4668
rect 280 5382 346 5425
rect 280 5348 296 5382
rect 330 5348 346 5382
rect 280 5314 346 5348
rect 280 5280 296 5314
rect 330 5280 346 5314
rect 280 5246 346 5280
rect 280 5212 296 5246
rect 330 5212 346 5246
rect 280 5178 346 5212
rect 280 5144 296 5178
rect 330 5144 346 5178
rect 280 5110 346 5144
rect 280 5076 296 5110
rect 330 5076 346 5110
rect 280 5042 346 5076
rect 280 5008 296 5042
rect 330 5008 346 5042
rect 280 4974 346 5008
rect 280 4940 296 4974
rect 330 4940 346 4974
rect 280 4906 346 4940
rect 280 4872 296 4906
rect 330 4872 346 4906
rect 280 4838 346 4872
rect 280 4804 296 4838
rect 330 4804 346 4838
rect 280 4770 346 4804
rect 280 4736 296 4770
rect 330 4736 346 4770
rect 280 4702 346 4736
rect 280 4668 296 4702
rect 330 4668 346 4702
rect 280 4625 346 4668
rect 376 5382 442 5425
rect 376 5348 392 5382
rect 426 5348 442 5382
rect 376 5314 442 5348
rect 376 5280 392 5314
rect 426 5280 442 5314
rect 376 5246 442 5280
rect 376 5212 392 5246
rect 426 5212 442 5246
rect 376 5178 442 5212
rect 376 5144 392 5178
rect 426 5144 442 5178
rect 376 5110 442 5144
rect 376 5076 392 5110
rect 426 5076 442 5110
rect 376 5042 442 5076
rect 376 5008 392 5042
rect 426 5008 442 5042
rect 376 4974 442 5008
rect 376 4940 392 4974
rect 426 4940 442 4974
rect 376 4906 442 4940
rect 376 4872 392 4906
rect 426 4872 442 4906
rect 376 4838 442 4872
rect 376 4804 392 4838
rect 426 4804 442 4838
rect 376 4770 442 4804
rect 376 4736 392 4770
rect 426 4736 442 4770
rect 376 4702 442 4736
rect 376 4668 392 4702
rect 426 4668 442 4702
rect 376 4625 442 4668
rect 472 5382 538 5425
rect 472 5348 488 5382
rect 522 5348 538 5382
rect 472 5314 538 5348
rect 472 5280 488 5314
rect 522 5280 538 5314
rect 472 5246 538 5280
rect 472 5212 488 5246
rect 522 5212 538 5246
rect 472 5178 538 5212
rect 472 5144 488 5178
rect 522 5144 538 5178
rect 472 5110 538 5144
rect 472 5076 488 5110
rect 522 5076 538 5110
rect 472 5042 538 5076
rect 472 5008 488 5042
rect 522 5008 538 5042
rect 472 4974 538 5008
rect 472 4940 488 4974
rect 522 4940 538 4974
rect 472 4906 538 4940
rect 472 4872 488 4906
rect 522 4872 538 4906
rect 472 4838 538 4872
rect 472 4804 488 4838
rect 522 4804 538 4838
rect 472 4770 538 4804
rect 472 4736 488 4770
rect 522 4736 538 4770
rect 472 4702 538 4736
rect 472 4668 488 4702
rect 522 4668 538 4702
rect 472 4625 538 4668
rect 568 5382 634 5425
rect 568 5348 584 5382
rect 618 5348 634 5382
rect 568 5314 634 5348
rect 568 5280 584 5314
rect 618 5280 634 5314
rect 568 5246 634 5280
rect 568 5212 584 5246
rect 618 5212 634 5246
rect 568 5178 634 5212
rect 568 5144 584 5178
rect 618 5144 634 5178
rect 568 5110 634 5144
rect 568 5076 584 5110
rect 618 5076 634 5110
rect 568 5042 634 5076
rect 568 5008 584 5042
rect 618 5008 634 5042
rect 568 4974 634 5008
rect 568 4940 584 4974
rect 618 4940 634 4974
rect 568 4906 634 4940
rect 568 4872 584 4906
rect 618 4872 634 4906
rect 568 4838 634 4872
rect 568 4804 584 4838
rect 618 4804 634 4838
rect 568 4770 634 4804
rect 568 4736 584 4770
rect 618 4736 634 4770
rect 568 4702 634 4736
rect 568 4668 584 4702
rect 618 4668 634 4702
rect 568 4625 634 4668
rect 664 5382 730 5425
rect 664 5348 680 5382
rect 714 5348 730 5382
rect 664 5314 730 5348
rect 664 5280 680 5314
rect 714 5280 730 5314
rect 664 5246 730 5280
rect 664 5212 680 5246
rect 714 5212 730 5246
rect 664 5178 730 5212
rect 664 5144 680 5178
rect 714 5144 730 5178
rect 664 5110 730 5144
rect 664 5076 680 5110
rect 714 5076 730 5110
rect 664 5042 730 5076
rect 664 5008 680 5042
rect 714 5008 730 5042
rect 664 4974 730 5008
rect 664 4940 680 4974
rect 714 4940 730 4974
rect 664 4906 730 4940
rect 664 4872 680 4906
rect 714 4872 730 4906
rect 664 4838 730 4872
rect 664 4804 680 4838
rect 714 4804 730 4838
rect 664 4770 730 4804
rect 664 4736 680 4770
rect 714 4736 730 4770
rect 664 4702 730 4736
rect 664 4668 680 4702
rect 714 4668 730 4702
rect 664 4625 730 4668
rect 760 5382 826 5425
rect 760 5348 776 5382
rect 810 5348 826 5382
rect 760 5314 826 5348
rect 760 5280 776 5314
rect 810 5280 826 5314
rect 760 5246 826 5280
rect 760 5212 776 5246
rect 810 5212 826 5246
rect 760 5178 826 5212
rect 760 5144 776 5178
rect 810 5144 826 5178
rect 760 5110 826 5144
rect 760 5076 776 5110
rect 810 5076 826 5110
rect 760 5042 826 5076
rect 760 5008 776 5042
rect 810 5008 826 5042
rect 760 4974 826 5008
rect 760 4940 776 4974
rect 810 4940 826 4974
rect 760 4906 826 4940
rect 760 4872 776 4906
rect 810 4872 826 4906
rect 760 4838 826 4872
rect 760 4804 776 4838
rect 810 4804 826 4838
rect 760 4770 826 4804
rect 760 4736 776 4770
rect 810 4736 826 4770
rect 760 4702 826 4736
rect 760 4668 776 4702
rect 810 4668 826 4702
rect 760 4625 826 4668
rect 856 5382 922 5425
rect 856 5348 872 5382
rect 906 5348 922 5382
rect 856 5314 922 5348
rect 856 5280 872 5314
rect 906 5280 922 5314
rect 856 5246 922 5280
rect 856 5212 872 5246
rect 906 5212 922 5246
rect 856 5178 922 5212
rect 856 5144 872 5178
rect 906 5144 922 5178
rect 856 5110 922 5144
rect 856 5076 872 5110
rect 906 5076 922 5110
rect 856 5042 922 5076
rect 856 5008 872 5042
rect 906 5008 922 5042
rect 856 4974 922 5008
rect 856 4940 872 4974
rect 906 4940 922 4974
rect 856 4906 922 4940
rect 856 4872 872 4906
rect 906 4872 922 4906
rect 856 4838 922 4872
rect 856 4804 872 4838
rect 906 4804 922 4838
rect 856 4770 922 4804
rect 856 4736 872 4770
rect 906 4736 922 4770
rect 856 4702 922 4736
rect 856 4668 872 4702
rect 906 4668 922 4702
rect 856 4625 922 4668
rect 952 5382 1018 5425
rect 952 5348 968 5382
rect 1002 5348 1018 5382
rect 952 5314 1018 5348
rect 952 5280 968 5314
rect 1002 5280 1018 5314
rect 952 5246 1018 5280
rect 952 5212 968 5246
rect 1002 5212 1018 5246
rect 952 5178 1018 5212
rect 952 5144 968 5178
rect 1002 5144 1018 5178
rect 952 5110 1018 5144
rect 952 5076 968 5110
rect 1002 5076 1018 5110
rect 952 5042 1018 5076
rect 952 5008 968 5042
rect 1002 5008 1018 5042
rect 952 4974 1018 5008
rect 952 4940 968 4974
rect 1002 4940 1018 4974
rect 952 4906 1018 4940
rect 952 4872 968 4906
rect 1002 4872 1018 4906
rect 952 4838 1018 4872
rect 952 4804 968 4838
rect 1002 4804 1018 4838
rect 952 4770 1018 4804
rect 952 4736 968 4770
rect 1002 4736 1018 4770
rect 952 4702 1018 4736
rect 952 4668 968 4702
rect 1002 4668 1018 4702
rect 952 4625 1018 4668
rect 1048 5382 1114 5425
rect 1048 5348 1064 5382
rect 1098 5348 1114 5382
rect 1048 5314 1114 5348
rect 1048 5280 1064 5314
rect 1098 5280 1114 5314
rect 1048 5246 1114 5280
rect 1048 5212 1064 5246
rect 1098 5212 1114 5246
rect 1048 5178 1114 5212
rect 1048 5144 1064 5178
rect 1098 5144 1114 5178
rect 1048 5110 1114 5144
rect 1048 5076 1064 5110
rect 1098 5076 1114 5110
rect 1048 5042 1114 5076
rect 1048 5008 1064 5042
rect 1098 5008 1114 5042
rect 1048 4974 1114 5008
rect 1048 4940 1064 4974
rect 1098 4940 1114 4974
rect 1048 4906 1114 4940
rect 1048 4872 1064 4906
rect 1098 4872 1114 4906
rect 1048 4838 1114 4872
rect 1048 4804 1064 4838
rect 1098 4804 1114 4838
rect 1048 4770 1114 4804
rect 1048 4736 1064 4770
rect 1098 4736 1114 4770
rect 1048 4702 1114 4736
rect 1048 4668 1064 4702
rect 1098 4668 1114 4702
rect 1048 4625 1114 4668
rect 1144 5382 1210 5425
rect 1144 5348 1160 5382
rect 1194 5348 1210 5382
rect 1144 5314 1210 5348
rect 1144 5280 1160 5314
rect 1194 5280 1210 5314
rect 1144 5246 1210 5280
rect 1144 5212 1160 5246
rect 1194 5212 1210 5246
rect 1144 5178 1210 5212
rect 1144 5144 1160 5178
rect 1194 5144 1210 5178
rect 1144 5110 1210 5144
rect 1144 5076 1160 5110
rect 1194 5076 1210 5110
rect 1144 5042 1210 5076
rect 1144 5008 1160 5042
rect 1194 5008 1210 5042
rect 1144 4974 1210 5008
rect 1144 4940 1160 4974
rect 1194 4940 1210 4974
rect 1144 4906 1210 4940
rect 1144 4872 1160 4906
rect 1194 4872 1210 4906
rect 1144 4838 1210 4872
rect 1144 4804 1160 4838
rect 1194 4804 1210 4838
rect 1144 4770 1210 4804
rect 1144 4736 1160 4770
rect 1194 4736 1210 4770
rect 1144 4702 1210 4736
rect 1144 4668 1160 4702
rect 1194 4668 1210 4702
rect 1144 4625 1210 4668
rect 1240 5382 1306 5425
rect 1240 5348 1256 5382
rect 1290 5348 1306 5382
rect 1240 5314 1306 5348
rect 1240 5280 1256 5314
rect 1290 5280 1306 5314
rect 1240 5246 1306 5280
rect 1240 5212 1256 5246
rect 1290 5212 1306 5246
rect 1240 5178 1306 5212
rect 1240 5144 1256 5178
rect 1290 5144 1306 5178
rect 1240 5110 1306 5144
rect 1240 5076 1256 5110
rect 1290 5076 1306 5110
rect 1240 5042 1306 5076
rect 1240 5008 1256 5042
rect 1290 5008 1306 5042
rect 1240 4974 1306 5008
rect 1240 4940 1256 4974
rect 1290 4940 1306 4974
rect 1240 4906 1306 4940
rect 1240 4872 1256 4906
rect 1290 4872 1306 4906
rect 1240 4838 1306 4872
rect 1240 4804 1256 4838
rect 1290 4804 1306 4838
rect 1240 4770 1306 4804
rect 1240 4736 1256 4770
rect 1290 4736 1306 4770
rect 1240 4702 1306 4736
rect 1240 4668 1256 4702
rect 1290 4668 1306 4702
rect 1240 4625 1306 4668
rect 1336 5382 1402 5425
rect 1336 5348 1352 5382
rect 1386 5348 1402 5382
rect 1336 5314 1402 5348
rect 1336 5280 1352 5314
rect 1386 5280 1402 5314
rect 1336 5246 1402 5280
rect 1336 5212 1352 5246
rect 1386 5212 1402 5246
rect 1336 5178 1402 5212
rect 1336 5144 1352 5178
rect 1386 5144 1402 5178
rect 1336 5110 1402 5144
rect 1336 5076 1352 5110
rect 1386 5076 1402 5110
rect 1336 5042 1402 5076
rect 1336 5008 1352 5042
rect 1386 5008 1402 5042
rect 1336 4974 1402 5008
rect 1336 4940 1352 4974
rect 1386 4940 1402 4974
rect 1336 4906 1402 4940
rect 1336 4872 1352 4906
rect 1386 4872 1402 4906
rect 1336 4838 1402 4872
rect 1336 4804 1352 4838
rect 1386 4804 1402 4838
rect 1336 4770 1402 4804
rect 1336 4736 1352 4770
rect 1386 4736 1402 4770
rect 1336 4702 1402 4736
rect 1336 4668 1352 4702
rect 1386 4668 1402 4702
rect 1336 4625 1402 4668
rect 1432 5382 1498 5425
rect 1432 5348 1448 5382
rect 1482 5348 1498 5382
rect 1432 5314 1498 5348
rect 1432 5280 1448 5314
rect 1482 5280 1498 5314
rect 1432 5246 1498 5280
rect 1432 5212 1448 5246
rect 1482 5212 1498 5246
rect 1432 5178 1498 5212
rect 1432 5144 1448 5178
rect 1482 5144 1498 5178
rect 1432 5110 1498 5144
rect 1432 5076 1448 5110
rect 1482 5076 1498 5110
rect 1432 5042 1498 5076
rect 1432 5008 1448 5042
rect 1482 5008 1498 5042
rect 1432 4974 1498 5008
rect 1432 4940 1448 4974
rect 1482 4940 1498 4974
rect 1432 4906 1498 4940
rect 1432 4872 1448 4906
rect 1482 4872 1498 4906
rect 1432 4838 1498 4872
rect 1432 4804 1448 4838
rect 1482 4804 1498 4838
rect 1432 4770 1498 4804
rect 1432 4736 1448 4770
rect 1482 4736 1498 4770
rect 1432 4702 1498 4736
rect 1432 4668 1448 4702
rect 1482 4668 1498 4702
rect 1432 4625 1498 4668
rect 1528 5382 1594 5425
rect 1528 5348 1544 5382
rect 1578 5348 1594 5382
rect 1528 5314 1594 5348
rect 1528 5280 1544 5314
rect 1578 5280 1594 5314
rect 1528 5246 1594 5280
rect 1528 5212 1544 5246
rect 1578 5212 1594 5246
rect 1528 5178 1594 5212
rect 1528 5144 1544 5178
rect 1578 5144 1594 5178
rect 1528 5110 1594 5144
rect 1528 5076 1544 5110
rect 1578 5076 1594 5110
rect 1528 5042 1594 5076
rect 1528 5008 1544 5042
rect 1578 5008 1594 5042
rect 1528 4974 1594 5008
rect 1528 4940 1544 4974
rect 1578 4940 1594 4974
rect 1528 4906 1594 4940
rect 1528 4872 1544 4906
rect 1578 4872 1594 4906
rect 1528 4838 1594 4872
rect 1528 4804 1544 4838
rect 1578 4804 1594 4838
rect 1528 4770 1594 4804
rect 1528 4736 1544 4770
rect 1578 4736 1594 4770
rect 1528 4702 1594 4736
rect 1528 4668 1544 4702
rect 1578 4668 1594 4702
rect 1528 4625 1594 4668
rect 1624 5382 1690 5425
rect 1624 5348 1640 5382
rect 1674 5348 1690 5382
rect 1624 5314 1690 5348
rect 1624 5280 1640 5314
rect 1674 5280 1690 5314
rect 1624 5246 1690 5280
rect 1624 5212 1640 5246
rect 1674 5212 1690 5246
rect 1624 5178 1690 5212
rect 1624 5144 1640 5178
rect 1674 5144 1690 5178
rect 1624 5110 1690 5144
rect 1624 5076 1640 5110
rect 1674 5076 1690 5110
rect 1624 5042 1690 5076
rect 1624 5008 1640 5042
rect 1674 5008 1690 5042
rect 1624 4974 1690 5008
rect 1624 4940 1640 4974
rect 1674 4940 1690 4974
rect 1624 4906 1690 4940
rect 1624 4872 1640 4906
rect 1674 4872 1690 4906
rect 1624 4838 1690 4872
rect 1624 4804 1640 4838
rect 1674 4804 1690 4838
rect 1624 4770 1690 4804
rect 1624 4736 1640 4770
rect 1674 4736 1690 4770
rect 1624 4702 1690 4736
rect 1624 4668 1640 4702
rect 1674 4668 1690 4702
rect 1624 4625 1690 4668
rect 1720 5382 1786 5425
rect 1720 5348 1736 5382
rect 1770 5348 1786 5382
rect 1720 5314 1786 5348
rect 1720 5280 1736 5314
rect 1770 5280 1786 5314
rect 1720 5246 1786 5280
rect 1720 5212 1736 5246
rect 1770 5212 1786 5246
rect 1720 5178 1786 5212
rect 1720 5144 1736 5178
rect 1770 5144 1786 5178
rect 1720 5110 1786 5144
rect 1720 5076 1736 5110
rect 1770 5076 1786 5110
rect 1720 5042 1786 5076
rect 1720 5008 1736 5042
rect 1770 5008 1786 5042
rect 1720 4974 1786 5008
rect 1720 4940 1736 4974
rect 1770 4940 1786 4974
rect 1720 4906 1786 4940
rect 1720 4872 1736 4906
rect 1770 4872 1786 4906
rect 1720 4838 1786 4872
rect 1720 4804 1736 4838
rect 1770 4804 1786 4838
rect 1720 4770 1786 4804
rect 1720 4736 1736 4770
rect 1770 4736 1786 4770
rect 1720 4702 1786 4736
rect 1720 4668 1736 4702
rect 1770 4668 1786 4702
rect 1720 4625 1786 4668
rect 1816 5382 1882 5425
rect 1816 5348 1832 5382
rect 1866 5348 1882 5382
rect 1816 5314 1882 5348
rect 1816 5280 1832 5314
rect 1866 5280 1882 5314
rect 1816 5246 1882 5280
rect 1816 5212 1832 5246
rect 1866 5212 1882 5246
rect 1816 5178 1882 5212
rect 1816 5144 1832 5178
rect 1866 5144 1882 5178
rect 1816 5110 1882 5144
rect 1816 5076 1832 5110
rect 1866 5076 1882 5110
rect 1816 5042 1882 5076
rect 1816 5008 1832 5042
rect 1866 5008 1882 5042
rect 1816 4974 1882 5008
rect 1816 4940 1832 4974
rect 1866 4940 1882 4974
rect 1816 4906 1882 4940
rect 1816 4872 1832 4906
rect 1866 4872 1882 4906
rect 1816 4838 1882 4872
rect 1816 4804 1832 4838
rect 1866 4804 1882 4838
rect 1816 4770 1882 4804
rect 1816 4736 1832 4770
rect 1866 4736 1882 4770
rect 1816 4702 1882 4736
rect 1816 4668 1832 4702
rect 1866 4668 1882 4702
rect 1816 4625 1882 4668
rect 1912 5382 1974 5425
rect 1912 5348 1928 5382
rect 1962 5348 1974 5382
rect 1912 5314 1974 5348
rect 1912 5280 1928 5314
rect 1962 5280 1974 5314
rect 1912 5246 1974 5280
rect 1912 5212 1928 5246
rect 1962 5212 1974 5246
rect 1912 5178 1974 5212
rect 1912 5144 1928 5178
rect 1962 5144 1974 5178
rect 1912 5110 1974 5144
rect 1912 5076 1928 5110
rect 1962 5076 1974 5110
rect 1912 5042 1974 5076
rect 1912 5008 1928 5042
rect 1962 5008 1974 5042
rect 1912 4974 1974 5008
rect 1912 4940 1928 4974
rect 1962 4940 1974 4974
rect 1912 4906 1974 4940
rect 1912 4872 1928 4906
rect 1962 4872 1974 4906
rect 1912 4838 1974 4872
rect 1912 4804 1928 4838
rect 1962 4804 1974 4838
rect 1912 4770 1974 4804
rect 1912 4736 1928 4770
rect 1962 4736 1974 4770
rect 1912 4702 1974 4736
rect 1912 4668 1928 4702
rect 1962 4668 1974 4702
rect 1912 4625 1974 4668
rect -42537 -4780 -42475 -4737
rect -42537 -4814 -42525 -4780
rect -42491 -4814 -42475 -4780
rect -42537 -4848 -42475 -4814
rect -42537 -4882 -42525 -4848
rect -42491 -4882 -42475 -4848
rect -42537 -4916 -42475 -4882
rect -42537 -4950 -42525 -4916
rect -42491 -4950 -42475 -4916
rect -42537 -4984 -42475 -4950
rect -42537 -5018 -42525 -4984
rect -42491 -5018 -42475 -4984
rect -42537 -5052 -42475 -5018
rect -42537 -5086 -42525 -5052
rect -42491 -5086 -42475 -5052
rect -42537 -5120 -42475 -5086
rect -42537 -5154 -42525 -5120
rect -42491 -5154 -42475 -5120
rect -42537 -5188 -42475 -5154
rect -42537 -5222 -42525 -5188
rect -42491 -5222 -42475 -5188
rect -42537 -5256 -42475 -5222
rect -42537 -5290 -42525 -5256
rect -42491 -5290 -42475 -5256
rect -42537 -5324 -42475 -5290
rect -42537 -5358 -42525 -5324
rect -42491 -5358 -42475 -5324
rect -42537 -5392 -42475 -5358
rect -42537 -5426 -42525 -5392
rect -42491 -5426 -42475 -5392
rect -42537 -5460 -42475 -5426
rect -42537 -5494 -42525 -5460
rect -42491 -5494 -42475 -5460
rect -42537 -5537 -42475 -5494
rect -42445 -4780 -42379 -4737
rect -42445 -4814 -42429 -4780
rect -42395 -4814 -42379 -4780
rect -42445 -4848 -42379 -4814
rect -42445 -4882 -42429 -4848
rect -42395 -4882 -42379 -4848
rect -42445 -4916 -42379 -4882
rect -42445 -4950 -42429 -4916
rect -42395 -4950 -42379 -4916
rect -42445 -4984 -42379 -4950
rect -42445 -5018 -42429 -4984
rect -42395 -5018 -42379 -4984
rect -42445 -5052 -42379 -5018
rect -42445 -5086 -42429 -5052
rect -42395 -5086 -42379 -5052
rect -42445 -5120 -42379 -5086
rect -42445 -5154 -42429 -5120
rect -42395 -5154 -42379 -5120
rect -42445 -5188 -42379 -5154
rect -42445 -5222 -42429 -5188
rect -42395 -5222 -42379 -5188
rect -42445 -5256 -42379 -5222
rect -42445 -5290 -42429 -5256
rect -42395 -5290 -42379 -5256
rect -42445 -5324 -42379 -5290
rect -42445 -5358 -42429 -5324
rect -42395 -5358 -42379 -5324
rect -42445 -5392 -42379 -5358
rect -42445 -5426 -42429 -5392
rect -42395 -5426 -42379 -5392
rect -42445 -5460 -42379 -5426
rect -42445 -5494 -42429 -5460
rect -42395 -5494 -42379 -5460
rect -42445 -5537 -42379 -5494
rect -42349 -4780 -42283 -4737
rect -42349 -4814 -42333 -4780
rect -42299 -4814 -42283 -4780
rect -42349 -4848 -42283 -4814
rect -42349 -4882 -42333 -4848
rect -42299 -4882 -42283 -4848
rect -42349 -4916 -42283 -4882
rect -42349 -4950 -42333 -4916
rect -42299 -4950 -42283 -4916
rect -42349 -4984 -42283 -4950
rect -42349 -5018 -42333 -4984
rect -42299 -5018 -42283 -4984
rect -42349 -5052 -42283 -5018
rect -42349 -5086 -42333 -5052
rect -42299 -5086 -42283 -5052
rect -42349 -5120 -42283 -5086
rect -42349 -5154 -42333 -5120
rect -42299 -5154 -42283 -5120
rect -42349 -5188 -42283 -5154
rect -42349 -5222 -42333 -5188
rect -42299 -5222 -42283 -5188
rect -42349 -5256 -42283 -5222
rect -42349 -5290 -42333 -5256
rect -42299 -5290 -42283 -5256
rect -42349 -5324 -42283 -5290
rect -42349 -5358 -42333 -5324
rect -42299 -5358 -42283 -5324
rect -42349 -5392 -42283 -5358
rect -42349 -5426 -42333 -5392
rect -42299 -5426 -42283 -5392
rect -42349 -5460 -42283 -5426
rect -42349 -5494 -42333 -5460
rect -42299 -5494 -42283 -5460
rect -42349 -5537 -42283 -5494
rect -42253 -4780 -42187 -4737
rect -42253 -4814 -42237 -4780
rect -42203 -4814 -42187 -4780
rect -42253 -4848 -42187 -4814
rect -42253 -4882 -42237 -4848
rect -42203 -4882 -42187 -4848
rect -42253 -4916 -42187 -4882
rect -42253 -4950 -42237 -4916
rect -42203 -4950 -42187 -4916
rect -42253 -4984 -42187 -4950
rect -42253 -5018 -42237 -4984
rect -42203 -5018 -42187 -4984
rect -42253 -5052 -42187 -5018
rect -42253 -5086 -42237 -5052
rect -42203 -5086 -42187 -5052
rect -42253 -5120 -42187 -5086
rect -42253 -5154 -42237 -5120
rect -42203 -5154 -42187 -5120
rect -42253 -5188 -42187 -5154
rect -42253 -5222 -42237 -5188
rect -42203 -5222 -42187 -5188
rect -42253 -5256 -42187 -5222
rect -42253 -5290 -42237 -5256
rect -42203 -5290 -42187 -5256
rect -42253 -5324 -42187 -5290
rect -42253 -5358 -42237 -5324
rect -42203 -5358 -42187 -5324
rect -42253 -5392 -42187 -5358
rect -42253 -5426 -42237 -5392
rect -42203 -5426 -42187 -5392
rect -42253 -5460 -42187 -5426
rect -42253 -5494 -42237 -5460
rect -42203 -5494 -42187 -5460
rect -42253 -5537 -42187 -5494
rect -42157 -4780 -42091 -4737
rect -42157 -4814 -42141 -4780
rect -42107 -4814 -42091 -4780
rect -42157 -4848 -42091 -4814
rect -42157 -4882 -42141 -4848
rect -42107 -4882 -42091 -4848
rect -42157 -4916 -42091 -4882
rect -42157 -4950 -42141 -4916
rect -42107 -4950 -42091 -4916
rect -42157 -4984 -42091 -4950
rect -42157 -5018 -42141 -4984
rect -42107 -5018 -42091 -4984
rect -42157 -5052 -42091 -5018
rect -42157 -5086 -42141 -5052
rect -42107 -5086 -42091 -5052
rect -42157 -5120 -42091 -5086
rect -42157 -5154 -42141 -5120
rect -42107 -5154 -42091 -5120
rect -42157 -5188 -42091 -5154
rect -42157 -5222 -42141 -5188
rect -42107 -5222 -42091 -5188
rect -42157 -5256 -42091 -5222
rect -42157 -5290 -42141 -5256
rect -42107 -5290 -42091 -5256
rect -42157 -5324 -42091 -5290
rect -42157 -5358 -42141 -5324
rect -42107 -5358 -42091 -5324
rect -42157 -5392 -42091 -5358
rect -42157 -5426 -42141 -5392
rect -42107 -5426 -42091 -5392
rect -42157 -5460 -42091 -5426
rect -42157 -5494 -42141 -5460
rect -42107 -5494 -42091 -5460
rect -42157 -5537 -42091 -5494
rect -42061 -4780 -41995 -4737
rect -42061 -4814 -42045 -4780
rect -42011 -4814 -41995 -4780
rect -42061 -4848 -41995 -4814
rect -42061 -4882 -42045 -4848
rect -42011 -4882 -41995 -4848
rect -42061 -4916 -41995 -4882
rect -42061 -4950 -42045 -4916
rect -42011 -4950 -41995 -4916
rect -42061 -4984 -41995 -4950
rect -42061 -5018 -42045 -4984
rect -42011 -5018 -41995 -4984
rect -42061 -5052 -41995 -5018
rect -42061 -5086 -42045 -5052
rect -42011 -5086 -41995 -5052
rect -42061 -5120 -41995 -5086
rect -42061 -5154 -42045 -5120
rect -42011 -5154 -41995 -5120
rect -42061 -5188 -41995 -5154
rect -42061 -5222 -42045 -5188
rect -42011 -5222 -41995 -5188
rect -42061 -5256 -41995 -5222
rect -42061 -5290 -42045 -5256
rect -42011 -5290 -41995 -5256
rect -42061 -5324 -41995 -5290
rect -42061 -5358 -42045 -5324
rect -42011 -5358 -41995 -5324
rect -42061 -5392 -41995 -5358
rect -42061 -5426 -42045 -5392
rect -42011 -5426 -41995 -5392
rect -42061 -5460 -41995 -5426
rect -42061 -5494 -42045 -5460
rect -42011 -5494 -41995 -5460
rect -42061 -5537 -41995 -5494
rect -41965 -4780 -41899 -4737
rect -41965 -4814 -41949 -4780
rect -41915 -4814 -41899 -4780
rect -41965 -4848 -41899 -4814
rect -41965 -4882 -41949 -4848
rect -41915 -4882 -41899 -4848
rect -41965 -4916 -41899 -4882
rect -41965 -4950 -41949 -4916
rect -41915 -4950 -41899 -4916
rect -41965 -4984 -41899 -4950
rect -41965 -5018 -41949 -4984
rect -41915 -5018 -41899 -4984
rect -41965 -5052 -41899 -5018
rect -41965 -5086 -41949 -5052
rect -41915 -5086 -41899 -5052
rect -41965 -5120 -41899 -5086
rect -41965 -5154 -41949 -5120
rect -41915 -5154 -41899 -5120
rect -41965 -5188 -41899 -5154
rect -41965 -5222 -41949 -5188
rect -41915 -5222 -41899 -5188
rect -41965 -5256 -41899 -5222
rect -41965 -5290 -41949 -5256
rect -41915 -5290 -41899 -5256
rect -41965 -5324 -41899 -5290
rect -41965 -5358 -41949 -5324
rect -41915 -5358 -41899 -5324
rect -41965 -5392 -41899 -5358
rect -41965 -5426 -41949 -5392
rect -41915 -5426 -41899 -5392
rect -41965 -5460 -41899 -5426
rect -41965 -5494 -41949 -5460
rect -41915 -5494 -41899 -5460
rect -41965 -5537 -41899 -5494
rect -41869 -4780 -41803 -4737
rect -41869 -4814 -41853 -4780
rect -41819 -4814 -41803 -4780
rect -41869 -4848 -41803 -4814
rect -41869 -4882 -41853 -4848
rect -41819 -4882 -41803 -4848
rect -41869 -4916 -41803 -4882
rect -41869 -4950 -41853 -4916
rect -41819 -4950 -41803 -4916
rect -41869 -4984 -41803 -4950
rect -41869 -5018 -41853 -4984
rect -41819 -5018 -41803 -4984
rect -41869 -5052 -41803 -5018
rect -41869 -5086 -41853 -5052
rect -41819 -5086 -41803 -5052
rect -41869 -5120 -41803 -5086
rect -41869 -5154 -41853 -5120
rect -41819 -5154 -41803 -5120
rect -41869 -5188 -41803 -5154
rect -41869 -5222 -41853 -5188
rect -41819 -5222 -41803 -5188
rect -41869 -5256 -41803 -5222
rect -41869 -5290 -41853 -5256
rect -41819 -5290 -41803 -5256
rect -41869 -5324 -41803 -5290
rect -41869 -5358 -41853 -5324
rect -41819 -5358 -41803 -5324
rect -41869 -5392 -41803 -5358
rect -41869 -5426 -41853 -5392
rect -41819 -5426 -41803 -5392
rect -41869 -5460 -41803 -5426
rect -41869 -5494 -41853 -5460
rect -41819 -5494 -41803 -5460
rect -41869 -5537 -41803 -5494
rect -41773 -4780 -41707 -4737
rect -41773 -4814 -41757 -4780
rect -41723 -4814 -41707 -4780
rect -41773 -4848 -41707 -4814
rect -41773 -4882 -41757 -4848
rect -41723 -4882 -41707 -4848
rect -41773 -4916 -41707 -4882
rect -41773 -4950 -41757 -4916
rect -41723 -4950 -41707 -4916
rect -41773 -4984 -41707 -4950
rect -41773 -5018 -41757 -4984
rect -41723 -5018 -41707 -4984
rect -41773 -5052 -41707 -5018
rect -41773 -5086 -41757 -5052
rect -41723 -5086 -41707 -5052
rect -41773 -5120 -41707 -5086
rect -41773 -5154 -41757 -5120
rect -41723 -5154 -41707 -5120
rect -41773 -5188 -41707 -5154
rect -41773 -5222 -41757 -5188
rect -41723 -5222 -41707 -5188
rect -41773 -5256 -41707 -5222
rect -41773 -5290 -41757 -5256
rect -41723 -5290 -41707 -5256
rect -41773 -5324 -41707 -5290
rect -41773 -5358 -41757 -5324
rect -41723 -5358 -41707 -5324
rect -41773 -5392 -41707 -5358
rect -41773 -5426 -41757 -5392
rect -41723 -5426 -41707 -5392
rect -41773 -5460 -41707 -5426
rect -41773 -5494 -41757 -5460
rect -41723 -5494 -41707 -5460
rect -41773 -5537 -41707 -5494
rect -41677 -4780 -41611 -4737
rect -41677 -4814 -41661 -4780
rect -41627 -4814 -41611 -4780
rect -41677 -4848 -41611 -4814
rect -41677 -4882 -41661 -4848
rect -41627 -4882 -41611 -4848
rect -41677 -4916 -41611 -4882
rect -41677 -4950 -41661 -4916
rect -41627 -4950 -41611 -4916
rect -41677 -4984 -41611 -4950
rect -41677 -5018 -41661 -4984
rect -41627 -5018 -41611 -4984
rect -41677 -5052 -41611 -5018
rect -41677 -5086 -41661 -5052
rect -41627 -5086 -41611 -5052
rect -41677 -5120 -41611 -5086
rect -41677 -5154 -41661 -5120
rect -41627 -5154 -41611 -5120
rect -41677 -5188 -41611 -5154
rect -41677 -5222 -41661 -5188
rect -41627 -5222 -41611 -5188
rect -41677 -5256 -41611 -5222
rect -41677 -5290 -41661 -5256
rect -41627 -5290 -41611 -5256
rect -41677 -5324 -41611 -5290
rect -41677 -5358 -41661 -5324
rect -41627 -5358 -41611 -5324
rect -41677 -5392 -41611 -5358
rect -41677 -5426 -41661 -5392
rect -41627 -5426 -41611 -5392
rect -41677 -5460 -41611 -5426
rect -41677 -5494 -41661 -5460
rect -41627 -5494 -41611 -5460
rect -41677 -5537 -41611 -5494
rect -41581 -4780 -41515 -4737
rect -41581 -4814 -41565 -4780
rect -41531 -4814 -41515 -4780
rect -41581 -4848 -41515 -4814
rect -41581 -4882 -41565 -4848
rect -41531 -4882 -41515 -4848
rect -41581 -4916 -41515 -4882
rect -41581 -4950 -41565 -4916
rect -41531 -4950 -41515 -4916
rect -41581 -4984 -41515 -4950
rect -41581 -5018 -41565 -4984
rect -41531 -5018 -41515 -4984
rect -41581 -5052 -41515 -5018
rect -41581 -5086 -41565 -5052
rect -41531 -5086 -41515 -5052
rect -41581 -5120 -41515 -5086
rect -41581 -5154 -41565 -5120
rect -41531 -5154 -41515 -5120
rect -41581 -5188 -41515 -5154
rect -41581 -5222 -41565 -5188
rect -41531 -5222 -41515 -5188
rect -41581 -5256 -41515 -5222
rect -41581 -5290 -41565 -5256
rect -41531 -5290 -41515 -5256
rect -41581 -5324 -41515 -5290
rect -41581 -5358 -41565 -5324
rect -41531 -5358 -41515 -5324
rect -41581 -5392 -41515 -5358
rect -41581 -5426 -41565 -5392
rect -41531 -5426 -41515 -5392
rect -41581 -5460 -41515 -5426
rect -41581 -5494 -41565 -5460
rect -41531 -5494 -41515 -5460
rect -41581 -5537 -41515 -5494
rect -41485 -4780 -41419 -4737
rect -41485 -4814 -41469 -4780
rect -41435 -4814 -41419 -4780
rect -41485 -4848 -41419 -4814
rect -41485 -4882 -41469 -4848
rect -41435 -4882 -41419 -4848
rect -41485 -4916 -41419 -4882
rect -41485 -4950 -41469 -4916
rect -41435 -4950 -41419 -4916
rect -41485 -4984 -41419 -4950
rect -41485 -5018 -41469 -4984
rect -41435 -5018 -41419 -4984
rect -41485 -5052 -41419 -5018
rect -41485 -5086 -41469 -5052
rect -41435 -5086 -41419 -5052
rect -41485 -5120 -41419 -5086
rect -41485 -5154 -41469 -5120
rect -41435 -5154 -41419 -5120
rect -41485 -5188 -41419 -5154
rect -41485 -5222 -41469 -5188
rect -41435 -5222 -41419 -5188
rect -41485 -5256 -41419 -5222
rect -41485 -5290 -41469 -5256
rect -41435 -5290 -41419 -5256
rect -41485 -5324 -41419 -5290
rect -41485 -5358 -41469 -5324
rect -41435 -5358 -41419 -5324
rect -41485 -5392 -41419 -5358
rect -41485 -5426 -41469 -5392
rect -41435 -5426 -41419 -5392
rect -41485 -5460 -41419 -5426
rect -41485 -5494 -41469 -5460
rect -41435 -5494 -41419 -5460
rect -41485 -5537 -41419 -5494
rect -41389 -4780 -41323 -4737
rect -41389 -4814 -41373 -4780
rect -41339 -4814 -41323 -4780
rect -41389 -4848 -41323 -4814
rect -41389 -4882 -41373 -4848
rect -41339 -4882 -41323 -4848
rect -41389 -4916 -41323 -4882
rect -41389 -4950 -41373 -4916
rect -41339 -4950 -41323 -4916
rect -41389 -4984 -41323 -4950
rect -41389 -5018 -41373 -4984
rect -41339 -5018 -41323 -4984
rect -41389 -5052 -41323 -5018
rect -41389 -5086 -41373 -5052
rect -41339 -5086 -41323 -5052
rect -41389 -5120 -41323 -5086
rect -41389 -5154 -41373 -5120
rect -41339 -5154 -41323 -5120
rect -41389 -5188 -41323 -5154
rect -41389 -5222 -41373 -5188
rect -41339 -5222 -41323 -5188
rect -41389 -5256 -41323 -5222
rect -41389 -5290 -41373 -5256
rect -41339 -5290 -41323 -5256
rect -41389 -5324 -41323 -5290
rect -41389 -5358 -41373 -5324
rect -41339 -5358 -41323 -5324
rect -41389 -5392 -41323 -5358
rect -41389 -5426 -41373 -5392
rect -41339 -5426 -41323 -5392
rect -41389 -5460 -41323 -5426
rect -41389 -5494 -41373 -5460
rect -41339 -5494 -41323 -5460
rect -41389 -5537 -41323 -5494
rect -41293 -4780 -41227 -4737
rect -41293 -4814 -41277 -4780
rect -41243 -4814 -41227 -4780
rect -41293 -4848 -41227 -4814
rect -41293 -4882 -41277 -4848
rect -41243 -4882 -41227 -4848
rect -41293 -4916 -41227 -4882
rect -41293 -4950 -41277 -4916
rect -41243 -4950 -41227 -4916
rect -41293 -4984 -41227 -4950
rect -41293 -5018 -41277 -4984
rect -41243 -5018 -41227 -4984
rect -41293 -5052 -41227 -5018
rect -41293 -5086 -41277 -5052
rect -41243 -5086 -41227 -5052
rect -41293 -5120 -41227 -5086
rect -41293 -5154 -41277 -5120
rect -41243 -5154 -41227 -5120
rect -41293 -5188 -41227 -5154
rect -41293 -5222 -41277 -5188
rect -41243 -5222 -41227 -5188
rect -41293 -5256 -41227 -5222
rect -41293 -5290 -41277 -5256
rect -41243 -5290 -41227 -5256
rect -41293 -5324 -41227 -5290
rect -41293 -5358 -41277 -5324
rect -41243 -5358 -41227 -5324
rect -41293 -5392 -41227 -5358
rect -41293 -5426 -41277 -5392
rect -41243 -5426 -41227 -5392
rect -41293 -5460 -41227 -5426
rect -41293 -5494 -41277 -5460
rect -41243 -5494 -41227 -5460
rect -41293 -5537 -41227 -5494
rect -41197 -4780 -41131 -4737
rect -41197 -4814 -41181 -4780
rect -41147 -4814 -41131 -4780
rect -41197 -4848 -41131 -4814
rect -41197 -4882 -41181 -4848
rect -41147 -4882 -41131 -4848
rect -41197 -4916 -41131 -4882
rect -41197 -4950 -41181 -4916
rect -41147 -4950 -41131 -4916
rect -41197 -4984 -41131 -4950
rect -41197 -5018 -41181 -4984
rect -41147 -5018 -41131 -4984
rect -41197 -5052 -41131 -5018
rect -41197 -5086 -41181 -5052
rect -41147 -5086 -41131 -5052
rect -41197 -5120 -41131 -5086
rect -41197 -5154 -41181 -5120
rect -41147 -5154 -41131 -5120
rect -41197 -5188 -41131 -5154
rect -41197 -5222 -41181 -5188
rect -41147 -5222 -41131 -5188
rect -41197 -5256 -41131 -5222
rect -41197 -5290 -41181 -5256
rect -41147 -5290 -41131 -5256
rect -41197 -5324 -41131 -5290
rect -41197 -5358 -41181 -5324
rect -41147 -5358 -41131 -5324
rect -41197 -5392 -41131 -5358
rect -41197 -5426 -41181 -5392
rect -41147 -5426 -41131 -5392
rect -41197 -5460 -41131 -5426
rect -41197 -5494 -41181 -5460
rect -41147 -5494 -41131 -5460
rect -41197 -5537 -41131 -5494
rect -41101 -4780 -41035 -4737
rect -41101 -4814 -41085 -4780
rect -41051 -4814 -41035 -4780
rect -41101 -4848 -41035 -4814
rect -41101 -4882 -41085 -4848
rect -41051 -4882 -41035 -4848
rect -41101 -4916 -41035 -4882
rect -41101 -4950 -41085 -4916
rect -41051 -4950 -41035 -4916
rect -41101 -4984 -41035 -4950
rect -41101 -5018 -41085 -4984
rect -41051 -5018 -41035 -4984
rect -41101 -5052 -41035 -5018
rect -41101 -5086 -41085 -5052
rect -41051 -5086 -41035 -5052
rect -41101 -5120 -41035 -5086
rect -41101 -5154 -41085 -5120
rect -41051 -5154 -41035 -5120
rect -41101 -5188 -41035 -5154
rect -41101 -5222 -41085 -5188
rect -41051 -5222 -41035 -5188
rect -41101 -5256 -41035 -5222
rect -41101 -5290 -41085 -5256
rect -41051 -5290 -41035 -5256
rect -41101 -5324 -41035 -5290
rect -41101 -5358 -41085 -5324
rect -41051 -5358 -41035 -5324
rect -41101 -5392 -41035 -5358
rect -41101 -5426 -41085 -5392
rect -41051 -5426 -41035 -5392
rect -41101 -5460 -41035 -5426
rect -41101 -5494 -41085 -5460
rect -41051 -5494 -41035 -5460
rect -41101 -5537 -41035 -5494
rect -41005 -4780 -40939 -4737
rect -41005 -4814 -40989 -4780
rect -40955 -4814 -40939 -4780
rect -41005 -4848 -40939 -4814
rect -41005 -4882 -40989 -4848
rect -40955 -4882 -40939 -4848
rect -41005 -4916 -40939 -4882
rect -41005 -4950 -40989 -4916
rect -40955 -4950 -40939 -4916
rect -41005 -4984 -40939 -4950
rect -41005 -5018 -40989 -4984
rect -40955 -5018 -40939 -4984
rect -41005 -5052 -40939 -5018
rect -41005 -5086 -40989 -5052
rect -40955 -5086 -40939 -5052
rect -41005 -5120 -40939 -5086
rect -41005 -5154 -40989 -5120
rect -40955 -5154 -40939 -5120
rect -41005 -5188 -40939 -5154
rect -41005 -5222 -40989 -5188
rect -40955 -5222 -40939 -5188
rect -41005 -5256 -40939 -5222
rect -41005 -5290 -40989 -5256
rect -40955 -5290 -40939 -5256
rect -41005 -5324 -40939 -5290
rect -41005 -5358 -40989 -5324
rect -40955 -5358 -40939 -5324
rect -41005 -5392 -40939 -5358
rect -41005 -5426 -40989 -5392
rect -40955 -5426 -40939 -5392
rect -41005 -5460 -40939 -5426
rect -41005 -5494 -40989 -5460
rect -40955 -5494 -40939 -5460
rect -41005 -5537 -40939 -5494
rect -40909 -4780 -40843 -4737
rect -40909 -4814 -40893 -4780
rect -40859 -4814 -40843 -4780
rect -40909 -4848 -40843 -4814
rect -40909 -4882 -40893 -4848
rect -40859 -4882 -40843 -4848
rect -40909 -4916 -40843 -4882
rect -40909 -4950 -40893 -4916
rect -40859 -4950 -40843 -4916
rect -40909 -4984 -40843 -4950
rect -40909 -5018 -40893 -4984
rect -40859 -5018 -40843 -4984
rect -40909 -5052 -40843 -5018
rect -40909 -5086 -40893 -5052
rect -40859 -5086 -40843 -5052
rect -40909 -5120 -40843 -5086
rect -40909 -5154 -40893 -5120
rect -40859 -5154 -40843 -5120
rect -40909 -5188 -40843 -5154
rect -40909 -5222 -40893 -5188
rect -40859 -5222 -40843 -5188
rect -40909 -5256 -40843 -5222
rect -40909 -5290 -40893 -5256
rect -40859 -5290 -40843 -5256
rect -40909 -5324 -40843 -5290
rect -40909 -5358 -40893 -5324
rect -40859 -5358 -40843 -5324
rect -40909 -5392 -40843 -5358
rect -40909 -5426 -40893 -5392
rect -40859 -5426 -40843 -5392
rect -40909 -5460 -40843 -5426
rect -40909 -5494 -40893 -5460
rect -40859 -5494 -40843 -5460
rect -40909 -5537 -40843 -5494
rect -40813 -4780 -40747 -4737
rect -40813 -4814 -40797 -4780
rect -40763 -4814 -40747 -4780
rect -40813 -4848 -40747 -4814
rect -40813 -4882 -40797 -4848
rect -40763 -4882 -40747 -4848
rect -40813 -4916 -40747 -4882
rect -40813 -4950 -40797 -4916
rect -40763 -4950 -40747 -4916
rect -40813 -4984 -40747 -4950
rect -40813 -5018 -40797 -4984
rect -40763 -5018 -40747 -4984
rect -40813 -5052 -40747 -5018
rect -40813 -5086 -40797 -5052
rect -40763 -5086 -40747 -5052
rect -40813 -5120 -40747 -5086
rect -40813 -5154 -40797 -5120
rect -40763 -5154 -40747 -5120
rect -40813 -5188 -40747 -5154
rect -40813 -5222 -40797 -5188
rect -40763 -5222 -40747 -5188
rect -40813 -5256 -40747 -5222
rect -40813 -5290 -40797 -5256
rect -40763 -5290 -40747 -5256
rect -40813 -5324 -40747 -5290
rect -40813 -5358 -40797 -5324
rect -40763 -5358 -40747 -5324
rect -40813 -5392 -40747 -5358
rect -40813 -5426 -40797 -5392
rect -40763 -5426 -40747 -5392
rect -40813 -5460 -40747 -5426
rect -40813 -5494 -40797 -5460
rect -40763 -5494 -40747 -5460
rect -40813 -5537 -40747 -5494
rect -40717 -4780 -40655 -4737
rect -40717 -4814 -40701 -4780
rect -40667 -4814 -40655 -4780
rect -40717 -4848 -40655 -4814
rect -40717 -4882 -40701 -4848
rect -40667 -4882 -40655 -4848
rect -40717 -4916 -40655 -4882
rect -40717 -4950 -40701 -4916
rect -40667 -4950 -40655 -4916
rect -40717 -4984 -40655 -4950
rect -40717 -5018 -40701 -4984
rect -40667 -5018 -40655 -4984
rect -40717 -5052 -40655 -5018
rect -40717 -5086 -40701 -5052
rect -40667 -5086 -40655 -5052
rect -40717 -5120 -40655 -5086
rect -40717 -5154 -40701 -5120
rect -40667 -5154 -40655 -5120
rect -40717 -5188 -40655 -5154
rect -40717 -5222 -40701 -5188
rect -40667 -5222 -40655 -5188
rect -40717 -5256 -40655 -5222
rect -40717 -5290 -40701 -5256
rect -40667 -5290 -40655 -5256
rect -40717 -5324 -40655 -5290
rect -40717 -5358 -40701 -5324
rect -40667 -5358 -40655 -5324
rect -40717 -5392 -40655 -5358
rect -40717 -5426 -40701 -5392
rect -40667 -5426 -40655 -5392
rect -40717 -5460 -40655 -5426
rect -40717 -5494 -40701 -5460
rect -40667 -5494 -40655 -5460
rect -40717 -5537 -40655 -5494
rect 104 -4806 166 -4763
rect 104 -4840 116 -4806
rect 150 -4840 166 -4806
rect 104 -4874 166 -4840
rect 104 -4908 116 -4874
rect 150 -4908 166 -4874
rect 104 -4942 166 -4908
rect 104 -4976 116 -4942
rect 150 -4976 166 -4942
rect 104 -5010 166 -4976
rect 104 -5044 116 -5010
rect 150 -5044 166 -5010
rect 104 -5078 166 -5044
rect 104 -5112 116 -5078
rect 150 -5112 166 -5078
rect 104 -5146 166 -5112
rect 104 -5180 116 -5146
rect 150 -5180 166 -5146
rect 104 -5214 166 -5180
rect 104 -5248 116 -5214
rect 150 -5248 166 -5214
rect 104 -5282 166 -5248
rect 104 -5316 116 -5282
rect 150 -5316 166 -5282
rect 104 -5350 166 -5316
rect 104 -5384 116 -5350
rect 150 -5384 166 -5350
rect 104 -5418 166 -5384
rect 104 -5452 116 -5418
rect 150 -5452 166 -5418
rect 104 -5486 166 -5452
rect 104 -5520 116 -5486
rect 150 -5520 166 -5486
rect 104 -5563 166 -5520
rect 196 -4806 262 -4763
rect 196 -4840 212 -4806
rect 246 -4840 262 -4806
rect 196 -4874 262 -4840
rect 196 -4908 212 -4874
rect 246 -4908 262 -4874
rect 196 -4942 262 -4908
rect 196 -4976 212 -4942
rect 246 -4976 262 -4942
rect 196 -5010 262 -4976
rect 196 -5044 212 -5010
rect 246 -5044 262 -5010
rect 196 -5078 262 -5044
rect 196 -5112 212 -5078
rect 246 -5112 262 -5078
rect 196 -5146 262 -5112
rect 196 -5180 212 -5146
rect 246 -5180 262 -5146
rect 196 -5214 262 -5180
rect 196 -5248 212 -5214
rect 246 -5248 262 -5214
rect 196 -5282 262 -5248
rect 196 -5316 212 -5282
rect 246 -5316 262 -5282
rect 196 -5350 262 -5316
rect 196 -5384 212 -5350
rect 246 -5384 262 -5350
rect 196 -5418 262 -5384
rect 196 -5452 212 -5418
rect 246 -5452 262 -5418
rect 196 -5486 262 -5452
rect 196 -5520 212 -5486
rect 246 -5520 262 -5486
rect 196 -5563 262 -5520
rect 292 -4806 358 -4763
rect 292 -4840 308 -4806
rect 342 -4840 358 -4806
rect 292 -4874 358 -4840
rect 292 -4908 308 -4874
rect 342 -4908 358 -4874
rect 292 -4942 358 -4908
rect 292 -4976 308 -4942
rect 342 -4976 358 -4942
rect 292 -5010 358 -4976
rect 292 -5044 308 -5010
rect 342 -5044 358 -5010
rect 292 -5078 358 -5044
rect 292 -5112 308 -5078
rect 342 -5112 358 -5078
rect 292 -5146 358 -5112
rect 292 -5180 308 -5146
rect 342 -5180 358 -5146
rect 292 -5214 358 -5180
rect 292 -5248 308 -5214
rect 342 -5248 358 -5214
rect 292 -5282 358 -5248
rect 292 -5316 308 -5282
rect 342 -5316 358 -5282
rect 292 -5350 358 -5316
rect 292 -5384 308 -5350
rect 342 -5384 358 -5350
rect 292 -5418 358 -5384
rect 292 -5452 308 -5418
rect 342 -5452 358 -5418
rect 292 -5486 358 -5452
rect 292 -5520 308 -5486
rect 342 -5520 358 -5486
rect 292 -5563 358 -5520
rect 388 -4806 454 -4763
rect 388 -4840 404 -4806
rect 438 -4840 454 -4806
rect 388 -4874 454 -4840
rect 388 -4908 404 -4874
rect 438 -4908 454 -4874
rect 388 -4942 454 -4908
rect 388 -4976 404 -4942
rect 438 -4976 454 -4942
rect 388 -5010 454 -4976
rect 388 -5044 404 -5010
rect 438 -5044 454 -5010
rect 388 -5078 454 -5044
rect 388 -5112 404 -5078
rect 438 -5112 454 -5078
rect 388 -5146 454 -5112
rect 388 -5180 404 -5146
rect 438 -5180 454 -5146
rect 388 -5214 454 -5180
rect 388 -5248 404 -5214
rect 438 -5248 454 -5214
rect 388 -5282 454 -5248
rect 388 -5316 404 -5282
rect 438 -5316 454 -5282
rect 388 -5350 454 -5316
rect 388 -5384 404 -5350
rect 438 -5384 454 -5350
rect 388 -5418 454 -5384
rect 388 -5452 404 -5418
rect 438 -5452 454 -5418
rect 388 -5486 454 -5452
rect 388 -5520 404 -5486
rect 438 -5520 454 -5486
rect 388 -5563 454 -5520
rect 484 -4806 550 -4763
rect 484 -4840 500 -4806
rect 534 -4840 550 -4806
rect 484 -4874 550 -4840
rect 484 -4908 500 -4874
rect 534 -4908 550 -4874
rect 484 -4942 550 -4908
rect 484 -4976 500 -4942
rect 534 -4976 550 -4942
rect 484 -5010 550 -4976
rect 484 -5044 500 -5010
rect 534 -5044 550 -5010
rect 484 -5078 550 -5044
rect 484 -5112 500 -5078
rect 534 -5112 550 -5078
rect 484 -5146 550 -5112
rect 484 -5180 500 -5146
rect 534 -5180 550 -5146
rect 484 -5214 550 -5180
rect 484 -5248 500 -5214
rect 534 -5248 550 -5214
rect 484 -5282 550 -5248
rect 484 -5316 500 -5282
rect 534 -5316 550 -5282
rect 484 -5350 550 -5316
rect 484 -5384 500 -5350
rect 534 -5384 550 -5350
rect 484 -5418 550 -5384
rect 484 -5452 500 -5418
rect 534 -5452 550 -5418
rect 484 -5486 550 -5452
rect 484 -5520 500 -5486
rect 534 -5520 550 -5486
rect 484 -5563 550 -5520
rect 580 -4806 646 -4763
rect 580 -4840 596 -4806
rect 630 -4840 646 -4806
rect 580 -4874 646 -4840
rect 580 -4908 596 -4874
rect 630 -4908 646 -4874
rect 580 -4942 646 -4908
rect 580 -4976 596 -4942
rect 630 -4976 646 -4942
rect 580 -5010 646 -4976
rect 580 -5044 596 -5010
rect 630 -5044 646 -5010
rect 580 -5078 646 -5044
rect 580 -5112 596 -5078
rect 630 -5112 646 -5078
rect 580 -5146 646 -5112
rect 580 -5180 596 -5146
rect 630 -5180 646 -5146
rect 580 -5214 646 -5180
rect 580 -5248 596 -5214
rect 630 -5248 646 -5214
rect 580 -5282 646 -5248
rect 580 -5316 596 -5282
rect 630 -5316 646 -5282
rect 580 -5350 646 -5316
rect 580 -5384 596 -5350
rect 630 -5384 646 -5350
rect 580 -5418 646 -5384
rect 580 -5452 596 -5418
rect 630 -5452 646 -5418
rect 580 -5486 646 -5452
rect 580 -5520 596 -5486
rect 630 -5520 646 -5486
rect 580 -5563 646 -5520
rect 676 -4806 742 -4763
rect 676 -4840 692 -4806
rect 726 -4840 742 -4806
rect 676 -4874 742 -4840
rect 676 -4908 692 -4874
rect 726 -4908 742 -4874
rect 676 -4942 742 -4908
rect 676 -4976 692 -4942
rect 726 -4976 742 -4942
rect 676 -5010 742 -4976
rect 676 -5044 692 -5010
rect 726 -5044 742 -5010
rect 676 -5078 742 -5044
rect 676 -5112 692 -5078
rect 726 -5112 742 -5078
rect 676 -5146 742 -5112
rect 676 -5180 692 -5146
rect 726 -5180 742 -5146
rect 676 -5214 742 -5180
rect 676 -5248 692 -5214
rect 726 -5248 742 -5214
rect 676 -5282 742 -5248
rect 676 -5316 692 -5282
rect 726 -5316 742 -5282
rect 676 -5350 742 -5316
rect 676 -5384 692 -5350
rect 726 -5384 742 -5350
rect 676 -5418 742 -5384
rect 676 -5452 692 -5418
rect 726 -5452 742 -5418
rect 676 -5486 742 -5452
rect 676 -5520 692 -5486
rect 726 -5520 742 -5486
rect 676 -5563 742 -5520
rect 772 -4806 838 -4763
rect 772 -4840 788 -4806
rect 822 -4840 838 -4806
rect 772 -4874 838 -4840
rect 772 -4908 788 -4874
rect 822 -4908 838 -4874
rect 772 -4942 838 -4908
rect 772 -4976 788 -4942
rect 822 -4976 838 -4942
rect 772 -5010 838 -4976
rect 772 -5044 788 -5010
rect 822 -5044 838 -5010
rect 772 -5078 838 -5044
rect 772 -5112 788 -5078
rect 822 -5112 838 -5078
rect 772 -5146 838 -5112
rect 772 -5180 788 -5146
rect 822 -5180 838 -5146
rect 772 -5214 838 -5180
rect 772 -5248 788 -5214
rect 822 -5248 838 -5214
rect 772 -5282 838 -5248
rect 772 -5316 788 -5282
rect 822 -5316 838 -5282
rect 772 -5350 838 -5316
rect 772 -5384 788 -5350
rect 822 -5384 838 -5350
rect 772 -5418 838 -5384
rect 772 -5452 788 -5418
rect 822 -5452 838 -5418
rect 772 -5486 838 -5452
rect 772 -5520 788 -5486
rect 822 -5520 838 -5486
rect 772 -5563 838 -5520
rect 868 -4806 934 -4763
rect 868 -4840 884 -4806
rect 918 -4840 934 -4806
rect 868 -4874 934 -4840
rect 868 -4908 884 -4874
rect 918 -4908 934 -4874
rect 868 -4942 934 -4908
rect 868 -4976 884 -4942
rect 918 -4976 934 -4942
rect 868 -5010 934 -4976
rect 868 -5044 884 -5010
rect 918 -5044 934 -5010
rect 868 -5078 934 -5044
rect 868 -5112 884 -5078
rect 918 -5112 934 -5078
rect 868 -5146 934 -5112
rect 868 -5180 884 -5146
rect 918 -5180 934 -5146
rect 868 -5214 934 -5180
rect 868 -5248 884 -5214
rect 918 -5248 934 -5214
rect 868 -5282 934 -5248
rect 868 -5316 884 -5282
rect 918 -5316 934 -5282
rect 868 -5350 934 -5316
rect 868 -5384 884 -5350
rect 918 -5384 934 -5350
rect 868 -5418 934 -5384
rect 868 -5452 884 -5418
rect 918 -5452 934 -5418
rect 868 -5486 934 -5452
rect 868 -5520 884 -5486
rect 918 -5520 934 -5486
rect 868 -5563 934 -5520
rect 964 -4806 1030 -4763
rect 964 -4840 980 -4806
rect 1014 -4840 1030 -4806
rect 964 -4874 1030 -4840
rect 964 -4908 980 -4874
rect 1014 -4908 1030 -4874
rect 964 -4942 1030 -4908
rect 964 -4976 980 -4942
rect 1014 -4976 1030 -4942
rect 964 -5010 1030 -4976
rect 964 -5044 980 -5010
rect 1014 -5044 1030 -5010
rect 964 -5078 1030 -5044
rect 964 -5112 980 -5078
rect 1014 -5112 1030 -5078
rect 964 -5146 1030 -5112
rect 964 -5180 980 -5146
rect 1014 -5180 1030 -5146
rect 964 -5214 1030 -5180
rect 964 -5248 980 -5214
rect 1014 -5248 1030 -5214
rect 964 -5282 1030 -5248
rect 964 -5316 980 -5282
rect 1014 -5316 1030 -5282
rect 964 -5350 1030 -5316
rect 964 -5384 980 -5350
rect 1014 -5384 1030 -5350
rect 964 -5418 1030 -5384
rect 964 -5452 980 -5418
rect 1014 -5452 1030 -5418
rect 964 -5486 1030 -5452
rect 964 -5520 980 -5486
rect 1014 -5520 1030 -5486
rect 964 -5563 1030 -5520
rect 1060 -4806 1126 -4763
rect 1060 -4840 1076 -4806
rect 1110 -4840 1126 -4806
rect 1060 -4874 1126 -4840
rect 1060 -4908 1076 -4874
rect 1110 -4908 1126 -4874
rect 1060 -4942 1126 -4908
rect 1060 -4976 1076 -4942
rect 1110 -4976 1126 -4942
rect 1060 -5010 1126 -4976
rect 1060 -5044 1076 -5010
rect 1110 -5044 1126 -5010
rect 1060 -5078 1126 -5044
rect 1060 -5112 1076 -5078
rect 1110 -5112 1126 -5078
rect 1060 -5146 1126 -5112
rect 1060 -5180 1076 -5146
rect 1110 -5180 1126 -5146
rect 1060 -5214 1126 -5180
rect 1060 -5248 1076 -5214
rect 1110 -5248 1126 -5214
rect 1060 -5282 1126 -5248
rect 1060 -5316 1076 -5282
rect 1110 -5316 1126 -5282
rect 1060 -5350 1126 -5316
rect 1060 -5384 1076 -5350
rect 1110 -5384 1126 -5350
rect 1060 -5418 1126 -5384
rect 1060 -5452 1076 -5418
rect 1110 -5452 1126 -5418
rect 1060 -5486 1126 -5452
rect 1060 -5520 1076 -5486
rect 1110 -5520 1126 -5486
rect 1060 -5563 1126 -5520
rect 1156 -4806 1222 -4763
rect 1156 -4840 1172 -4806
rect 1206 -4840 1222 -4806
rect 1156 -4874 1222 -4840
rect 1156 -4908 1172 -4874
rect 1206 -4908 1222 -4874
rect 1156 -4942 1222 -4908
rect 1156 -4976 1172 -4942
rect 1206 -4976 1222 -4942
rect 1156 -5010 1222 -4976
rect 1156 -5044 1172 -5010
rect 1206 -5044 1222 -5010
rect 1156 -5078 1222 -5044
rect 1156 -5112 1172 -5078
rect 1206 -5112 1222 -5078
rect 1156 -5146 1222 -5112
rect 1156 -5180 1172 -5146
rect 1206 -5180 1222 -5146
rect 1156 -5214 1222 -5180
rect 1156 -5248 1172 -5214
rect 1206 -5248 1222 -5214
rect 1156 -5282 1222 -5248
rect 1156 -5316 1172 -5282
rect 1206 -5316 1222 -5282
rect 1156 -5350 1222 -5316
rect 1156 -5384 1172 -5350
rect 1206 -5384 1222 -5350
rect 1156 -5418 1222 -5384
rect 1156 -5452 1172 -5418
rect 1206 -5452 1222 -5418
rect 1156 -5486 1222 -5452
rect 1156 -5520 1172 -5486
rect 1206 -5520 1222 -5486
rect 1156 -5563 1222 -5520
rect 1252 -4806 1318 -4763
rect 1252 -4840 1268 -4806
rect 1302 -4840 1318 -4806
rect 1252 -4874 1318 -4840
rect 1252 -4908 1268 -4874
rect 1302 -4908 1318 -4874
rect 1252 -4942 1318 -4908
rect 1252 -4976 1268 -4942
rect 1302 -4976 1318 -4942
rect 1252 -5010 1318 -4976
rect 1252 -5044 1268 -5010
rect 1302 -5044 1318 -5010
rect 1252 -5078 1318 -5044
rect 1252 -5112 1268 -5078
rect 1302 -5112 1318 -5078
rect 1252 -5146 1318 -5112
rect 1252 -5180 1268 -5146
rect 1302 -5180 1318 -5146
rect 1252 -5214 1318 -5180
rect 1252 -5248 1268 -5214
rect 1302 -5248 1318 -5214
rect 1252 -5282 1318 -5248
rect 1252 -5316 1268 -5282
rect 1302 -5316 1318 -5282
rect 1252 -5350 1318 -5316
rect 1252 -5384 1268 -5350
rect 1302 -5384 1318 -5350
rect 1252 -5418 1318 -5384
rect 1252 -5452 1268 -5418
rect 1302 -5452 1318 -5418
rect 1252 -5486 1318 -5452
rect 1252 -5520 1268 -5486
rect 1302 -5520 1318 -5486
rect 1252 -5563 1318 -5520
rect 1348 -4806 1414 -4763
rect 1348 -4840 1364 -4806
rect 1398 -4840 1414 -4806
rect 1348 -4874 1414 -4840
rect 1348 -4908 1364 -4874
rect 1398 -4908 1414 -4874
rect 1348 -4942 1414 -4908
rect 1348 -4976 1364 -4942
rect 1398 -4976 1414 -4942
rect 1348 -5010 1414 -4976
rect 1348 -5044 1364 -5010
rect 1398 -5044 1414 -5010
rect 1348 -5078 1414 -5044
rect 1348 -5112 1364 -5078
rect 1398 -5112 1414 -5078
rect 1348 -5146 1414 -5112
rect 1348 -5180 1364 -5146
rect 1398 -5180 1414 -5146
rect 1348 -5214 1414 -5180
rect 1348 -5248 1364 -5214
rect 1398 -5248 1414 -5214
rect 1348 -5282 1414 -5248
rect 1348 -5316 1364 -5282
rect 1398 -5316 1414 -5282
rect 1348 -5350 1414 -5316
rect 1348 -5384 1364 -5350
rect 1398 -5384 1414 -5350
rect 1348 -5418 1414 -5384
rect 1348 -5452 1364 -5418
rect 1398 -5452 1414 -5418
rect 1348 -5486 1414 -5452
rect 1348 -5520 1364 -5486
rect 1398 -5520 1414 -5486
rect 1348 -5563 1414 -5520
rect 1444 -4806 1510 -4763
rect 1444 -4840 1460 -4806
rect 1494 -4840 1510 -4806
rect 1444 -4874 1510 -4840
rect 1444 -4908 1460 -4874
rect 1494 -4908 1510 -4874
rect 1444 -4942 1510 -4908
rect 1444 -4976 1460 -4942
rect 1494 -4976 1510 -4942
rect 1444 -5010 1510 -4976
rect 1444 -5044 1460 -5010
rect 1494 -5044 1510 -5010
rect 1444 -5078 1510 -5044
rect 1444 -5112 1460 -5078
rect 1494 -5112 1510 -5078
rect 1444 -5146 1510 -5112
rect 1444 -5180 1460 -5146
rect 1494 -5180 1510 -5146
rect 1444 -5214 1510 -5180
rect 1444 -5248 1460 -5214
rect 1494 -5248 1510 -5214
rect 1444 -5282 1510 -5248
rect 1444 -5316 1460 -5282
rect 1494 -5316 1510 -5282
rect 1444 -5350 1510 -5316
rect 1444 -5384 1460 -5350
rect 1494 -5384 1510 -5350
rect 1444 -5418 1510 -5384
rect 1444 -5452 1460 -5418
rect 1494 -5452 1510 -5418
rect 1444 -5486 1510 -5452
rect 1444 -5520 1460 -5486
rect 1494 -5520 1510 -5486
rect 1444 -5563 1510 -5520
rect 1540 -4806 1606 -4763
rect 1540 -4840 1556 -4806
rect 1590 -4840 1606 -4806
rect 1540 -4874 1606 -4840
rect 1540 -4908 1556 -4874
rect 1590 -4908 1606 -4874
rect 1540 -4942 1606 -4908
rect 1540 -4976 1556 -4942
rect 1590 -4976 1606 -4942
rect 1540 -5010 1606 -4976
rect 1540 -5044 1556 -5010
rect 1590 -5044 1606 -5010
rect 1540 -5078 1606 -5044
rect 1540 -5112 1556 -5078
rect 1590 -5112 1606 -5078
rect 1540 -5146 1606 -5112
rect 1540 -5180 1556 -5146
rect 1590 -5180 1606 -5146
rect 1540 -5214 1606 -5180
rect 1540 -5248 1556 -5214
rect 1590 -5248 1606 -5214
rect 1540 -5282 1606 -5248
rect 1540 -5316 1556 -5282
rect 1590 -5316 1606 -5282
rect 1540 -5350 1606 -5316
rect 1540 -5384 1556 -5350
rect 1590 -5384 1606 -5350
rect 1540 -5418 1606 -5384
rect 1540 -5452 1556 -5418
rect 1590 -5452 1606 -5418
rect 1540 -5486 1606 -5452
rect 1540 -5520 1556 -5486
rect 1590 -5520 1606 -5486
rect 1540 -5563 1606 -5520
rect 1636 -4806 1702 -4763
rect 1636 -4840 1652 -4806
rect 1686 -4840 1702 -4806
rect 1636 -4874 1702 -4840
rect 1636 -4908 1652 -4874
rect 1686 -4908 1702 -4874
rect 1636 -4942 1702 -4908
rect 1636 -4976 1652 -4942
rect 1686 -4976 1702 -4942
rect 1636 -5010 1702 -4976
rect 1636 -5044 1652 -5010
rect 1686 -5044 1702 -5010
rect 1636 -5078 1702 -5044
rect 1636 -5112 1652 -5078
rect 1686 -5112 1702 -5078
rect 1636 -5146 1702 -5112
rect 1636 -5180 1652 -5146
rect 1686 -5180 1702 -5146
rect 1636 -5214 1702 -5180
rect 1636 -5248 1652 -5214
rect 1686 -5248 1702 -5214
rect 1636 -5282 1702 -5248
rect 1636 -5316 1652 -5282
rect 1686 -5316 1702 -5282
rect 1636 -5350 1702 -5316
rect 1636 -5384 1652 -5350
rect 1686 -5384 1702 -5350
rect 1636 -5418 1702 -5384
rect 1636 -5452 1652 -5418
rect 1686 -5452 1702 -5418
rect 1636 -5486 1702 -5452
rect 1636 -5520 1652 -5486
rect 1686 -5520 1702 -5486
rect 1636 -5563 1702 -5520
rect 1732 -4806 1798 -4763
rect 1732 -4840 1748 -4806
rect 1782 -4840 1798 -4806
rect 1732 -4874 1798 -4840
rect 1732 -4908 1748 -4874
rect 1782 -4908 1798 -4874
rect 1732 -4942 1798 -4908
rect 1732 -4976 1748 -4942
rect 1782 -4976 1798 -4942
rect 1732 -5010 1798 -4976
rect 1732 -5044 1748 -5010
rect 1782 -5044 1798 -5010
rect 1732 -5078 1798 -5044
rect 1732 -5112 1748 -5078
rect 1782 -5112 1798 -5078
rect 1732 -5146 1798 -5112
rect 1732 -5180 1748 -5146
rect 1782 -5180 1798 -5146
rect 1732 -5214 1798 -5180
rect 1732 -5248 1748 -5214
rect 1782 -5248 1798 -5214
rect 1732 -5282 1798 -5248
rect 1732 -5316 1748 -5282
rect 1782 -5316 1798 -5282
rect 1732 -5350 1798 -5316
rect 1732 -5384 1748 -5350
rect 1782 -5384 1798 -5350
rect 1732 -5418 1798 -5384
rect 1732 -5452 1748 -5418
rect 1782 -5452 1798 -5418
rect 1732 -5486 1798 -5452
rect 1732 -5520 1748 -5486
rect 1782 -5520 1798 -5486
rect 1732 -5563 1798 -5520
rect 1828 -4806 1894 -4763
rect 1828 -4840 1844 -4806
rect 1878 -4840 1894 -4806
rect 1828 -4874 1894 -4840
rect 1828 -4908 1844 -4874
rect 1878 -4908 1894 -4874
rect 1828 -4942 1894 -4908
rect 1828 -4976 1844 -4942
rect 1878 -4976 1894 -4942
rect 1828 -5010 1894 -4976
rect 1828 -5044 1844 -5010
rect 1878 -5044 1894 -5010
rect 1828 -5078 1894 -5044
rect 1828 -5112 1844 -5078
rect 1878 -5112 1894 -5078
rect 1828 -5146 1894 -5112
rect 1828 -5180 1844 -5146
rect 1878 -5180 1894 -5146
rect 1828 -5214 1894 -5180
rect 1828 -5248 1844 -5214
rect 1878 -5248 1894 -5214
rect 1828 -5282 1894 -5248
rect 1828 -5316 1844 -5282
rect 1878 -5316 1894 -5282
rect 1828 -5350 1894 -5316
rect 1828 -5384 1844 -5350
rect 1878 -5384 1894 -5350
rect 1828 -5418 1894 -5384
rect 1828 -5452 1844 -5418
rect 1878 -5452 1894 -5418
rect 1828 -5486 1894 -5452
rect 1828 -5520 1844 -5486
rect 1878 -5520 1894 -5486
rect 1828 -5563 1894 -5520
rect 1924 -4806 1986 -4763
rect 1924 -4840 1940 -4806
rect 1974 -4840 1986 -4806
rect 1924 -4874 1986 -4840
rect 1924 -4908 1940 -4874
rect 1974 -4908 1986 -4874
rect 1924 -4942 1986 -4908
rect 1924 -4976 1940 -4942
rect 1974 -4976 1986 -4942
rect 1924 -5010 1986 -4976
rect 1924 -5044 1940 -5010
rect 1974 -5044 1986 -5010
rect 1924 -5078 1986 -5044
rect 1924 -5112 1940 -5078
rect 1974 -5112 1986 -5078
rect 1924 -5146 1986 -5112
rect 1924 -5180 1940 -5146
rect 1974 -5180 1986 -5146
rect 1924 -5214 1986 -5180
rect 1924 -5248 1940 -5214
rect 1974 -5248 1986 -5214
rect 1924 -5282 1986 -5248
rect 1924 -5316 1940 -5282
rect 1974 -5316 1986 -5282
rect 1924 -5350 1986 -5316
rect 1924 -5384 1940 -5350
rect 1974 -5384 1986 -5350
rect 1924 -5418 1986 -5384
rect 1924 -5452 1940 -5418
rect 1974 -5452 1986 -5418
rect 1924 -5486 1986 -5452
rect 1924 -5520 1940 -5486
rect 1974 -5520 1986 -5486
rect 1924 -5563 1986 -5520
<< pdiff >>
rect -50459 33299 -50401 33312
rect -50459 33265 -50447 33299
rect -50413 33265 -50401 33299
rect -50459 33231 -50401 33265
rect -50459 33197 -50447 33231
rect -50413 33197 -50401 33231
rect -50459 33163 -50401 33197
rect -50459 33129 -50447 33163
rect -50413 33129 -50401 33163
rect -50459 33095 -50401 33129
rect -50459 33061 -50447 33095
rect -50413 33061 -50401 33095
rect -50459 33027 -50401 33061
rect -50459 32993 -50447 33027
rect -50413 32993 -50401 33027
rect -50459 32959 -50401 32993
rect -50459 32925 -50447 32959
rect -50413 32925 -50401 32959
rect -50459 32912 -50401 32925
rect -50301 33299 -50243 33312
rect -50301 33265 -50289 33299
rect -50255 33265 -50243 33299
rect -50301 33231 -50243 33265
rect -50301 33197 -50289 33231
rect -50255 33197 -50243 33231
rect -50301 33163 -50243 33197
rect -50301 33129 -50289 33163
rect -50255 33129 -50243 33163
rect -50301 33095 -50243 33129
rect -50301 33061 -50289 33095
rect -50255 33061 -50243 33095
rect -50301 33027 -50243 33061
rect -50301 32993 -50289 33027
rect -50255 32993 -50243 33027
rect -50301 32959 -50243 32993
rect -50301 32925 -50289 32959
rect -50255 32925 -50243 32959
rect -50301 32912 -50243 32925
rect -50143 33299 -50085 33312
rect -50143 33265 -50131 33299
rect -50097 33265 -50085 33299
rect -50143 33231 -50085 33265
rect -50143 33197 -50131 33231
rect -50097 33197 -50085 33231
rect -50143 33163 -50085 33197
rect -50143 33129 -50131 33163
rect -50097 33129 -50085 33163
rect -50143 33095 -50085 33129
rect -50143 33061 -50131 33095
rect -50097 33061 -50085 33095
rect -50143 33027 -50085 33061
rect -50143 32993 -50131 33027
rect -50097 32993 -50085 33027
rect -50143 32959 -50085 32993
rect -50143 32925 -50131 32959
rect -50097 32925 -50085 32959
rect -50143 32912 -50085 32925
rect -49985 33299 -49927 33312
rect -49985 33265 -49973 33299
rect -49939 33265 -49927 33299
rect -49985 33231 -49927 33265
rect -49985 33197 -49973 33231
rect -49939 33197 -49927 33231
rect -49985 33163 -49927 33197
rect -49985 33129 -49973 33163
rect -49939 33129 -49927 33163
rect -49985 33095 -49927 33129
rect -49985 33061 -49973 33095
rect -49939 33061 -49927 33095
rect -49985 33027 -49927 33061
rect -49985 32993 -49973 33027
rect -49939 32993 -49927 33027
rect -49985 32959 -49927 32993
rect -49985 32925 -49973 32959
rect -49939 32925 -49927 32959
rect -49985 32912 -49927 32925
rect -49827 33299 -49769 33312
rect -49827 33265 -49815 33299
rect -49781 33265 -49769 33299
rect -49827 33231 -49769 33265
rect -49827 33197 -49815 33231
rect -49781 33197 -49769 33231
rect -49827 33163 -49769 33197
rect -49827 33129 -49815 33163
rect -49781 33129 -49769 33163
rect -49827 33095 -49769 33129
rect -49827 33061 -49815 33095
rect -49781 33061 -49769 33095
rect -49827 33027 -49769 33061
rect -49827 32993 -49815 33027
rect -49781 32993 -49769 33027
rect -49827 32959 -49769 32993
rect -49827 32925 -49815 32959
rect -49781 32925 -49769 32959
rect -49827 32912 -49769 32925
rect -49669 33299 -49611 33312
rect -49669 33265 -49657 33299
rect -49623 33265 -49611 33299
rect -49669 33231 -49611 33265
rect -49669 33197 -49657 33231
rect -49623 33197 -49611 33231
rect -49669 33163 -49611 33197
rect -49669 33129 -49657 33163
rect -49623 33129 -49611 33163
rect -49669 33095 -49611 33129
rect -49669 33061 -49657 33095
rect -49623 33061 -49611 33095
rect -49669 33027 -49611 33061
rect -49669 32993 -49657 33027
rect -49623 32993 -49611 33027
rect -49669 32959 -49611 32993
rect -49669 32925 -49657 32959
rect -49623 32925 -49611 32959
rect -49669 32912 -49611 32925
rect -49511 33299 -49453 33312
rect -49511 33265 -49499 33299
rect -49465 33265 -49453 33299
rect -49511 33231 -49453 33265
rect -49511 33197 -49499 33231
rect -49465 33197 -49453 33231
rect -49511 33163 -49453 33197
rect -49511 33129 -49499 33163
rect -49465 33129 -49453 33163
rect -49511 33095 -49453 33129
rect -49511 33061 -49499 33095
rect -49465 33061 -49453 33095
rect -49511 33027 -49453 33061
rect -49511 32993 -49499 33027
rect -49465 32993 -49453 33027
rect -49511 32959 -49453 32993
rect -49511 32925 -49499 32959
rect -49465 32925 -49453 32959
rect -49511 32912 -49453 32925
rect -49353 33299 -49295 33312
rect -49353 33265 -49341 33299
rect -49307 33265 -49295 33299
rect -49353 33231 -49295 33265
rect -49353 33197 -49341 33231
rect -49307 33197 -49295 33231
rect -49353 33163 -49295 33197
rect -49353 33129 -49341 33163
rect -49307 33129 -49295 33163
rect -49353 33095 -49295 33129
rect -49353 33061 -49341 33095
rect -49307 33061 -49295 33095
rect -49353 33027 -49295 33061
rect -49353 32993 -49341 33027
rect -49307 32993 -49295 33027
rect -49353 32959 -49295 32993
rect -49353 32925 -49341 32959
rect -49307 32925 -49295 32959
rect -49353 32912 -49295 32925
rect -49195 33299 -49137 33312
rect -49195 33265 -49183 33299
rect -49149 33265 -49137 33299
rect -49195 33231 -49137 33265
rect -49195 33197 -49183 33231
rect -49149 33197 -49137 33231
rect -49195 33163 -49137 33197
rect -49195 33129 -49183 33163
rect -49149 33129 -49137 33163
rect -49195 33095 -49137 33129
rect -49195 33061 -49183 33095
rect -49149 33061 -49137 33095
rect -49195 33027 -49137 33061
rect -49195 32993 -49183 33027
rect -49149 32993 -49137 33027
rect -49195 32959 -49137 32993
rect -49195 32925 -49183 32959
rect -49149 32925 -49137 32959
rect -49195 32912 -49137 32925
rect -49037 33299 -48979 33312
rect -49037 33265 -49025 33299
rect -48991 33265 -48979 33299
rect -49037 33231 -48979 33265
rect -49037 33197 -49025 33231
rect -48991 33197 -48979 33231
rect -49037 33163 -48979 33197
rect -49037 33129 -49025 33163
rect -48991 33129 -48979 33163
rect -49037 33095 -48979 33129
rect -49037 33061 -49025 33095
rect -48991 33061 -48979 33095
rect -49037 33027 -48979 33061
rect -49037 32993 -49025 33027
rect -48991 32993 -48979 33027
rect -49037 32959 -48979 32993
rect -49037 32925 -49025 32959
rect -48991 32925 -48979 32959
rect -49037 32912 -48979 32925
rect -48879 33299 -48821 33312
rect -48879 33265 -48867 33299
rect -48833 33265 -48821 33299
rect -48879 33231 -48821 33265
rect -48879 33197 -48867 33231
rect -48833 33197 -48821 33231
rect -48879 33163 -48821 33197
rect -48879 33129 -48867 33163
rect -48833 33129 -48821 33163
rect -48879 33095 -48821 33129
rect -48879 33061 -48867 33095
rect -48833 33061 -48821 33095
rect -48879 33027 -48821 33061
rect -48879 32993 -48867 33027
rect -48833 32993 -48821 33027
rect -48879 32959 -48821 32993
rect -48879 32925 -48867 32959
rect -48833 32925 -48821 32959
rect -48879 32912 -48821 32925
rect 2888 33299 2946 33312
rect 2888 33265 2900 33299
rect 2934 33265 2946 33299
rect 2888 33231 2946 33265
rect 2888 33197 2900 33231
rect 2934 33197 2946 33231
rect 2888 33163 2946 33197
rect 2888 33129 2900 33163
rect 2934 33129 2946 33163
rect 2888 33095 2946 33129
rect 2888 33061 2900 33095
rect 2934 33061 2946 33095
rect 2888 33027 2946 33061
rect 2888 32993 2900 33027
rect 2934 32993 2946 33027
rect 2888 32959 2946 32993
rect 2888 32925 2900 32959
rect 2934 32925 2946 32959
rect 2888 32912 2946 32925
rect 3046 33299 3104 33312
rect 3046 33265 3058 33299
rect 3092 33265 3104 33299
rect 3046 33231 3104 33265
rect 3046 33197 3058 33231
rect 3092 33197 3104 33231
rect 3046 33163 3104 33197
rect 3046 33129 3058 33163
rect 3092 33129 3104 33163
rect 3046 33095 3104 33129
rect 3046 33061 3058 33095
rect 3092 33061 3104 33095
rect 3046 33027 3104 33061
rect 3046 32993 3058 33027
rect 3092 32993 3104 33027
rect 3046 32959 3104 32993
rect 3046 32925 3058 32959
rect 3092 32925 3104 32959
rect 3046 32912 3104 32925
rect 3204 33299 3262 33312
rect 3204 33265 3216 33299
rect 3250 33265 3262 33299
rect 3204 33231 3262 33265
rect 3204 33197 3216 33231
rect 3250 33197 3262 33231
rect 3204 33163 3262 33197
rect 3204 33129 3216 33163
rect 3250 33129 3262 33163
rect 3204 33095 3262 33129
rect 3204 33061 3216 33095
rect 3250 33061 3262 33095
rect 3204 33027 3262 33061
rect 3204 32993 3216 33027
rect 3250 32993 3262 33027
rect 3204 32959 3262 32993
rect 3204 32925 3216 32959
rect 3250 32925 3262 32959
rect 3204 32912 3262 32925
rect 3362 33299 3420 33312
rect 3362 33265 3374 33299
rect 3408 33265 3420 33299
rect 3362 33231 3420 33265
rect 3362 33197 3374 33231
rect 3408 33197 3420 33231
rect 3362 33163 3420 33197
rect 3362 33129 3374 33163
rect 3408 33129 3420 33163
rect 3362 33095 3420 33129
rect 3362 33061 3374 33095
rect 3408 33061 3420 33095
rect 3362 33027 3420 33061
rect 3362 32993 3374 33027
rect 3408 32993 3420 33027
rect 3362 32959 3420 32993
rect 3362 32925 3374 32959
rect 3408 32925 3420 32959
rect 3362 32912 3420 32925
rect 3520 33299 3578 33312
rect 3520 33265 3532 33299
rect 3566 33265 3578 33299
rect 3520 33231 3578 33265
rect 3520 33197 3532 33231
rect 3566 33197 3578 33231
rect 3520 33163 3578 33197
rect 3520 33129 3532 33163
rect 3566 33129 3578 33163
rect 3520 33095 3578 33129
rect 3520 33061 3532 33095
rect 3566 33061 3578 33095
rect 3520 33027 3578 33061
rect 3520 32993 3532 33027
rect 3566 32993 3578 33027
rect 3520 32959 3578 32993
rect 3520 32925 3532 32959
rect 3566 32925 3578 32959
rect 3520 32912 3578 32925
rect 3678 33299 3736 33312
rect 3678 33265 3690 33299
rect 3724 33265 3736 33299
rect 3678 33231 3736 33265
rect 3678 33197 3690 33231
rect 3724 33197 3736 33231
rect 3678 33163 3736 33197
rect 3678 33129 3690 33163
rect 3724 33129 3736 33163
rect 3678 33095 3736 33129
rect 3678 33061 3690 33095
rect 3724 33061 3736 33095
rect 3678 33027 3736 33061
rect 3678 32993 3690 33027
rect 3724 32993 3736 33027
rect 3678 32959 3736 32993
rect 3678 32925 3690 32959
rect 3724 32925 3736 32959
rect 3678 32912 3736 32925
rect 3836 33299 3894 33312
rect 3836 33265 3848 33299
rect 3882 33265 3894 33299
rect 3836 33231 3894 33265
rect 3836 33197 3848 33231
rect 3882 33197 3894 33231
rect 3836 33163 3894 33197
rect 3836 33129 3848 33163
rect 3882 33129 3894 33163
rect 3836 33095 3894 33129
rect 3836 33061 3848 33095
rect 3882 33061 3894 33095
rect 3836 33027 3894 33061
rect 3836 32993 3848 33027
rect 3882 32993 3894 33027
rect 3836 32959 3894 32993
rect 3836 32925 3848 32959
rect 3882 32925 3894 32959
rect 3836 32912 3894 32925
rect 3994 33299 4052 33312
rect 3994 33265 4006 33299
rect 4040 33265 4052 33299
rect 3994 33231 4052 33265
rect 3994 33197 4006 33231
rect 4040 33197 4052 33231
rect 3994 33163 4052 33197
rect 3994 33129 4006 33163
rect 4040 33129 4052 33163
rect 3994 33095 4052 33129
rect 3994 33061 4006 33095
rect 4040 33061 4052 33095
rect 3994 33027 4052 33061
rect 3994 32993 4006 33027
rect 4040 32993 4052 33027
rect 3994 32959 4052 32993
rect 3994 32925 4006 32959
rect 4040 32925 4052 32959
rect 3994 32912 4052 32925
rect 4152 33299 4210 33312
rect 4152 33265 4164 33299
rect 4198 33265 4210 33299
rect 4152 33231 4210 33265
rect 4152 33197 4164 33231
rect 4198 33197 4210 33231
rect 4152 33163 4210 33197
rect 4152 33129 4164 33163
rect 4198 33129 4210 33163
rect 4152 33095 4210 33129
rect 4152 33061 4164 33095
rect 4198 33061 4210 33095
rect 4152 33027 4210 33061
rect 4152 32993 4164 33027
rect 4198 32993 4210 33027
rect 4152 32959 4210 32993
rect 4152 32925 4164 32959
rect 4198 32925 4210 32959
rect 4152 32912 4210 32925
rect 4310 33299 4368 33312
rect 4310 33265 4322 33299
rect 4356 33265 4368 33299
rect 4310 33231 4368 33265
rect 4310 33197 4322 33231
rect 4356 33197 4368 33231
rect 4310 33163 4368 33197
rect 4310 33129 4322 33163
rect 4356 33129 4368 33163
rect 4310 33095 4368 33129
rect 4310 33061 4322 33095
rect 4356 33061 4368 33095
rect 4310 33027 4368 33061
rect 4310 32993 4322 33027
rect 4356 32993 4368 33027
rect 4310 32959 4368 32993
rect 4310 32925 4322 32959
rect 4356 32925 4368 32959
rect 4310 32912 4368 32925
rect 4468 33299 4526 33312
rect 4468 33265 4480 33299
rect 4514 33265 4526 33299
rect 4468 33231 4526 33265
rect 4468 33197 4480 33231
rect 4514 33197 4526 33231
rect 4468 33163 4526 33197
rect 4468 33129 4480 33163
rect 4514 33129 4526 33163
rect 4468 33095 4526 33129
rect 4468 33061 4480 33095
rect 4514 33061 4526 33095
rect 4468 33027 4526 33061
rect 4468 32993 4480 33027
rect 4514 32993 4526 33027
rect 4468 32959 4526 32993
rect 4468 32925 4480 32959
rect 4514 32925 4526 32959
rect 4468 32912 4526 32925
<< ndiffc >>
rect -50447 32606 -50413 32640
rect -50447 32538 -50413 32572
rect -50447 32470 -50413 32504
rect -50289 32606 -50255 32640
rect -50289 32538 -50255 32572
rect -50289 32470 -50255 32504
rect -50131 32606 -50097 32640
rect -50131 32538 -50097 32572
rect -50131 32470 -50097 32504
rect -49973 32606 -49939 32640
rect -49973 32538 -49939 32572
rect -49973 32470 -49939 32504
rect -49815 32606 -49781 32640
rect -49815 32538 -49781 32572
rect -49815 32470 -49781 32504
rect -49657 32606 -49623 32640
rect -49657 32538 -49623 32572
rect -49657 32470 -49623 32504
rect -49499 32606 -49465 32640
rect -49499 32538 -49465 32572
rect -49499 32470 -49465 32504
rect -49341 32606 -49307 32640
rect -49341 32538 -49307 32572
rect -49341 32470 -49307 32504
rect -49183 32606 -49149 32640
rect -49183 32538 -49149 32572
rect -49183 32470 -49149 32504
rect -49025 32606 -48991 32640
rect -49025 32538 -48991 32572
rect -49025 32470 -48991 32504
rect -48867 32606 -48833 32640
rect -48867 32538 -48833 32572
rect -48867 32470 -48833 32504
rect 2900 32606 2934 32640
rect 2900 32538 2934 32572
rect 2900 32470 2934 32504
rect 3058 32606 3092 32640
rect 3058 32538 3092 32572
rect 3058 32470 3092 32504
rect 3216 32606 3250 32640
rect 3216 32538 3250 32572
rect 3216 32470 3250 32504
rect 3374 32606 3408 32640
rect 3374 32538 3408 32572
rect 3374 32470 3408 32504
rect 3532 32606 3566 32640
rect 3532 32538 3566 32572
rect 3532 32470 3566 32504
rect 3690 32606 3724 32640
rect 3690 32538 3724 32572
rect 3690 32470 3724 32504
rect 3848 32606 3882 32640
rect 3848 32538 3882 32572
rect 3848 32470 3882 32504
rect 4006 32606 4040 32640
rect 4006 32538 4040 32572
rect 4006 32470 4040 32504
rect 4164 32606 4198 32640
rect 4164 32538 4198 32572
rect 4164 32470 4198 32504
rect 4322 32606 4356 32640
rect 4322 32538 4356 32572
rect 4322 32470 4356 32504
rect 4480 32606 4514 32640
rect 4480 32538 4514 32572
rect 4480 32470 4514 32504
rect -42524 5360 -42490 5394
rect -42524 5292 -42490 5326
rect -42524 5224 -42490 5258
rect -42524 5156 -42490 5190
rect -42524 5088 -42490 5122
rect -42524 5020 -42490 5054
rect -42524 4952 -42490 4986
rect -42524 4884 -42490 4918
rect -42524 4816 -42490 4850
rect -42524 4748 -42490 4782
rect -42524 4680 -42490 4714
rect -42428 5360 -42394 5394
rect -42428 5292 -42394 5326
rect -42428 5224 -42394 5258
rect -42428 5156 -42394 5190
rect -42428 5088 -42394 5122
rect -42428 5020 -42394 5054
rect -42428 4952 -42394 4986
rect -42428 4884 -42394 4918
rect -42428 4816 -42394 4850
rect -42428 4748 -42394 4782
rect -42428 4680 -42394 4714
rect -42332 5360 -42298 5394
rect -42332 5292 -42298 5326
rect -42332 5224 -42298 5258
rect -42332 5156 -42298 5190
rect -42332 5088 -42298 5122
rect -42332 5020 -42298 5054
rect -42332 4952 -42298 4986
rect -42332 4884 -42298 4918
rect -42332 4816 -42298 4850
rect -42332 4748 -42298 4782
rect -42332 4680 -42298 4714
rect -42236 5360 -42202 5394
rect -42236 5292 -42202 5326
rect -42236 5224 -42202 5258
rect -42236 5156 -42202 5190
rect -42236 5088 -42202 5122
rect -42236 5020 -42202 5054
rect -42236 4952 -42202 4986
rect -42236 4884 -42202 4918
rect -42236 4816 -42202 4850
rect -42236 4748 -42202 4782
rect -42236 4680 -42202 4714
rect -42140 5360 -42106 5394
rect -42140 5292 -42106 5326
rect -42140 5224 -42106 5258
rect -42140 5156 -42106 5190
rect -42140 5088 -42106 5122
rect -42140 5020 -42106 5054
rect -42140 4952 -42106 4986
rect -42140 4884 -42106 4918
rect -42140 4816 -42106 4850
rect -42140 4748 -42106 4782
rect -42140 4680 -42106 4714
rect -42044 5360 -42010 5394
rect -42044 5292 -42010 5326
rect -42044 5224 -42010 5258
rect -42044 5156 -42010 5190
rect -42044 5088 -42010 5122
rect -42044 5020 -42010 5054
rect -42044 4952 -42010 4986
rect -42044 4884 -42010 4918
rect -42044 4816 -42010 4850
rect -42044 4748 -42010 4782
rect -42044 4680 -42010 4714
rect -41948 5360 -41914 5394
rect -41948 5292 -41914 5326
rect -41948 5224 -41914 5258
rect -41948 5156 -41914 5190
rect -41948 5088 -41914 5122
rect -41948 5020 -41914 5054
rect -41948 4952 -41914 4986
rect -41948 4884 -41914 4918
rect -41948 4816 -41914 4850
rect -41948 4748 -41914 4782
rect -41948 4680 -41914 4714
rect -41852 5360 -41818 5394
rect -41852 5292 -41818 5326
rect -41852 5224 -41818 5258
rect -41852 5156 -41818 5190
rect -41852 5088 -41818 5122
rect -41852 5020 -41818 5054
rect -41852 4952 -41818 4986
rect -41852 4884 -41818 4918
rect -41852 4816 -41818 4850
rect -41852 4748 -41818 4782
rect -41852 4680 -41818 4714
rect -41756 5360 -41722 5394
rect -41756 5292 -41722 5326
rect -41756 5224 -41722 5258
rect -41756 5156 -41722 5190
rect -41756 5088 -41722 5122
rect -41756 5020 -41722 5054
rect -41756 4952 -41722 4986
rect -41756 4884 -41722 4918
rect -41756 4816 -41722 4850
rect -41756 4748 -41722 4782
rect -41756 4680 -41722 4714
rect -41660 5360 -41626 5394
rect -41660 5292 -41626 5326
rect -41660 5224 -41626 5258
rect -41660 5156 -41626 5190
rect -41660 5088 -41626 5122
rect -41660 5020 -41626 5054
rect -41660 4952 -41626 4986
rect -41660 4884 -41626 4918
rect -41660 4816 -41626 4850
rect -41660 4748 -41626 4782
rect -41660 4680 -41626 4714
rect -41564 5360 -41530 5394
rect -41564 5292 -41530 5326
rect -41564 5224 -41530 5258
rect -41564 5156 -41530 5190
rect -41564 5088 -41530 5122
rect -41564 5020 -41530 5054
rect -41564 4952 -41530 4986
rect -41564 4884 -41530 4918
rect -41564 4816 -41530 4850
rect -41564 4748 -41530 4782
rect -41564 4680 -41530 4714
rect -41468 5360 -41434 5394
rect -41468 5292 -41434 5326
rect -41468 5224 -41434 5258
rect -41468 5156 -41434 5190
rect -41468 5088 -41434 5122
rect -41468 5020 -41434 5054
rect -41468 4952 -41434 4986
rect -41468 4884 -41434 4918
rect -41468 4816 -41434 4850
rect -41468 4748 -41434 4782
rect -41468 4680 -41434 4714
rect -41372 5360 -41338 5394
rect -41372 5292 -41338 5326
rect -41372 5224 -41338 5258
rect -41372 5156 -41338 5190
rect -41372 5088 -41338 5122
rect -41372 5020 -41338 5054
rect -41372 4952 -41338 4986
rect -41372 4884 -41338 4918
rect -41372 4816 -41338 4850
rect -41372 4748 -41338 4782
rect -41372 4680 -41338 4714
rect -41276 5360 -41242 5394
rect -41276 5292 -41242 5326
rect -41276 5224 -41242 5258
rect -41276 5156 -41242 5190
rect -41276 5088 -41242 5122
rect -41276 5020 -41242 5054
rect -41276 4952 -41242 4986
rect -41276 4884 -41242 4918
rect -41276 4816 -41242 4850
rect -41276 4748 -41242 4782
rect -41276 4680 -41242 4714
rect -41180 5360 -41146 5394
rect -41180 5292 -41146 5326
rect -41180 5224 -41146 5258
rect -41180 5156 -41146 5190
rect -41180 5088 -41146 5122
rect -41180 5020 -41146 5054
rect -41180 4952 -41146 4986
rect -41180 4884 -41146 4918
rect -41180 4816 -41146 4850
rect -41180 4748 -41146 4782
rect -41180 4680 -41146 4714
rect -41084 5360 -41050 5394
rect -41084 5292 -41050 5326
rect -41084 5224 -41050 5258
rect -41084 5156 -41050 5190
rect -41084 5088 -41050 5122
rect -41084 5020 -41050 5054
rect -41084 4952 -41050 4986
rect -41084 4884 -41050 4918
rect -41084 4816 -41050 4850
rect -41084 4748 -41050 4782
rect -41084 4680 -41050 4714
rect -40988 5360 -40954 5394
rect -40988 5292 -40954 5326
rect -40988 5224 -40954 5258
rect -40988 5156 -40954 5190
rect -40988 5088 -40954 5122
rect -40988 5020 -40954 5054
rect -40988 4952 -40954 4986
rect -40988 4884 -40954 4918
rect -40988 4816 -40954 4850
rect -40988 4748 -40954 4782
rect -40988 4680 -40954 4714
rect -40892 5360 -40858 5394
rect -40892 5292 -40858 5326
rect -40892 5224 -40858 5258
rect -40892 5156 -40858 5190
rect -40892 5088 -40858 5122
rect -40892 5020 -40858 5054
rect -40892 4952 -40858 4986
rect -40892 4884 -40858 4918
rect -40892 4816 -40858 4850
rect -40892 4748 -40858 4782
rect -40892 4680 -40858 4714
rect -40796 5360 -40762 5394
rect -40796 5292 -40762 5326
rect -40796 5224 -40762 5258
rect -40796 5156 -40762 5190
rect -40796 5088 -40762 5122
rect -40796 5020 -40762 5054
rect -40796 4952 -40762 4986
rect -40796 4884 -40762 4918
rect -40796 4816 -40762 4850
rect -40796 4748 -40762 4782
rect -40796 4680 -40762 4714
rect -40700 5360 -40666 5394
rect -40700 5292 -40666 5326
rect -40700 5224 -40666 5258
rect -40700 5156 -40666 5190
rect -40700 5088 -40666 5122
rect -40700 5020 -40666 5054
rect -40700 4952 -40666 4986
rect -40700 4884 -40666 4918
rect -40700 4816 -40666 4850
rect -40700 4748 -40666 4782
rect -40700 4680 -40666 4714
rect 104 5348 138 5382
rect 104 5280 138 5314
rect 104 5212 138 5246
rect 104 5144 138 5178
rect 104 5076 138 5110
rect 104 5008 138 5042
rect 104 4940 138 4974
rect 104 4872 138 4906
rect 104 4804 138 4838
rect 104 4736 138 4770
rect 104 4668 138 4702
rect 200 5348 234 5382
rect 200 5280 234 5314
rect 200 5212 234 5246
rect 200 5144 234 5178
rect 200 5076 234 5110
rect 200 5008 234 5042
rect 200 4940 234 4974
rect 200 4872 234 4906
rect 200 4804 234 4838
rect 200 4736 234 4770
rect 200 4668 234 4702
rect 296 5348 330 5382
rect 296 5280 330 5314
rect 296 5212 330 5246
rect 296 5144 330 5178
rect 296 5076 330 5110
rect 296 5008 330 5042
rect 296 4940 330 4974
rect 296 4872 330 4906
rect 296 4804 330 4838
rect 296 4736 330 4770
rect 296 4668 330 4702
rect 392 5348 426 5382
rect 392 5280 426 5314
rect 392 5212 426 5246
rect 392 5144 426 5178
rect 392 5076 426 5110
rect 392 5008 426 5042
rect 392 4940 426 4974
rect 392 4872 426 4906
rect 392 4804 426 4838
rect 392 4736 426 4770
rect 392 4668 426 4702
rect 488 5348 522 5382
rect 488 5280 522 5314
rect 488 5212 522 5246
rect 488 5144 522 5178
rect 488 5076 522 5110
rect 488 5008 522 5042
rect 488 4940 522 4974
rect 488 4872 522 4906
rect 488 4804 522 4838
rect 488 4736 522 4770
rect 488 4668 522 4702
rect 584 5348 618 5382
rect 584 5280 618 5314
rect 584 5212 618 5246
rect 584 5144 618 5178
rect 584 5076 618 5110
rect 584 5008 618 5042
rect 584 4940 618 4974
rect 584 4872 618 4906
rect 584 4804 618 4838
rect 584 4736 618 4770
rect 584 4668 618 4702
rect 680 5348 714 5382
rect 680 5280 714 5314
rect 680 5212 714 5246
rect 680 5144 714 5178
rect 680 5076 714 5110
rect 680 5008 714 5042
rect 680 4940 714 4974
rect 680 4872 714 4906
rect 680 4804 714 4838
rect 680 4736 714 4770
rect 680 4668 714 4702
rect 776 5348 810 5382
rect 776 5280 810 5314
rect 776 5212 810 5246
rect 776 5144 810 5178
rect 776 5076 810 5110
rect 776 5008 810 5042
rect 776 4940 810 4974
rect 776 4872 810 4906
rect 776 4804 810 4838
rect 776 4736 810 4770
rect 776 4668 810 4702
rect 872 5348 906 5382
rect 872 5280 906 5314
rect 872 5212 906 5246
rect 872 5144 906 5178
rect 872 5076 906 5110
rect 872 5008 906 5042
rect 872 4940 906 4974
rect 872 4872 906 4906
rect 872 4804 906 4838
rect 872 4736 906 4770
rect 872 4668 906 4702
rect 968 5348 1002 5382
rect 968 5280 1002 5314
rect 968 5212 1002 5246
rect 968 5144 1002 5178
rect 968 5076 1002 5110
rect 968 5008 1002 5042
rect 968 4940 1002 4974
rect 968 4872 1002 4906
rect 968 4804 1002 4838
rect 968 4736 1002 4770
rect 968 4668 1002 4702
rect 1064 5348 1098 5382
rect 1064 5280 1098 5314
rect 1064 5212 1098 5246
rect 1064 5144 1098 5178
rect 1064 5076 1098 5110
rect 1064 5008 1098 5042
rect 1064 4940 1098 4974
rect 1064 4872 1098 4906
rect 1064 4804 1098 4838
rect 1064 4736 1098 4770
rect 1064 4668 1098 4702
rect 1160 5348 1194 5382
rect 1160 5280 1194 5314
rect 1160 5212 1194 5246
rect 1160 5144 1194 5178
rect 1160 5076 1194 5110
rect 1160 5008 1194 5042
rect 1160 4940 1194 4974
rect 1160 4872 1194 4906
rect 1160 4804 1194 4838
rect 1160 4736 1194 4770
rect 1160 4668 1194 4702
rect 1256 5348 1290 5382
rect 1256 5280 1290 5314
rect 1256 5212 1290 5246
rect 1256 5144 1290 5178
rect 1256 5076 1290 5110
rect 1256 5008 1290 5042
rect 1256 4940 1290 4974
rect 1256 4872 1290 4906
rect 1256 4804 1290 4838
rect 1256 4736 1290 4770
rect 1256 4668 1290 4702
rect 1352 5348 1386 5382
rect 1352 5280 1386 5314
rect 1352 5212 1386 5246
rect 1352 5144 1386 5178
rect 1352 5076 1386 5110
rect 1352 5008 1386 5042
rect 1352 4940 1386 4974
rect 1352 4872 1386 4906
rect 1352 4804 1386 4838
rect 1352 4736 1386 4770
rect 1352 4668 1386 4702
rect 1448 5348 1482 5382
rect 1448 5280 1482 5314
rect 1448 5212 1482 5246
rect 1448 5144 1482 5178
rect 1448 5076 1482 5110
rect 1448 5008 1482 5042
rect 1448 4940 1482 4974
rect 1448 4872 1482 4906
rect 1448 4804 1482 4838
rect 1448 4736 1482 4770
rect 1448 4668 1482 4702
rect 1544 5348 1578 5382
rect 1544 5280 1578 5314
rect 1544 5212 1578 5246
rect 1544 5144 1578 5178
rect 1544 5076 1578 5110
rect 1544 5008 1578 5042
rect 1544 4940 1578 4974
rect 1544 4872 1578 4906
rect 1544 4804 1578 4838
rect 1544 4736 1578 4770
rect 1544 4668 1578 4702
rect 1640 5348 1674 5382
rect 1640 5280 1674 5314
rect 1640 5212 1674 5246
rect 1640 5144 1674 5178
rect 1640 5076 1674 5110
rect 1640 5008 1674 5042
rect 1640 4940 1674 4974
rect 1640 4872 1674 4906
rect 1640 4804 1674 4838
rect 1640 4736 1674 4770
rect 1640 4668 1674 4702
rect 1736 5348 1770 5382
rect 1736 5280 1770 5314
rect 1736 5212 1770 5246
rect 1736 5144 1770 5178
rect 1736 5076 1770 5110
rect 1736 5008 1770 5042
rect 1736 4940 1770 4974
rect 1736 4872 1770 4906
rect 1736 4804 1770 4838
rect 1736 4736 1770 4770
rect 1736 4668 1770 4702
rect 1832 5348 1866 5382
rect 1832 5280 1866 5314
rect 1832 5212 1866 5246
rect 1832 5144 1866 5178
rect 1832 5076 1866 5110
rect 1832 5008 1866 5042
rect 1832 4940 1866 4974
rect 1832 4872 1866 4906
rect 1832 4804 1866 4838
rect 1832 4736 1866 4770
rect 1832 4668 1866 4702
rect 1928 5348 1962 5382
rect 1928 5280 1962 5314
rect 1928 5212 1962 5246
rect 1928 5144 1962 5178
rect 1928 5076 1962 5110
rect 1928 5008 1962 5042
rect 1928 4940 1962 4974
rect 1928 4872 1962 4906
rect 1928 4804 1962 4838
rect 1928 4736 1962 4770
rect 1928 4668 1962 4702
rect -42525 -4814 -42491 -4780
rect -42525 -4882 -42491 -4848
rect -42525 -4950 -42491 -4916
rect -42525 -5018 -42491 -4984
rect -42525 -5086 -42491 -5052
rect -42525 -5154 -42491 -5120
rect -42525 -5222 -42491 -5188
rect -42525 -5290 -42491 -5256
rect -42525 -5358 -42491 -5324
rect -42525 -5426 -42491 -5392
rect -42525 -5494 -42491 -5460
rect -42429 -4814 -42395 -4780
rect -42429 -4882 -42395 -4848
rect -42429 -4950 -42395 -4916
rect -42429 -5018 -42395 -4984
rect -42429 -5086 -42395 -5052
rect -42429 -5154 -42395 -5120
rect -42429 -5222 -42395 -5188
rect -42429 -5290 -42395 -5256
rect -42429 -5358 -42395 -5324
rect -42429 -5426 -42395 -5392
rect -42429 -5494 -42395 -5460
rect -42333 -4814 -42299 -4780
rect -42333 -4882 -42299 -4848
rect -42333 -4950 -42299 -4916
rect -42333 -5018 -42299 -4984
rect -42333 -5086 -42299 -5052
rect -42333 -5154 -42299 -5120
rect -42333 -5222 -42299 -5188
rect -42333 -5290 -42299 -5256
rect -42333 -5358 -42299 -5324
rect -42333 -5426 -42299 -5392
rect -42333 -5494 -42299 -5460
rect -42237 -4814 -42203 -4780
rect -42237 -4882 -42203 -4848
rect -42237 -4950 -42203 -4916
rect -42237 -5018 -42203 -4984
rect -42237 -5086 -42203 -5052
rect -42237 -5154 -42203 -5120
rect -42237 -5222 -42203 -5188
rect -42237 -5290 -42203 -5256
rect -42237 -5358 -42203 -5324
rect -42237 -5426 -42203 -5392
rect -42237 -5494 -42203 -5460
rect -42141 -4814 -42107 -4780
rect -42141 -4882 -42107 -4848
rect -42141 -4950 -42107 -4916
rect -42141 -5018 -42107 -4984
rect -42141 -5086 -42107 -5052
rect -42141 -5154 -42107 -5120
rect -42141 -5222 -42107 -5188
rect -42141 -5290 -42107 -5256
rect -42141 -5358 -42107 -5324
rect -42141 -5426 -42107 -5392
rect -42141 -5494 -42107 -5460
rect -42045 -4814 -42011 -4780
rect -42045 -4882 -42011 -4848
rect -42045 -4950 -42011 -4916
rect -42045 -5018 -42011 -4984
rect -42045 -5086 -42011 -5052
rect -42045 -5154 -42011 -5120
rect -42045 -5222 -42011 -5188
rect -42045 -5290 -42011 -5256
rect -42045 -5358 -42011 -5324
rect -42045 -5426 -42011 -5392
rect -42045 -5494 -42011 -5460
rect -41949 -4814 -41915 -4780
rect -41949 -4882 -41915 -4848
rect -41949 -4950 -41915 -4916
rect -41949 -5018 -41915 -4984
rect -41949 -5086 -41915 -5052
rect -41949 -5154 -41915 -5120
rect -41949 -5222 -41915 -5188
rect -41949 -5290 -41915 -5256
rect -41949 -5358 -41915 -5324
rect -41949 -5426 -41915 -5392
rect -41949 -5494 -41915 -5460
rect -41853 -4814 -41819 -4780
rect -41853 -4882 -41819 -4848
rect -41853 -4950 -41819 -4916
rect -41853 -5018 -41819 -4984
rect -41853 -5086 -41819 -5052
rect -41853 -5154 -41819 -5120
rect -41853 -5222 -41819 -5188
rect -41853 -5290 -41819 -5256
rect -41853 -5358 -41819 -5324
rect -41853 -5426 -41819 -5392
rect -41853 -5494 -41819 -5460
rect -41757 -4814 -41723 -4780
rect -41757 -4882 -41723 -4848
rect -41757 -4950 -41723 -4916
rect -41757 -5018 -41723 -4984
rect -41757 -5086 -41723 -5052
rect -41757 -5154 -41723 -5120
rect -41757 -5222 -41723 -5188
rect -41757 -5290 -41723 -5256
rect -41757 -5358 -41723 -5324
rect -41757 -5426 -41723 -5392
rect -41757 -5494 -41723 -5460
rect -41661 -4814 -41627 -4780
rect -41661 -4882 -41627 -4848
rect -41661 -4950 -41627 -4916
rect -41661 -5018 -41627 -4984
rect -41661 -5086 -41627 -5052
rect -41661 -5154 -41627 -5120
rect -41661 -5222 -41627 -5188
rect -41661 -5290 -41627 -5256
rect -41661 -5358 -41627 -5324
rect -41661 -5426 -41627 -5392
rect -41661 -5494 -41627 -5460
rect -41565 -4814 -41531 -4780
rect -41565 -4882 -41531 -4848
rect -41565 -4950 -41531 -4916
rect -41565 -5018 -41531 -4984
rect -41565 -5086 -41531 -5052
rect -41565 -5154 -41531 -5120
rect -41565 -5222 -41531 -5188
rect -41565 -5290 -41531 -5256
rect -41565 -5358 -41531 -5324
rect -41565 -5426 -41531 -5392
rect -41565 -5494 -41531 -5460
rect -41469 -4814 -41435 -4780
rect -41469 -4882 -41435 -4848
rect -41469 -4950 -41435 -4916
rect -41469 -5018 -41435 -4984
rect -41469 -5086 -41435 -5052
rect -41469 -5154 -41435 -5120
rect -41469 -5222 -41435 -5188
rect -41469 -5290 -41435 -5256
rect -41469 -5358 -41435 -5324
rect -41469 -5426 -41435 -5392
rect -41469 -5494 -41435 -5460
rect -41373 -4814 -41339 -4780
rect -41373 -4882 -41339 -4848
rect -41373 -4950 -41339 -4916
rect -41373 -5018 -41339 -4984
rect -41373 -5086 -41339 -5052
rect -41373 -5154 -41339 -5120
rect -41373 -5222 -41339 -5188
rect -41373 -5290 -41339 -5256
rect -41373 -5358 -41339 -5324
rect -41373 -5426 -41339 -5392
rect -41373 -5494 -41339 -5460
rect -41277 -4814 -41243 -4780
rect -41277 -4882 -41243 -4848
rect -41277 -4950 -41243 -4916
rect -41277 -5018 -41243 -4984
rect -41277 -5086 -41243 -5052
rect -41277 -5154 -41243 -5120
rect -41277 -5222 -41243 -5188
rect -41277 -5290 -41243 -5256
rect -41277 -5358 -41243 -5324
rect -41277 -5426 -41243 -5392
rect -41277 -5494 -41243 -5460
rect -41181 -4814 -41147 -4780
rect -41181 -4882 -41147 -4848
rect -41181 -4950 -41147 -4916
rect -41181 -5018 -41147 -4984
rect -41181 -5086 -41147 -5052
rect -41181 -5154 -41147 -5120
rect -41181 -5222 -41147 -5188
rect -41181 -5290 -41147 -5256
rect -41181 -5358 -41147 -5324
rect -41181 -5426 -41147 -5392
rect -41181 -5494 -41147 -5460
rect -41085 -4814 -41051 -4780
rect -41085 -4882 -41051 -4848
rect -41085 -4950 -41051 -4916
rect -41085 -5018 -41051 -4984
rect -41085 -5086 -41051 -5052
rect -41085 -5154 -41051 -5120
rect -41085 -5222 -41051 -5188
rect -41085 -5290 -41051 -5256
rect -41085 -5358 -41051 -5324
rect -41085 -5426 -41051 -5392
rect -41085 -5494 -41051 -5460
rect -40989 -4814 -40955 -4780
rect -40989 -4882 -40955 -4848
rect -40989 -4950 -40955 -4916
rect -40989 -5018 -40955 -4984
rect -40989 -5086 -40955 -5052
rect -40989 -5154 -40955 -5120
rect -40989 -5222 -40955 -5188
rect -40989 -5290 -40955 -5256
rect -40989 -5358 -40955 -5324
rect -40989 -5426 -40955 -5392
rect -40989 -5494 -40955 -5460
rect -40893 -4814 -40859 -4780
rect -40893 -4882 -40859 -4848
rect -40893 -4950 -40859 -4916
rect -40893 -5018 -40859 -4984
rect -40893 -5086 -40859 -5052
rect -40893 -5154 -40859 -5120
rect -40893 -5222 -40859 -5188
rect -40893 -5290 -40859 -5256
rect -40893 -5358 -40859 -5324
rect -40893 -5426 -40859 -5392
rect -40893 -5494 -40859 -5460
rect -40797 -4814 -40763 -4780
rect -40797 -4882 -40763 -4848
rect -40797 -4950 -40763 -4916
rect -40797 -5018 -40763 -4984
rect -40797 -5086 -40763 -5052
rect -40797 -5154 -40763 -5120
rect -40797 -5222 -40763 -5188
rect -40797 -5290 -40763 -5256
rect -40797 -5358 -40763 -5324
rect -40797 -5426 -40763 -5392
rect -40797 -5494 -40763 -5460
rect -40701 -4814 -40667 -4780
rect -40701 -4882 -40667 -4848
rect -40701 -4950 -40667 -4916
rect -40701 -5018 -40667 -4984
rect -40701 -5086 -40667 -5052
rect -40701 -5154 -40667 -5120
rect -40701 -5222 -40667 -5188
rect -40701 -5290 -40667 -5256
rect -40701 -5358 -40667 -5324
rect -40701 -5426 -40667 -5392
rect -40701 -5494 -40667 -5460
rect 116 -4840 150 -4806
rect 116 -4908 150 -4874
rect 116 -4976 150 -4942
rect 116 -5044 150 -5010
rect 116 -5112 150 -5078
rect 116 -5180 150 -5146
rect 116 -5248 150 -5214
rect 116 -5316 150 -5282
rect 116 -5384 150 -5350
rect 116 -5452 150 -5418
rect 116 -5520 150 -5486
rect 212 -4840 246 -4806
rect 212 -4908 246 -4874
rect 212 -4976 246 -4942
rect 212 -5044 246 -5010
rect 212 -5112 246 -5078
rect 212 -5180 246 -5146
rect 212 -5248 246 -5214
rect 212 -5316 246 -5282
rect 212 -5384 246 -5350
rect 212 -5452 246 -5418
rect 212 -5520 246 -5486
rect 308 -4840 342 -4806
rect 308 -4908 342 -4874
rect 308 -4976 342 -4942
rect 308 -5044 342 -5010
rect 308 -5112 342 -5078
rect 308 -5180 342 -5146
rect 308 -5248 342 -5214
rect 308 -5316 342 -5282
rect 308 -5384 342 -5350
rect 308 -5452 342 -5418
rect 308 -5520 342 -5486
rect 404 -4840 438 -4806
rect 404 -4908 438 -4874
rect 404 -4976 438 -4942
rect 404 -5044 438 -5010
rect 404 -5112 438 -5078
rect 404 -5180 438 -5146
rect 404 -5248 438 -5214
rect 404 -5316 438 -5282
rect 404 -5384 438 -5350
rect 404 -5452 438 -5418
rect 404 -5520 438 -5486
rect 500 -4840 534 -4806
rect 500 -4908 534 -4874
rect 500 -4976 534 -4942
rect 500 -5044 534 -5010
rect 500 -5112 534 -5078
rect 500 -5180 534 -5146
rect 500 -5248 534 -5214
rect 500 -5316 534 -5282
rect 500 -5384 534 -5350
rect 500 -5452 534 -5418
rect 500 -5520 534 -5486
rect 596 -4840 630 -4806
rect 596 -4908 630 -4874
rect 596 -4976 630 -4942
rect 596 -5044 630 -5010
rect 596 -5112 630 -5078
rect 596 -5180 630 -5146
rect 596 -5248 630 -5214
rect 596 -5316 630 -5282
rect 596 -5384 630 -5350
rect 596 -5452 630 -5418
rect 596 -5520 630 -5486
rect 692 -4840 726 -4806
rect 692 -4908 726 -4874
rect 692 -4976 726 -4942
rect 692 -5044 726 -5010
rect 692 -5112 726 -5078
rect 692 -5180 726 -5146
rect 692 -5248 726 -5214
rect 692 -5316 726 -5282
rect 692 -5384 726 -5350
rect 692 -5452 726 -5418
rect 692 -5520 726 -5486
rect 788 -4840 822 -4806
rect 788 -4908 822 -4874
rect 788 -4976 822 -4942
rect 788 -5044 822 -5010
rect 788 -5112 822 -5078
rect 788 -5180 822 -5146
rect 788 -5248 822 -5214
rect 788 -5316 822 -5282
rect 788 -5384 822 -5350
rect 788 -5452 822 -5418
rect 788 -5520 822 -5486
rect 884 -4840 918 -4806
rect 884 -4908 918 -4874
rect 884 -4976 918 -4942
rect 884 -5044 918 -5010
rect 884 -5112 918 -5078
rect 884 -5180 918 -5146
rect 884 -5248 918 -5214
rect 884 -5316 918 -5282
rect 884 -5384 918 -5350
rect 884 -5452 918 -5418
rect 884 -5520 918 -5486
rect 980 -4840 1014 -4806
rect 980 -4908 1014 -4874
rect 980 -4976 1014 -4942
rect 980 -5044 1014 -5010
rect 980 -5112 1014 -5078
rect 980 -5180 1014 -5146
rect 980 -5248 1014 -5214
rect 980 -5316 1014 -5282
rect 980 -5384 1014 -5350
rect 980 -5452 1014 -5418
rect 980 -5520 1014 -5486
rect 1076 -4840 1110 -4806
rect 1076 -4908 1110 -4874
rect 1076 -4976 1110 -4942
rect 1076 -5044 1110 -5010
rect 1076 -5112 1110 -5078
rect 1076 -5180 1110 -5146
rect 1076 -5248 1110 -5214
rect 1076 -5316 1110 -5282
rect 1076 -5384 1110 -5350
rect 1076 -5452 1110 -5418
rect 1076 -5520 1110 -5486
rect 1172 -4840 1206 -4806
rect 1172 -4908 1206 -4874
rect 1172 -4976 1206 -4942
rect 1172 -5044 1206 -5010
rect 1172 -5112 1206 -5078
rect 1172 -5180 1206 -5146
rect 1172 -5248 1206 -5214
rect 1172 -5316 1206 -5282
rect 1172 -5384 1206 -5350
rect 1172 -5452 1206 -5418
rect 1172 -5520 1206 -5486
rect 1268 -4840 1302 -4806
rect 1268 -4908 1302 -4874
rect 1268 -4976 1302 -4942
rect 1268 -5044 1302 -5010
rect 1268 -5112 1302 -5078
rect 1268 -5180 1302 -5146
rect 1268 -5248 1302 -5214
rect 1268 -5316 1302 -5282
rect 1268 -5384 1302 -5350
rect 1268 -5452 1302 -5418
rect 1268 -5520 1302 -5486
rect 1364 -4840 1398 -4806
rect 1364 -4908 1398 -4874
rect 1364 -4976 1398 -4942
rect 1364 -5044 1398 -5010
rect 1364 -5112 1398 -5078
rect 1364 -5180 1398 -5146
rect 1364 -5248 1398 -5214
rect 1364 -5316 1398 -5282
rect 1364 -5384 1398 -5350
rect 1364 -5452 1398 -5418
rect 1364 -5520 1398 -5486
rect 1460 -4840 1494 -4806
rect 1460 -4908 1494 -4874
rect 1460 -4976 1494 -4942
rect 1460 -5044 1494 -5010
rect 1460 -5112 1494 -5078
rect 1460 -5180 1494 -5146
rect 1460 -5248 1494 -5214
rect 1460 -5316 1494 -5282
rect 1460 -5384 1494 -5350
rect 1460 -5452 1494 -5418
rect 1460 -5520 1494 -5486
rect 1556 -4840 1590 -4806
rect 1556 -4908 1590 -4874
rect 1556 -4976 1590 -4942
rect 1556 -5044 1590 -5010
rect 1556 -5112 1590 -5078
rect 1556 -5180 1590 -5146
rect 1556 -5248 1590 -5214
rect 1556 -5316 1590 -5282
rect 1556 -5384 1590 -5350
rect 1556 -5452 1590 -5418
rect 1556 -5520 1590 -5486
rect 1652 -4840 1686 -4806
rect 1652 -4908 1686 -4874
rect 1652 -4976 1686 -4942
rect 1652 -5044 1686 -5010
rect 1652 -5112 1686 -5078
rect 1652 -5180 1686 -5146
rect 1652 -5248 1686 -5214
rect 1652 -5316 1686 -5282
rect 1652 -5384 1686 -5350
rect 1652 -5452 1686 -5418
rect 1652 -5520 1686 -5486
rect 1748 -4840 1782 -4806
rect 1748 -4908 1782 -4874
rect 1748 -4976 1782 -4942
rect 1748 -5044 1782 -5010
rect 1748 -5112 1782 -5078
rect 1748 -5180 1782 -5146
rect 1748 -5248 1782 -5214
rect 1748 -5316 1782 -5282
rect 1748 -5384 1782 -5350
rect 1748 -5452 1782 -5418
rect 1748 -5520 1782 -5486
rect 1844 -4840 1878 -4806
rect 1844 -4908 1878 -4874
rect 1844 -4976 1878 -4942
rect 1844 -5044 1878 -5010
rect 1844 -5112 1878 -5078
rect 1844 -5180 1878 -5146
rect 1844 -5248 1878 -5214
rect 1844 -5316 1878 -5282
rect 1844 -5384 1878 -5350
rect 1844 -5452 1878 -5418
rect 1844 -5520 1878 -5486
rect 1940 -4840 1974 -4806
rect 1940 -4908 1974 -4874
rect 1940 -4976 1974 -4942
rect 1940 -5044 1974 -5010
rect 1940 -5112 1974 -5078
rect 1940 -5180 1974 -5146
rect 1940 -5248 1974 -5214
rect 1940 -5316 1974 -5282
rect 1940 -5384 1974 -5350
rect 1940 -5452 1974 -5418
rect 1940 -5520 1974 -5486
<< pdiffc >>
rect -50447 33265 -50413 33299
rect -50447 33197 -50413 33231
rect -50447 33129 -50413 33163
rect -50447 33061 -50413 33095
rect -50447 32993 -50413 33027
rect -50447 32925 -50413 32959
rect -50289 33265 -50255 33299
rect -50289 33197 -50255 33231
rect -50289 33129 -50255 33163
rect -50289 33061 -50255 33095
rect -50289 32993 -50255 33027
rect -50289 32925 -50255 32959
rect -50131 33265 -50097 33299
rect -50131 33197 -50097 33231
rect -50131 33129 -50097 33163
rect -50131 33061 -50097 33095
rect -50131 32993 -50097 33027
rect -50131 32925 -50097 32959
rect -49973 33265 -49939 33299
rect -49973 33197 -49939 33231
rect -49973 33129 -49939 33163
rect -49973 33061 -49939 33095
rect -49973 32993 -49939 33027
rect -49973 32925 -49939 32959
rect -49815 33265 -49781 33299
rect -49815 33197 -49781 33231
rect -49815 33129 -49781 33163
rect -49815 33061 -49781 33095
rect -49815 32993 -49781 33027
rect -49815 32925 -49781 32959
rect -49657 33265 -49623 33299
rect -49657 33197 -49623 33231
rect -49657 33129 -49623 33163
rect -49657 33061 -49623 33095
rect -49657 32993 -49623 33027
rect -49657 32925 -49623 32959
rect -49499 33265 -49465 33299
rect -49499 33197 -49465 33231
rect -49499 33129 -49465 33163
rect -49499 33061 -49465 33095
rect -49499 32993 -49465 33027
rect -49499 32925 -49465 32959
rect -49341 33265 -49307 33299
rect -49341 33197 -49307 33231
rect -49341 33129 -49307 33163
rect -49341 33061 -49307 33095
rect -49341 32993 -49307 33027
rect -49341 32925 -49307 32959
rect -49183 33265 -49149 33299
rect -49183 33197 -49149 33231
rect -49183 33129 -49149 33163
rect -49183 33061 -49149 33095
rect -49183 32993 -49149 33027
rect -49183 32925 -49149 32959
rect -49025 33265 -48991 33299
rect -49025 33197 -48991 33231
rect -49025 33129 -48991 33163
rect -49025 33061 -48991 33095
rect -49025 32993 -48991 33027
rect -49025 32925 -48991 32959
rect -48867 33265 -48833 33299
rect -48867 33197 -48833 33231
rect -48867 33129 -48833 33163
rect -48867 33061 -48833 33095
rect -48867 32993 -48833 33027
rect -48867 32925 -48833 32959
rect 2900 33265 2934 33299
rect 2900 33197 2934 33231
rect 2900 33129 2934 33163
rect 2900 33061 2934 33095
rect 2900 32993 2934 33027
rect 2900 32925 2934 32959
rect 3058 33265 3092 33299
rect 3058 33197 3092 33231
rect 3058 33129 3092 33163
rect 3058 33061 3092 33095
rect 3058 32993 3092 33027
rect 3058 32925 3092 32959
rect 3216 33265 3250 33299
rect 3216 33197 3250 33231
rect 3216 33129 3250 33163
rect 3216 33061 3250 33095
rect 3216 32993 3250 33027
rect 3216 32925 3250 32959
rect 3374 33265 3408 33299
rect 3374 33197 3408 33231
rect 3374 33129 3408 33163
rect 3374 33061 3408 33095
rect 3374 32993 3408 33027
rect 3374 32925 3408 32959
rect 3532 33265 3566 33299
rect 3532 33197 3566 33231
rect 3532 33129 3566 33163
rect 3532 33061 3566 33095
rect 3532 32993 3566 33027
rect 3532 32925 3566 32959
rect 3690 33265 3724 33299
rect 3690 33197 3724 33231
rect 3690 33129 3724 33163
rect 3690 33061 3724 33095
rect 3690 32993 3724 33027
rect 3690 32925 3724 32959
rect 3848 33265 3882 33299
rect 3848 33197 3882 33231
rect 3848 33129 3882 33163
rect 3848 33061 3882 33095
rect 3848 32993 3882 33027
rect 3848 32925 3882 32959
rect 4006 33265 4040 33299
rect 4006 33197 4040 33231
rect 4006 33129 4040 33163
rect 4006 33061 4040 33095
rect 4006 32993 4040 33027
rect 4006 32925 4040 32959
rect 4164 33265 4198 33299
rect 4164 33197 4198 33231
rect 4164 33129 4198 33163
rect 4164 33061 4198 33095
rect 4164 32993 4198 33027
rect 4164 32925 4198 32959
rect 4322 33265 4356 33299
rect 4322 33197 4356 33231
rect 4322 33129 4356 33163
rect 4322 33061 4356 33095
rect 4322 32993 4356 33027
rect 4322 32925 4356 32959
rect 4480 33265 4514 33299
rect 4480 33197 4514 33231
rect 4480 33129 4514 33163
rect 4480 33061 4514 33095
rect 4480 32993 4514 33027
rect 4480 32925 4514 32959
<< psubdiff >>
rect 2023 32635 2119 32669
rect 2153 32635 2187 32669
rect 2221 32635 2317 32669
rect 2023 32573 2057 32635
rect 2283 32573 2317 32635
rect 2023 32505 2057 32539
rect 2283 32505 2317 32539
rect 2023 32409 2057 32471
rect 2283 32409 2317 32471
rect 2023 32375 2119 32409
rect 2153 32375 2187 32409
rect 2221 32375 2317 32409
rect -50473 32349 -48807 32373
rect -50473 32315 -50449 32349
rect -50415 32315 -50377 32349
rect -50343 32315 -50305 32349
rect -50271 32315 -50233 32349
rect -50199 32315 -50161 32349
rect -50127 32315 -50089 32349
rect -50055 32315 -50017 32349
rect -49983 32315 -49945 32349
rect -49911 32315 -49873 32349
rect -49839 32315 -49801 32349
rect -49767 32315 -49729 32349
rect -49695 32315 -49657 32349
rect -49623 32315 -49585 32349
rect -49551 32315 -49513 32349
rect -49479 32315 -49441 32349
rect -49407 32315 -49369 32349
rect -49335 32315 -49297 32349
rect -49263 32315 -49225 32349
rect -49191 32315 -49153 32349
rect -49119 32315 -49081 32349
rect -49047 32315 -49009 32349
rect -48975 32315 -48937 32349
rect -48903 32315 -48865 32349
rect -48831 32315 -48807 32349
rect -50473 32277 -48807 32315
rect -50473 32243 -50449 32277
rect -50415 32243 -50377 32277
rect -50343 32243 -50305 32277
rect -50271 32243 -50233 32277
rect -50199 32243 -50161 32277
rect -50127 32243 -50089 32277
rect -50055 32243 -50017 32277
rect -49983 32243 -49945 32277
rect -49911 32243 -49873 32277
rect -49839 32243 -49801 32277
rect -49767 32243 -49729 32277
rect -49695 32243 -49657 32277
rect -49623 32243 -49585 32277
rect -49551 32243 -49513 32277
rect -49479 32243 -49441 32277
rect -49407 32243 -49369 32277
rect -49335 32243 -49297 32277
rect -49263 32243 -49225 32277
rect -49191 32243 -49153 32277
rect -49119 32243 -49081 32277
rect -49047 32243 -49009 32277
rect -48975 32243 -48937 32277
rect -48903 32243 -48865 32277
rect -48831 32243 -48807 32277
rect -50473 32219 -48807 32243
rect 2874 32349 4540 32373
rect 2874 32315 2898 32349
rect 2932 32315 2970 32349
rect 3004 32315 3042 32349
rect 3076 32315 3114 32349
rect 3148 32315 3186 32349
rect 3220 32315 3258 32349
rect 3292 32315 3330 32349
rect 3364 32315 3402 32349
rect 3436 32315 3474 32349
rect 3508 32315 3546 32349
rect 3580 32315 3618 32349
rect 3652 32315 3690 32349
rect 3724 32315 3762 32349
rect 3796 32315 3834 32349
rect 3868 32315 3906 32349
rect 3940 32315 3978 32349
rect 4012 32315 4050 32349
rect 4084 32315 4122 32349
rect 4156 32315 4194 32349
rect 4228 32315 4266 32349
rect 4300 32315 4338 32349
rect 4372 32315 4410 32349
rect 4444 32315 4482 32349
rect 4516 32315 4540 32349
rect 2874 32277 4540 32315
rect 2874 32243 2898 32277
rect 2932 32243 2970 32277
rect 3004 32243 3042 32277
rect 3076 32243 3114 32277
rect 3148 32243 3186 32277
rect 3220 32243 3258 32277
rect 3292 32243 3330 32277
rect 3364 32243 3402 32277
rect 3436 32243 3474 32277
rect 3508 32243 3546 32277
rect 3580 32243 3618 32277
rect 3652 32243 3690 32277
rect 3724 32243 3762 32277
rect 3796 32243 3834 32277
rect 3868 32243 3906 32277
rect 3940 32243 3978 32277
rect 4012 32243 4050 32277
rect 4084 32243 4122 32277
rect 4156 32243 4194 32277
rect 4228 32243 4266 32277
rect 4300 32243 4338 32277
rect 4372 32243 4410 32277
rect 4444 32243 4482 32277
rect 4516 32243 4540 32277
rect 2874 32219 4540 32243
rect -50899 32131 -50803 32165
rect -50769 32131 -50735 32165
rect -50701 32131 -50605 32165
rect -50899 32069 -50865 32131
rect -50639 32069 -50605 32131
rect -50899 32001 -50865 32035
rect -50639 32001 -50605 32035
rect -50899 31905 -50865 31967
rect -50639 31905 -50605 31967
rect -50899 31871 -50803 31905
rect -50769 31871 -50735 31905
rect -50701 31871 -50605 31905
<< nsubdiff >>
rect -50473 33524 -48807 33548
rect -50473 33490 -50449 33524
rect -50415 33490 -50377 33524
rect -50343 33490 -50305 33524
rect -50271 33490 -50233 33524
rect -50199 33490 -50161 33524
rect -50127 33490 -50089 33524
rect -50055 33490 -50017 33524
rect -49983 33490 -49945 33524
rect -49911 33490 -49873 33524
rect -49839 33490 -49801 33524
rect -49767 33490 -49729 33524
rect -49695 33490 -49657 33524
rect -49623 33490 -49585 33524
rect -49551 33490 -49513 33524
rect -49479 33490 -49441 33524
rect -49407 33490 -49369 33524
rect -49335 33490 -49297 33524
rect -49263 33490 -49225 33524
rect -49191 33490 -49153 33524
rect -49119 33490 -49081 33524
rect -49047 33490 -49009 33524
rect -48975 33490 -48937 33524
rect -48903 33490 -48865 33524
rect -48831 33490 -48807 33524
rect -50473 33452 -48807 33490
rect -50473 33418 -50449 33452
rect -50415 33418 -50377 33452
rect -50343 33418 -50305 33452
rect -50271 33418 -50233 33452
rect -50199 33418 -50161 33452
rect -50127 33418 -50089 33452
rect -50055 33418 -50017 33452
rect -49983 33418 -49945 33452
rect -49911 33418 -49873 33452
rect -49839 33418 -49801 33452
rect -49767 33418 -49729 33452
rect -49695 33418 -49657 33452
rect -49623 33418 -49585 33452
rect -49551 33418 -49513 33452
rect -49479 33418 -49441 33452
rect -49407 33418 -49369 33452
rect -49335 33418 -49297 33452
rect -49263 33418 -49225 33452
rect -49191 33418 -49153 33452
rect -49119 33418 -49081 33452
rect -49047 33418 -49009 33452
rect -48975 33418 -48937 33452
rect -48903 33418 -48865 33452
rect -48831 33418 -48807 33452
rect -50473 33394 -48807 33418
rect 2874 33524 4540 33548
rect 2874 33490 2898 33524
rect 2932 33490 2970 33524
rect 3004 33490 3042 33524
rect 3076 33490 3114 33524
rect 3148 33490 3186 33524
rect 3220 33490 3258 33524
rect 3292 33490 3330 33524
rect 3364 33490 3402 33524
rect 3436 33490 3474 33524
rect 3508 33490 3546 33524
rect 3580 33490 3618 33524
rect 3652 33490 3690 33524
rect 3724 33490 3762 33524
rect 3796 33490 3834 33524
rect 3868 33490 3906 33524
rect 3940 33490 3978 33524
rect 4012 33490 4050 33524
rect 4084 33490 4122 33524
rect 4156 33490 4194 33524
rect 4228 33490 4266 33524
rect 4300 33490 4338 33524
rect 4372 33490 4410 33524
rect 4444 33490 4482 33524
rect 4516 33490 4540 33524
rect 2874 33452 4540 33490
rect 2874 33418 2898 33452
rect 2932 33418 2970 33452
rect 3004 33418 3042 33452
rect 3076 33418 3114 33452
rect 3148 33418 3186 33452
rect 3220 33418 3258 33452
rect 3292 33418 3330 33452
rect 3364 33418 3402 33452
rect 3436 33418 3474 33452
rect 3508 33418 3546 33452
rect 3580 33418 3618 33452
rect 3652 33418 3690 33452
rect 3724 33418 3762 33452
rect 3796 33418 3834 33452
rect 3868 33418 3906 33452
rect 3940 33418 3978 33452
rect 4012 33418 4050 33452
rect 4084 33418 4122 33452
rect 4156 33418 4194 33452
rect 4228 33418 4266 33452
rect 4300 33418 4338 33452
rect 4372 33418 4410 33452
rect 4444 33418 4482 33452
rect 4516 33418 4540 33452
rect 2874 33394 4540 33418
<< psubdiffcont >>
rect 2119 32635 2153 32669
rect 2187 32635 2221 32669
rect 2023 32539 2057 32573
rect 2023 32471 2057 32505
rect 2283 32539 2317 32573
rect 2283 32471 2317 32505
rect 2119 32375 2153 32409
rect 2187 32375 2221 32409
rect -50449 32315 -50415 32349
rect -50377 32315 -50343 32349
rect -50305 32315 -50271 32349
rect -50233 32315 -50199 32349
rect -50161 32315 -50127 32349
rect -50089 32315 -50055 32349
rect -50017 32315 -49983 32349
rect -49945 32315 -49911 32349
rect -49873 32315 -49839 32349
rect -49801 32315 -49767 32349
rect -49729 32315 -49695 32349
rect -49657 32315 -49623 32349
rect -49585 32315 -49551 32349
rect -49513 32315 -49479 32349
rect -49441 32315 -49407 32349
rect -49369 32315 -49335 32349
rect -49297 32315 -49263 32349
rect -49225 32315 -49191 32349
rect -49153 32315 -49119 32349
rect -49081 32315 -49047 32349
rect -49009 32315 -48975 32349
rect -48937 32315 -48903 32349
rect -48865 32315 -48831 32349
rect -50449 32243 -50415 32277
rect -50377 32243 -50343 32277
rect -50305 32243 -50271 32277
rect -50233 32243 -50199 32277
rect -50161 32243 -50127 32277
rect -50089 32243 -50055 32277
rect -50017 32243 -49983 32277
rect -49945 32243 -49911 32277
rect -49873 32243 -49839 32277
rect -49801 32243 -49767 32277
rect -49729 32243 -49695 32277
rect -49657 32243 -49623 32277
rect -49585 32243 -49551 32277
rect -49513 32243 -49479 32277
rect -49441 32243 -49407 32277
rect -49369 32243 -49335 32277
rect -49297 32243 -49263 32277
rect -49225 32243 -49191 32277
rect -49153 32243 -49119 32277
rect -49081 32243 -49047 32277
rect -49009 32243 -48975 32277
rect -48937 32243 -48903 32277
rect -48865 32243 -48831 32277
rect 2898 32315 2932 32349
rect 2970 32315 3004 32349
rect 3042 32315 3076 32349
rect 3114 32315 3148 32349
rect 3186 32315 3220 32349
rect 3258 32315 3292 32349
rect 3330 32315 3364 32349
rect 3402 32315 3436 32349
rect 3474 32315 3508 32349
rect 3546 32315 3580 32349
rect 3618 32315 3652 32349
rect 3690 32315 3724 32349
rect 3762 32315 3796 32349
rect 3834 32315 3868 32349
rect 3906 32315 3940 32349
rect 3978 32315 4012 32349
rect 4050 32315 4084 32349
rect 4122 32315 4156 32349
rect 4194 32315 4228 32349
rect 4266 32315 4300 32349
rect 4338 32315 4372 32349
rect 4410 32315 4444 32349
rect 4482 32315 4516 32349
rect 2898 32243 2932 32277
rect 2970 32243 3004 32277
rect 3042 32243 3076 32277
rect 3114 32243 3148 32277
rect 3186 32243 3220 32277
rect 3258 32243 3292 32277
rect 3330 32243 3364 32277
rect 3402 32243 3436 32277
rect 3474 32243 3508 32277
rect 3546 32243 3580 32277
rect 3618 32243 3652 32277
rect 3690 32243 3724 32277
rect 3762 32243 3796 32277
rect 3834 32243 3868 32277
rect 3906 32243 3940 32277
rect 3978 32243 4012 32277
rect 4050 32243 4084 32277
rect 4122 32243 4156 32277
rect 4194 32243 4228 32277
rect 4266 32243 4300 32277
rect 4338 32243 4372 32277
rect 4410 32243 4444 32277
rect 4482 32243 4516 32277
rect -50803 32131 -50769 32165
rect -50735 32131 -50701 32165
rect -50899 32035 -50865 32069
rect -50899 31967 -50865 32001
rect -50639 32035 -50605 32069
rect -50639 31967 -50605 32001
rect -50803 31871 -50769 31905
rect -50735 31871 -50701 31905
<< nsubdiffcont >>
rect -50449 33490 -50415 33524
rect -50377 33490 -50343 33524
rect -50305 33490 -50271 33524
rect -50233 33490 -50199 33524
rect -50161 33490 -50127 33524
rect -50089 33490 -50055 33524
rect -50017 33490 -49983 33524
rect -49945 33490 -49911 33524
rect -49873 33490 -49839 33524
rect -49801 33490 -49767 33524
rect -49729 33490 -49695 33524
rect -49657 33490 -49623 33524
rect -49585 33490 -49551 33524
rect -49513 33490 -49479 33524
rect -49441 33490 -49407 33524
rect -49369 33490 -49335 33524
rect -49297 33490 -49263 33524
rect -49225 33490 -49191 33524
rect -49153 33490 -49119 33524
rect -49081 33490 -49047 33524
rect -49009 33490 -48975 33524
rect -48937 33490 -48903 33524
rect -48865 33490 -48831 33524
rect -50449 33418 -50415 33452
rect -50377 33418 -50343 33452
rect -50305 33418 -50271 33452
rect -50233 33418 -50199 33452
rect -50161 33418 -50127 33452
rect -50089 33418 -50055 33452
rect -50017 33418 -49983 33452
rect -49945 33418 -49911 33452
rect -49873 33418 -49839 33452
rect -49801 33418 -49767 33452
rect -49729 33418 -49695 33452
rect -49657 33418 -49623 33452
rect -49585 33418 -49551 33452
rect -49513 33418 -49479 33452
rect -49441 33418 -49407 33452
rect -49369 33418 -49335 33452
rect -49297 33418 -49263 33452
rect -49225 33418 -49191 33452
rect -49153 33418 -49119 33452
rect -49081 33418 -49047 33452
rect -49009 33418 -48975 33452
rect -48937 33418 -48903 33452
rect -48865 33418 -48831 33452
rect 2898 33490 2932 33524
rect 2970 33490 3004 33524
rect 3042 33490 3076 33524
rect 3114 33490 3148 33524
rect 3186 33490 3220 33524
rect 3258 33490 3292 33524
rect 3330 33490 3364 33524
rect 3402 33490 3436 33524
rect 3474 33490 3508 33524
rect 3546 33490 3580 33524
rect 3618 33490 3652 33524
rect 3690 33490 3724 33524
rect 3762 33490 3796 33524
rect 3834 33490 3868 33524
rect 3906 33490 3940 33524
rect 3978 33490 4012 33524
rect 4050 33490 4084 33524
rect 4122 33490 4156 33524
rect 4194 33490 4228 33524
rect 4266 33490 4300 33524
rect 4338 33490 4372 33524
rect 4410 33490 4444 33524
rect 4482 33490 4516 33524
rect 2898 33418 2932 33452
rect 2970 33418 3004 33452
rect 3042 33418 3076 33452
rect 3114 33418 3148 33452
rect 3186 33418 3220 33452
rect 3258 33418 3292 33452
rect 3330 33418 3364 33452
rect 3402 33418 3436 33452
rect 3474 33418 3508 33452
rect 3546 33418 3580 33452
rect 3618 33418 3652 33452
rect 3690 33418 3724 33452
rect 3762 33418 3796 33452
rect 3834 33418 3868 33452
rect 3906 33418 3940 33452
rect 3978 33418 4012 33452
rect 4050 33418 4084 33452
rect 4122 33418 4156 33452
rect 4194 33418 4228 33452
rect 4266 33418 4300 33452
rect 4338 33418 4372 33452
rect 4410 33418 4444 33452
rect 4482 33418 4516 33452
<< poly >>
rect -50401 33312 -50301 33338
rect -50243 33312 -50143 33338
rect -50085 33312 -49985 33338
rect -49927 33312 -49827 33338
rect -49769 33312 -49669 33338
rect -49611 33312 -49511 33338
rect -49453 33312 -49353 33338
rect -49295 33312 -49195 33338
rect -49137 33312 -49037 33338
rect -48979 33312 -48879 33338
rect 2946 33312 3046 33338
rect 3104 33312 3204 33338
rect 3262 33312 3362 33338
rect 3420 33312 3520 33338
rect 3578 33312 3678 33338
rect 3736 33312 3836 33338
rect 3894 33312 3994 33338
rect 4052 33312 4152 33338
rect 4210 33312 4310 33338
rect 4368 33312 4468 33338
rect -50401 32865 -50301 32912
rect -50401 32831 -50368 32865
rect -50334 32831 -50301 32865
rect -50401 32815 -50301 32831
rect -50243 32865 -50143 32912
rect -50243 32831 -50210 32865
rect -50176 32831 -50143 32865
rect -50243 32815 -50143 32831
rect -50085 32865 -49985 32912
rect -50085 32831 -50052 32865
rect -50018 32831 -49985 32865
rect -50085 32815 -49985 32831
rect -49927 32865 -49827 32912
rect -49927 32831 -49894 32865
rect -49860 32831 -49827 32865
rect -49927 32815 -49827 32831
rect -49769 32865 -49669 32912
rect -49769 32831 -49736 32865
rect -49702 32831 -49669 32865
rect -49769 32815 -49669 32831
rect -49611 32865 -49511 32912
rect -49611 32831 -49578 32865
rect -49544 32831 -49511 32865
rect -49611 32815 -49511 32831
rect -49453 32865 -49353 32912
rect -49453 32831 -49420 32865
rect -49386 32831 -49353 32865
rect -49453 32815 -49353 32831
rect -49295 32865 -49195 32912
rect -49295 32831 -49262 32865
rect -49228 32831 -49195 32865
rect -49295 32815 -49195 32831
rect -49137 32865 -49037 32912
rect -49137 32831 -49104 32865
rect -49070 32831 -49037 32865
rect -49137 32815 -49037 32831
rect -48979 32865 -48879 32912
rect -48979 32831 -48946 32865
rect -48912 32831 -48879 32865
rect -48979 32815 -48879 32831
rect 2946 32865 3046 32912
rect 2946 32831 2979 32865
rect 3013 32831 3046 32865
rect 2946 32815 3046 32831
rect 3104 32865 3204 32912
rect 3104 32831 3137 32865
rect 3171 32831 3204 32865
rect 3104 32815 3204 32831
rect 3262 32865 3362 32912
rect 3262 32831 3295 32865
rect 3329 32831 3362 32865
rect 3262 32815 3362 32831
rect 3420 32865 3520 32912
rect 3420 32831 3453 32865
rect 3487 32831 3520 32865
rect 3420 32815 3520 32831
rect 3578 32865 3678 32912
rect 3578 32831 3611 32865
rect 3645 32831 3678 32865
rect 3578 32815 3678 32831
rect 3736 32865 3836 32912
rect 3736 32831 3769 32865
rect 3803 32831 3836 32865
rect 3736 32815 3836 32831
rect 3894 32865 3994 32912
rect 3894 32831 3927 32865
rect 3961 32831 3994 32865
rect 3894 32815 3994 32831
rect 4052 32865 4152 32912
rect 4052 32831 4085 32865
rect 4119 32831 4152 32865
rect 4052 32815 4152 32831
rect 4210 32865 4310 32912
rect 4210 32831 4243 32865
rect 4277 32831 4310 32865
rect 4210 32815 4310 32831
rect 4368 32865 4468 32912
rect 4368 32831 4401 32865
rect 4435 32831 4468 32865
rect 4368 32815 4468 32831
rect -50401 32727 -50301 32743
rect -50401 32693 -50368 32727
rect -50334 32693 -50301 32727
rect -50401 32655 -50301 32693
rect -50243 32727 -50143 32743
rect -50243 32693 -50210 32727
rect -50176 32693 -50143 32727
rect -50243 32655 -50143 32693
rect -50085 32727 -49985 32743
rect -50085 32693 -50052 32727
rect -50018 32693 -49985 32727
rect -50085 32655 -49985 32693
rect -49927 32727 -49827 32743
rect -49927 32693 -49894 32727
rect -49860 32693 -49827 32727
rect -49927 32655 -49827 32693
rect -49769 32727 -49669 32743
rect -49769 32693 -49736 32727
rect -49702 32693 -49669 32727
rect -49769 32655 -49669 32693
rect -49611 32727 -49511 32743
rect -49611 32693 -49578 32727
rect -49544 32693 -49511 32727
rect -49611 32655 -49511 32693
rect -49453 32727 -49353 32743
rect -49453 32693 -49420 32727
rect -49386 32693 -49353 32727
rect -49453 32655 -49353 32693
rect -49295 32727 -49195 32743
rect -49295 32693 -49262 32727
rect -49228 32693 -49195 32727
rect -49295 32655 -49195 32693
rect -49137 32727 -49037 32743
rect -49137 32693 -49104 32727
rect -49070 32693 -49037 32727
rect -49137 32655 -49037 32693
rect -48979 32727 -48879 32743
rect -48979 32693 -48946 32727
rect -48912 32693 -48879 32727
rect -48979 32655 -48879 32693
rect 2946 32727 3046 32743
rect 2946 32693 2979 32727
rect 3013 32693 3046 32727
rect 2946 32655 3046 32693
rect 3104 32727 3204 32743
rect 3104 32693 3137 32727
rect 3171 32693 3204 32727
rect 3104 32655 3204 32693
rect 3262 32727 3362 32743
rect 3262 32693 3295 32727
rect 3329 32693 3362 32727
rect 3262 32655 3362 32693
rect 3420 32727 3520 32743
rect 3420 32693 3453 32727
rect 3487 32693 3520 32727
rect 3420 32655 3520 32693
rect 3578 32727 3678 32743
rect 3578 32693 3611 32727
rect 3645 32693 3678 32727
rect 3578 32655 3678 32693
rect 3736 32727 3836 32743
rect 3736 32693 3769 32727
rect 3803 32693 3836 32727
rect 3736 32655 3836 32693
rect 3894 32727 3994 32743
rect 3894 32693 3927 32727
rect 3961 32693 3994 32727
rect 3894 32655 3994 32693
rect 4052 32727 4152 32743
rect 4052 32693 4085 32727
rect 4119 32693 4152 32727
rect 4052 32655 4152 32693
rect 4210 32727 4310 32743
rect 4210 32693 4243 32727
rect 4277 32693 4310 32727
rect 4210 32655 4310 32693
rect 4368 32727 4468 32743
rect 4368 32693 4401 32727
rect 4435 32693 4468 32727
rect 4368 32655 4468 32693
rect -50401 32429 -50301 32455
rect -50243 32429 -50143 32455
rect -50085 32429 -49985 32455
rect -49927 32429 -49827 32455
rect -49769 32429 -49669 32455
rect -49611 32429 -49511 32455
rect -49453 32429 -49353 32455
rect -49295 32429 -49195 32455
rect -49137 32429 -49037 32455
rect -48979 32429 -48879 32455
rect 2946 32429 3046 32455
rect 3104 32429 3204 32455
rect 3262 32429 3362 32455
rect 3420 32429 3520 32455
rect 3578 32429 3678 32455
rect 3736 32429 3836 32455
rect 3894 32429 3994 32455
rect 4052 32429 4152 32455
rect 4210 32429 4310 32455
rect 4368 32429 4468 32455
rect -42474 5437 -42444 5463
rect -42378 5437 -42348 5463
rect -42282 5437 -42252 5463
rect -42186 5437 -42156 5463
rect -42090 5437 -42060 5463
rect -41994 5437 -41964 5463
rect -41898 5437 -41868 5463
rect -41802 5437 -41772 5463
rect -41706 5437 -41676 5463
rect -41610 5437 -41580 5463
rect -41514 5437 -41484 5463
rect -41418 5437 -41388 5463
rect -41322 5437 -41292 5463
rect -41226 5437 -41196 5463
rect -41130 5437 -41100 5463
rect -41034 5437 -41004 5463
rect -40938 5437 -40908 5463
rect -40842 5437 -40812 5463
rect -40746 5437 -40716 5463
rect 154 5425 184 5451
rect 250 5425 280 5451
rect 346 5425 376 5451
rect 442 5425 472 5451
rect 538 5425 568 5451
rect 634 5425 664 5451
rect 730 5425 760 5451
rect 826 5425 856 5451
rect 922 5425 952 5451
rect 1018 5425 1048 5451
rect 1114 5425 1144 5451
rect 1210 5425 1240 5451
rect 1306 5425 1336 5451
rect 1402 5425 1432 5451
rect 1498 5425 1528 5451
rect 1594 5425 1624 5451
rect 1690 5425 1720 5451
rect 1786 5425 1816 5451
rect 1882 5425 1912 5451
rect -42474 4607 -42444 4637
rect -42378 4607 -42348 4637
rect -42282 4607 -42252 4637
rect -42186 4607 -42156 4637
rect -42090 4607 -42060 4637
rect -41994 4607 -41964 4637
rect -41898 4607 -41868 4637
rect -41802 4607 -41772 4637
rect -41706 4607 -41676 4637
rect -41610 4607 -41580 4637
rect -41514 4607 -41484 4637
rect -41418 4607 -41388 4637
rect -41322 4607 -41292 4637
rect -41226 4607 -41196 4637
rect -41130 4607 -41100 4637
rect -41034 4607 -41004 4637
rect -40938 4607 -40908 4637
rect -40842 4607 -40812 4637
rect -40746 4607 -40716 4637
rect -42474 4567 -40716 4607
rect -42474 4533 -42440 4567
rect -42406 4533 -42368 4567
rect -42334 4533 -42296 4567
rect -42262 4533 -42224 4567
rect -42190 4533 -42152 4567
rect -42118 4533 -42080 4567
rect -42046 4533 -42008 4567
rect -41974 4533 -41936 4567
rect -41902 4533 -41864 4567
rect -41830 4533 -41792 4567
rect -41758 4533 -41720 4567
rect -41686 4533 -41648 4567
rect -41614 4533 -41576 4567
rect -41542 4533 -41504 4567
rect -41470 4533 -41432 4567
rect -41398 4533 -41360 4567
rect -41326 4533 -41288 4567
rect -41254 4533 -41216 4567
rect -41182 4533 -41144 4567
rect -41110 4533 -41072 4567
rect -41038 4533 -41000 4567
rect -40966 4533 -40928 4567
rect -40894 4533 -40856 4567
rect -40822 4533 -40784 4567
rect -40750 4533 -40716 4567
rect -42474 4495 -40716 4533
rect -42474 4461 -42440 4495
rect -42406 4461 -42368 4495
rect -42334 4461 -42296 4495
rect -42262 4461 -42224 4495
rect -42190 4461 -42152 4495
rect -42118 4461 -42080 4495
rect -42046 4461 -42008 4495
rect -41974 4461 -41936 4495
rect -41902 4461 -41864 4495
rect -41830 4461 -41792 4495
rect -41758 4461 -41720 4495
rect -41686 4461 -41648 4495
rect -41614 4461 -41576 4495
rect -41542 4461 -41504 4495
rect -41470 4461 -41432 4495
rect -41398 4461 -41360 4495
rect -41326 4461 -41288 4495
rect -41254 4461 -41216 4495
rect -41182 4461 -41144 4495
rect -41110 4461 -41072 4495
rect -41038 4461 -41000 4495
rect -40966 4461 -40928 4495
rect -40894 4461 -40856 4495
rect -40822 4461 -40784 4495
rect -40750 4461 -40716 4495
rect -42474 4451 -40716 4461
rect 154 4600 184 4625
rect 250 4600 280 4625
rect 346 4600 376 4625
rect 442 4600 472 4625
rect 538 4600 568 4625
rect 634 4600 664 4625
rect 730 4600 760 4625
rect 826 4600 856 4625
rect 922 4600 952 4625
rect 1018 4600 1048 4625
rect 1114 4600 1144 4625
rect 1210 4600 1240 4625
rect 1306 4600 1336 4625
rect 1402 4600 1432 4625
rect 1498 4600 1528 4625
rect 1594 4600 1624 4625
rect 1690 4600 1720 4625
rect 1786 4600 1816 4625
rect 1882 4600 1912 4625
rect 154 4560 1912 4600
rect 154 4526 188 4560
rect 222 4526 260 4560
rect 294 4526 332 4560
rect 366 4526 404 4560
rect 438 4526 476 4560
rect 510 4526 548 4560
rect 582 4526 620 4560
rect 654 4526 692 4560
rect 726 4526 764 4560
rect 798 4526 836 4560
rect 870 4526 908 4560
rect 942 4526 980 4560
rect 1014 4526 1052 4560
rect 1086 4526 1124 4560
rect 1158 4526 1196 4560
rect 1230 4526 1268 4560
rect 1302 4526 1340 4560
rect 1374 4526 1412 4560
rect 1446 4526 1484 4560
rect 1518 4526 1556 4560
rect 1590 4526 1628 4560
rect 1662 4526 1700 4560
rect 1734 4526 1772 4560
rect 1806 4526 1844 4560
rect 1878 4526 1912 4560
rect 154 4488 1912 4526
rect 154 4454 188 4488
rect 222 4454 260 4488
rect 294 4454 332 4488
rect 366 4454 404 4488
rect 438 4454 476 4488
rect 510 4454 548 4488
rect 582 4454 620 4488
rect 654 4454 692 4488
rect 726 4454 764 4488
rect 798 4454 836 4488
rect 870 4454 908 4488
rect 942 4454 980 4488
rect 1014 4454 1052 4488
rect 1086 4454 1124 4488
rect 1158 4454 1196 4488
rect 1230 4454 1268 4488
rect 1302 4454 1340 4488
rect 1374 4454 1412 4488
rect 1446 4454 1484 4488
rect 1518 4454 1556 4488
rect 1590 4454 1628 4488
rect 1662 4454 1700 4488
rect 1734 4454 1772 4488
rect 1806 4454 1844 4488
rect 1878 4454 1912 4488
rect 154 4444 1912 4454
rect -42475 -4737 -42445 -4711
rect -42379 -4737 -42349 -4711
rect -42283 -4737 -42253 -4711
rect -42187 -4737 -42157 -4711
rect -42091 -4737 -42061 -4711
rect -41995 -4737 -41965 -4711
rect -41899 -4737 -41869 -4711
rect -41803 -4737 -41773 -4711
rect -41707 -4737 -41677 -4711
rect -41611 -4737 -41581 -4711
rect -41515 -4737 -41485 -4711
rect -41419 -4737 -41389 -4711
rect -41323 -4737 -41293 -4711
rect -41227 -4737 -41197 -4711
rect -41131 -4737 -41101 -4711
rect -41035 -4737 -41005 -4711
rect -40939 -4737 -40909 -4711
rect -40843 -4737 -40813 -4711
rect -40747 -4737 -40717 -4711
rect 166 -4763 196 -4737
rect 262 -4763 292 -4737
rect 358 -4763 388 -4737
rect 454 -4763 484 -4737
rect 550 -4763 580 -4737
rect 646 -4763 676 -4737
rect 742 -4763 772 -4737
rect 838 -4763 868 -4737
rect 934 -4763 964 -4737
rect 1030 -4763 1060 -4737
rect 1126 -4763 1156 -4737
rect 1222 -4763 1252 -4737
rect 1318 -4763 1348 -4737
rect 1414 -4763 1444 -4737
rect 1510 -4763 1540 -4737
rect 1606 -4763 1636 -4737
rect 1702 -4763 1732 -4737
rect 1798 -4763 1828 -4737
rect 1894 -4763 1924 -4737
rect -42475 -5567 -42445 -5537
rect -42379 -5567 -42349 -5537
rect -42283 -5567 -42253 -5537
rect -42187 -5567 -42157 -5537
rect -42091 -5567 -42061 -5537
rect -41995 -5567 -41965 -5537
rect -41899 -5567 -41869 -5537
rect -41803 -5567 -41773 -5537
rect -41707 -5567 -41677 -5537
rect -41611 -5567 -41581 -5537
rect -41515 -5567 -41485 -5537
rect -41419 -5567 -41389 -5537
rect -41323 -5567 -41293 -5537
rect -41227 -5567 -41197 -5537
rect -41131 -5567 -41101 -5537
rect -41035 -5567 -41005 -5537
rect -40939 -5567 -40909 -5537
rect -40843 -5567 -40813 -5537
rect -40747 -5567 -40717 -5537
rect -42475 -5607 -40717 -5567
rect -42475 -5641 -42441 -5607
rect -42407 -5641 -42369 -5607
rect -42335 -5641 -42297 -5607
rect -42263 -5641 -42225 -5607
rect -42191 -5641 -42153 -5607
rect -42119 -5641 -42081 -5607
rect -42047 -5641 -42009 -5607
rect -41975 -5641 -41937 -5607
rect -41903 -5641 -41865 -5607
rect -41831 -5641 -41793 -5607
rect -41759 -5641 -41721 -5607
rect -41687 -5641 -41649 -5607
rect -41615 -5641 -41577 -5607
rect -41543 -5641 -41505 -5607
rect -41471 -5641 -41433 -5607
rect -41399 -5641 -41361 -5607
rect -41327 -5641 -41289 -5607
rect -41255 -5641 -41217 -5607
rect -41183 -5641 -41145 -5607
rect -41111 -5641 -41073 -5607
rect -41039 -5641 -41001 -5607
rect -40967 -5641 -40929 -5607
rect -40895 -5641 -40857 -5607
rect -40823 -5641 -40785 -5607
rect -40751 -5641 -40717 -5607
rect -42475 -5679 -40717 -5641
rect -42475 -5713 -42441 -5679
rect -42407 -5713 -42369 -5679
rect -42335 -5713 -42297 -5679
rect -42263 -5713 -42225 -5679
rect -42191 -5713 -42153 -5679
rect -42119 -5713 -42081 -5679
rect -42047 -5713 -42009 -5679
rect -41975 -5713 -41937 -5679
rect -41903 -5713 -41865 -5679
rect -41831 -5713 -41793 -5679
rect -41759 -5713 -41721 -5679
rect -41687 -5713 -41649 -5679
rect -41615 -5713 -41577 -5679
rect -41543 -5713 -41505 -5679
rect -41471 -5713 -41433 -5679
rect -41399 -5713 -41361 -5679
rect -41327 -5713 -41289 -5679
rect -41255 -5713 -41217 -5679
rect -41183 -5713 -41145 -5679
rect -41111 -5713 -41073 -5679
rect -41039 -5713 -41001 -5679
rect -40967 -5713 -40929 -5679
rect -40895 -5713 -40857 -5679
rect -40823 -5713 -40785 -5679
rect -40751 -5713 -40717 -5679
rect -42475 -5723 -40717 -5713
rect 166 -5593 196 -5563
rect 262 -5593 292 -5563
rect 358 -5593 388 -5563
rect 454 -5593 484 -5563
rect 550 -5593 580 -5563
rect 646 -5593 676 -5563
rect 742 -5593 772 -5563
rect 838 -5593 868 -5563
rect 934 -5593 964 -5563
rect 1030 -5593 1060 -5563
rect 1126 -5593 1156 -5563
rect 1222 -5593 1252 -5563
rect 1318 -5593 1348 -5563
rect 1414 -5593 1444 -5563
rect 1510 -5593 1540 -5563
rect 1606 -5593 1636 -5563
rect 1702 -5593 1732 -5563
rect 1798 -5593 1828 -5563
rect 1894 -5593 1924 -5563
rect 166 -5633 1924 -5593
rect 166 -5667 200 -5633
rect 234 -5667 272 -5633
rect 306 -5667 344 -5633
rect 378 -5667 416 -5633
rect 450 -5667 488 -5633
rect 522 -5667 560 -5633
rect 594 -5667 632 -5633
rect 666 -5667 704 -5633
rect 738 -5667 776 -5633
rect 810 -5667 848 -5633
rect 882 -5667 920 -5633
rect 954 -5667 992 -5633
rect 1026 -5667 1064 -5633
rect 1098 -5667 1136 -5633
rect 1170 -5667 1208 -5633
rect 1242 -5667 1280 -5633
rect 1314 -5667 1352 -5633
rect 1386 -5667 1424 -5633
rect 1458 -5667 1496 -5633
rect 1530 -5667 1568 -5633
rect 1602 -5667 1640 -5633
rect 1674 -5667 1712 -5633
rect 1746 -5667 1784 -5633
rect 1818 -5667 1856 -5633
rect 1890 -5667 1924 -5633
rect 166 -5705 1924 -5667
rect 166 -5739 200 -5705
rect 234 -5739 272 -5705
rect 306 -5739 344 -5705
rect 378 -5739 416 -5705
rect 450 -5739 488 -5705
rect 522 -5739 560 -5705
rect 594 -5739 632 -5705
rect 666 -5739 704 -5705
rect 738 -5739 776 -5705
rect 810 -5739 848 -5705
rect 882 -5739 920 -5705
rect 954 -5739 992 -5705
rect 1026 -5739 1064 -5705
rect 1098 -5739 1136 -5705
rect 1170 -5739 1208 -5705
rect 1242 -5739 1280 -5705
rect 1314 -5739 1352 -5705
rect 1386 -5739 1424 -5705
rect 1458 -5739 1496 -5705
rect 1530 -5739 1568 -5705
rect 1602 -5739 1640 -5705
rect 1674 -5739 1712 -5705
rect 1746 -5739 1784 -5705
rect 1818 -5739 1856 -5705
rect 1890 -5739 1924 -5705
rect 166 -5749 1924 -5739
<< polycont >>
rect -50368 32831 -50334 32865
rect -50210 32831 -50176 32865
rect -50052 32831 -50018 32865
rect -49894 32831 -49860 32865
rect -49736 32831 -49702 32865
rect -49578 32831 -49544 32865
rect -49420 32831 -49386 32865
rect -49262 32831 -49228 32865
rect -49104 32831 -49070 32865
rect -48946 32831 -48912 32865
rect 2979 32831 3013 32865
rect 3137 32831 3171 32865
rect 3295 32831 3329 32865
rect 3453 32831 3487 32865
rect 3611 32831 3645 32865
rect 3769 32831 3803 32865
rect 3927 32831 3961 32865
rect 4085 32831 4119 32865
rect 4243 32831 4277 32865
rect 4401 32831 4435 32865
rect -50368 32693 -50334 32727
rect -50210 32693 -50176 32727
rect -50052 32693 -50018 32727
rect -49894 32693 -49860 32727
rect -49736 32693 -49702 32727
rect -49578 32693 -49544 32727
rect -49420 32693 -49386 32727
rect -49262 32693 -49228 32727
rect -49104 32693 -49070 32727
rect -48946 32693 -48912 32727
rect 2979 32693 3013 32727
rect 3137 32693 3171 32727
rect 3295 32693 3329 32727
rect 3453 32693 3487 32727
rect 3611 32693 3645 32727
rect 3769 32693 3803 32727
rect 3927 32693 3961 32727
rect 4085 32693 4119 32727
rect 4243 32693 4277 32727
rect 4401 32693 4435 32727
rect -42440 4533 -42406 4567
rect -42368 4533 -42334 4567
rect -42296 4533 -42262 4567
rect -42224 4533 -42190 4567
rect -42152 4533 -42118 4567
rect -42080 4533 -42046 4567
rect -42008 4533 -41974 4567
rect -41936 4533 -41902 4567
rect -41864 4533 -41830 4567
rect -41792 4533 -41758 4567
rect -41720 4533 -41686 4567
rect -41648 4533 -41614 4567
rect -41576 4533 -41542 4567
rect -41504 4533 -41470 4567
rect -41432 4533 -41398 4567
rect -41360 4533 -41326 4567
rect -41288 4533 -41254 4567
rect -41216 4533 -41182 4567
rect -41144 4533 -41110 4567
rect -41072 4533 -41038 4567
rect -41000 4533 -40966 4567
rect -40928 4533 -40894 4567
rect -40856 4533 -40822 4567
rect -40784 4533 -40750 4567
rect -42440 4461 -42406 4495
rect -42368 4461 -42334 4495
rect -42296 4461 -42262 4495
rect -42224 4461 -42190 4495
rect -42152 4461 -42118 4495
rect -42080 4461 -42046 4495
rect -42008 4461 -41974 4495
rect -41936 4461 -41902 4495
rect -41864 4461 -41830 4495
rect -41792 4461 -41758 4495
rect -41720 4461 -41686 4495
rect -41648 4461 -41614 4495
rect -41576 4461 -41542 4495
rect -41504 4461 -41470 4495
rect -41432 4461 -41398 4495
rect -41360 4461 -41326 4495
rect -41288 4461 -41254 4495
rect -41216 4461 -41182 4495
rect -41144 4461 -41110 4495
rect -41072 4461 -41038 4495
rect -41000 4461 -40966 4495
rect -40928 4461 -40894 4495
rect -40856 4461 -40822 4495
rect -40784 4461 -40750 4495
rect 188 4526 222 4560
rect 260 4526 294 4560
rect 332 4526 366 4560
rect 404 4526 438 4560
rect 476 4526 510 4560
rect 548 4526 582 4560
rect 620 4526 654 4560
rect 692 4526 726 4560
rect 764 4526 798 4560
rect 836 4526 870 4560
rect 908 4526 942 4560
rect 980 4526 1014 4560
rect 1052 4526 1086 4560
rect 1124 4526 1158 4560
rect 1196 4526 1230 4560
rect 1268 4526 1302 4560
rect 1340 4526 1374 4560
rect 1412 4526 1446 4560
rect 1484 4526 1518 4560
rect 1556 4526 1590 4560
rect 1628 4526 1662 4560
rect 1700 4526 1734 4560
rect 1772 4526 1806 4560
rect 1844 4526 1878 4560
rect 188 4454 222 4488
rect 260 4454 294 4488
rect 332 4454 366 4488
rect 404 4454 438 4488
rect 476 4454 510 4488
rect 548 4454 582 4488
rect 620 4454 654 4488
rect 692 4454 726 4488
rect 764 4454 798 4488
rect 836 4454 870 4488
rect 908 4454 942 4488
rect 980 4454 1014 4488
rect 1052 4454 1086 4488
rect 1124 4454 1158 4488
rect 1196 4454 1230 4488
rect 1268 4454 1302 4488
rect 1340 4454 1374 4488
rect 1412 4454 1446 4488
rect 1484 4454 1518 4488
rect 1556 4454 1590 4488
rect 1628 4454 1662 4488
rect 1700 4454 1734 4488
rect 1772 4454 1806 4488
rect 1844 4454 1878 4488
rect -42441 -5641 -42407 -5607
rect -42369 -5641 -42335 -5607
rect -42297 -5641 -42263 -5607
rect -42225 -5641 -42191 -5607
rect -42153 -5641 -42119 -5607
rect -42081 -5641 -42047 -5607
rect -42009 -5641 -41975 -5607
rect -41937 -5641 -41903 -5607
rect -41865 -5641 -41831 -5607
rect -41793 -5641 -41759 -5607
rect -41721 -5641 -41687 -5607
rect -41649 -5641 -41615 -5607
rect -41577 -5641 -41543 -5607
rect -41505 -5641 -41471 -5607
rect -41433 -5641 -41399 -5607
rect -41361 -5641 -41327 -5607
rect -41289 -5641 -41255 -5607
rect -41217 -5641 -41183 -5607
rect -41145 -5641 -41111 -5607
rect -41073 -5641 -41039 -5607
rect -41001 -5641 -40967 -5607
rect -40929 -5641 -40895 -5607
rect -40857 -5641 -40823 -5607
rect -40785 -5641 -40751 -5607
rect -42441 -5713 -42407 -5679
rect -42369 -5713 -42335 -5679
rect -42297 -5713 -42263 -5679
rect -42225 -5713 -42191 -5679
rect -42153 -5713 -42119 -5679
rect -42081 -5713 -42047 -5679
rect -42009 -5713 -41975 -5679
rect -41937 -5713 -41903 -5679
rect -41865 -5713 -41831 -5679
rect -41793 -5713 -41759 -5679
rect -41721 -5713 -41687 -5679
rect -41649 -5713 -41615 -5679
rect -41577 -5713 -41543 -5679
rect -41505 -5713 -41471 -5679
rect -41433 -5713 -41399 -5679
rect -41361 -5713 -41327 -5679
rect -41289 -5713 -41255 -5679
rect -41217 -5713 -41183 -5679
rect -41145 -5713 -41111 -5679
rect -41073 -5713 -41039 -5679
rect -41001 -5713 -40967 -5679
rect -40929 -5713 -40895 -5679
rect -40857 -5713 -40823 -5679
rect -40785 -5713 -40751 -5679
rect 200 -5667 234 -5633
rect 272 -5667 306 -5633
rect 344 -5667 378 -5633
rect 416 -5667 450 -5633
rect 488 -5667 522 -5633
rect 560 -5667 594 -5633
rect 632 -5667 666 -5633
rect 704 -5667 738 -5633
rect 776 -5667 810 -5633
rect 848 -5667 882 -5633
rect 920 -5667 954 -5633
rect 992 -5667 1026 -5633
rect 1064 -5667 1098 -5633
rect 1136 -5667 1170 -5633
rect 1208 -5667 1242 -5633
rect 1280 -5667 1314 -5633
rect 1352 -5667 1386 -5633
rect 1424 -5667 1458 -5633
rect 1496 -5667 1530 -5633
rect 1568 -5667 1602 -5633
rect 1640 -5667 1674 -5633
rect 1712 -5667 1746 -5633
rect 1784 -5667 1818 -5633
rect 1856 -5667 1890 -5633
rect 200 -5739 234 -5705
rect 272 -5739 306 -5705
rect 344 -5739 378 -5705
rect 416 -5739 450 -5705
rect 488 -5739 522 -5705
rect 560 -5739 594 -5705
rect 632 -5739 666 -5705
rect 704 -5739 738 -5705
rect 776 -5739 810 -5705
rect 848 -5739 882 -5705
rect 920 -5739 954 -5705
rect 992 -5739 1026 -5705
rect 1064 -5739 1098 -5705
rect 1136 -5739 1170 -5705
rect 1208 -5739 1242 -5705
rect 1280 -5739 1314 -5705
rect 1352 -5739 1386 -5705
rect 1424 -5739 1458 -5705
rect 1496 -5739 1530 -5705
rect 1568 -5739 1602 -5705
rect 1640 -5739 1674 -5705
rect 1712 -5739 1746 -5705
rect 1784 -5739 1818 -5705
rect 1856 -5739 1890 -5705
<< xpolycontact >>
rect -47356 24522 -47286 24954
rect -47356 15160 -47286 15522
rect -47038 24884 -46650 24954
rect -47038 24522 -46968 24884
rect -47038 15160 -46968 15522
rect -47356 15090 -46968 15160
rect -46720 24522 -46650 24884
rect -46720 15160 -46650 15522
rect -46402 24884 -46014 24954
rect -46402 24522 -46332 24884
rect -46402 15160 -46332 15522
rect -46720 15090 -46332 15160
rect -46084 24522 -46014 24884
rect -46084 15160 -46014 15522
rect -45766 24884 -45378 24954
rect -45766 24522 -45696 24884
rect -45766 15160 -45696 15522
rect -46084 15090 -45696 15160
rect -45448 24522 -45378 24884
rect -45448 15160 -45378 15522
rect -45130 24884 -44742 24954
rect -45130 24522 -45060 24884
rect -45130 15160 -45060 15522
rect -45448 15090 -45060 15160
rect -44812 24522 -44742 24884
rect -44812 15160 -44742 15522
rect -44494 24884 -44106 24954
rect -44494 24522 -44424 24884
rect -44494 15160 -44424 15522
rect -44812 15090 -44424 15160
rect -44176 24522 -44106 24884
rect -44176 15160 -44106 15522
rect -43858 24884 -43470 24954
rect -43858 24522 -43788 24884
rect -43858 15160 -43788 15522
rect -44176 15090 -43788 15160
rect -43540 24522 -43470 24884
rect -43540 15160 -43470 15522
rect -43222 24884 -42834 24954
rect -43222 24522 -43152 24884
rect -43222 15160 -43152 15522
rect -43540 15090 -43152 15160
rect -42904 24522 -42834 24884
rect -42904 15090 -42834 15522
rect 2404 24884 2792 24954
rect 2404 24522 2474 24884
rect 2404 15090 2474 15522
rect 2722 24522 2792 24884
rect 2722 15160 2792 15522
rect 3040 24884 3428 24954
rect 3040 24522 3110 24884
rect 3040 15160 3110 15522
rect 2722 15090 3110 15160
rect 3358 24522 3428 24884
rect 3358 15160 3428 15522
rect 3676 24884 4064 24954
rect 3676 24522 3746 24884
rect 3676 15160 3746 15522
rect 3358 15090 3746 15160
rect 3994 24522 4064 24884
rect 3994 15160 4064 15522
rect 4312 24884 4700 24954
rect 4312 24522 4382 24884
rect 4312 15160 4382 15522
rect 3994 15090 4382 15160
rect 4630 24522 4700 24884
rect 4630 15160 4700 15522
rect 4948 24884 5336 24954
rect 4948 24522 5018 24884
rect 4948 15160 5018 15522
rect 4630 15090 5018 15160
rect 5266 24522 5336 24884
rect 5266 15160 5336 15522
rect 5584 24884 5972 24954
rect 5584 24522 5654 24884
rect 5584 15160 5654 15522
rect 5266 15090 5654 15160
rect 5902 24522 5972 24884
rect 5902 15160 5972 15522
rect 6220 24884 6608 24954
rect 6220 24522 6290 24884
rect 6220 15160 6290 15522
rect 5902 15090 6290 15160
rect 6538 24522 6608 24884
rect 6538 15160 6608 15522
rect 6856 24522 6926 24954
rect 6856 15160 6926 15522
rect 6538 15090 6926 15160
rect -42904 4445 -42834 5003
rect 2404 4438 2474 4991
rect -42904 -5603 -42834 -5171
rect 2404 -5623 2474 -5191
<< xpolyres >>
rect -47356 15522 -47286 24522
rect -47038 15522 -46968 24522
rect -46720 15522 -46650 24522
rect -46402 15522 -46332 24522
rect -46084 15522 -46014 24522
rect -45766 15522 -45696 24522
rect -45448 15522 -45378 24522
rect -45130 15522 -45060 24522
rect -44812 15522 -44742 24522
rect -44494 15522 -44424 24522
rect -44176 15522 -44106 24522
rect -43858 15522 -43788 24522
rect -43540 15522 -43470 24522
rect -43222 15522 -43152 24522
rect -42904 15522 -42834 24522
rect -42904 5003 -42834 15090
rect 2404 15522 2474 24522
rect 2722 15522 2792 24522
rect 3040 15522 3110 24522
rect 3358 15522 3428 24522
rect 3676 15522 3746 24522
rect 3994 15522 4064 24522
rect 4312 15522 4382 24522
rect 4630 15522 4700 24522
rect 4948 15522 5018 24522
rect 5266 15522 5336 24522
rect 5584 15522 5654 24522
rect 5902 15522 5972 24522
rect 6220 15522 6290 24522
rect 6538 15522 6608 24522
rect 6856 15522 6926 24522
rect 2404 4991 2474 15090
rect -42904 -5171 -42834 4445
rect 2404 -5191 2474 4438
<< ndiode >>
rect 2125 32539 2215 32567
rect 2125 32505 2153 32539
rect 2187 32505 2215 32539
rect 2125 32477 2215 32505
rect -50797 32035 -50707 32063
rect -50797 32001 -50769 32035
rect -50735 32001 -50707 32035
rect -50797 31973 -50707 32001
<< ndiodec >>
rect 2153 32505 2187 32539
rect -50769 32001 -50735 32035
<< locali >>
rect -50465 33524 -48815 33540
rect -50465 33418 -50449 33524
rect -48831 33418 -48815 33524
rect -50465 33402 -48815 33418
rect 2882 33524 4532 33540
rect 2882 33418 2898 33524
rect 4516 33418 4532 33524
rect 2882 33402 4532 33418
rect -50447 33299 -50413 33316
rect -50447 33231 -50413 33239
rect -50447 33163 -50413 33167
rect -50447 33057 -50413 33061
rect -50447 32985 -50413 32993
rect -50942 32940 -50588 32956
rect -50942 32618 -50926 32940
rect -50604 32831 -50588 32940
rect -50447 32908 -50413 32925
rect -50289 33299 -50255 33316
rect -50289 33231 -50255 33239
rect -50289 33163 -50255 33167
rect -50289 33057 -50255 33061
rect -50289 32985 -50255 32993
rect -50289 32908 -50255 32925
rect -50131 33299 -50097 33316
rect -50131 33231 -50097 33239
rect -50131 33163 -50097 33167
rect -50131 33057 -50097 33061
rect -50131 32985 -50097 32993
rect -50131 32908 -50097 32925
rect -49973 33299 -49939 33316
rect -49973 33231 -49939 33239
rect -49973 33163 -49939 33167
rect -49973 33057 -49939 33061
rect -49973 32985 -49939 32993
rect -49973 32908 -49939 32925
rect -49815 33299 -49781 33316
rect -49815 33231 -49781 33239
rect -49815 33163 -49781 33167
rect -49815 33057 -49781 33061
rect -49815 32985 -49781 32993
rect -49815 32908 -49781 32925
rect -49657 33299 -49623 33316
rect -49657 33231 -49623 33239
rect -49657 33163 -49623 33167
rect -49657 33057 -49623 33061
rect -49657 32985 -49623 32993
rect -49657 32908 -49623 32925
rect -49499 33299 -49465 33316
rect -49499 33231 -49465 33239
rect -49499 33163 -49465 33167
rect -49499 33057 -49465 33061
rect -49499 32985 -49465 32993
rect -49499 32908 -49465 32925
rect -49341 33299 -49307 33316
rect -49341 33231 -49307 33239
rect -49341 33163 -49307 33167
rect -49341 33057 -49307 33061
rect -49341 32985 -49307 32993
rect -49341 32908 -49307 32925
rect -49183 33299 -49149 33316
rect -49183 33231 -49149 33239
rect -49183 33163 -49149 33167
rect -49183 33057 -49149 33061
rect -49183 32985 -49149 32993
rect -49183 32908 -49149 32925
rect -49025 33299 -48991 33316
rect -49025 33231 -48991 33239
rect -49025 33163 -48991 33167
rect -49025 33057 -48991 33061
rect -49025 32985 -48991 32993
rect -49025 32908 -48991 32925
rect -48867 33299 -48833 33316
rect -48867 33231 -48833 33239
rect -48867 33163 -48833 33167
rect -48867 33057 -48833 33061
rect -48867 32985 -48833 32993
rect 2900 33299 2934 33316
rect 2900 33231 2934 33239
rect 2900 33163 2934 33167
rect 2900 33057 2934 33061
rect 2900 32985 2934 32993
rect -48867 32908 -48833 32925
rect 2405 32940 2759 32956
rect -50401 32831 -50368 32865
rect -50334 32831 -50301 32865
rect -50243 32831 -50210 32865
rect -50176 32831 -50143 32865
rect -50085 32831 -50052 32865
rect -50018 32831 -49985 32865
rect -49927 32831 -49894 32865
rect -49860 32831 -49827 32865
rect -49769 32831 -49736 32865
rect -49702 32831 -49669 32865
rect -49611 32831 -49578 32865
rect -49544 32831 -49511 32865
rect -49453 32831 -49420 32865
rect -49386 32831 -49353 32865
rect -49295 32831 -49262 32865
rect -49228 32831 -49195 32865
rect -49137 32831 -49104 32865
rect -49070 32831 -49037 32865
rect -48979 32831 -48946 32865
rect -48912 32831 -48879 32865
rect -50604 32727 -48879 32831
rect -50604 32618 -50588 32727
rect -50401 32693 -50368 32727
rect -50334 32693 -50301 32727
rect -50243 32693 -50210 32727
rect -50176 32693 -50143 32727
rect -50085 32693 -50052 32727
rect -50018 32693 -49985 32727
rect -49927 32693 -49894 32727
rect -49860 32693 -49827 32727
rect -49769 32693 -49736 32727
rect -49702 32693 -49669 32727
rect -49611 32693 -49578 32727
rect -49544 32693 -49511 32727
rect -49453 32693 -49420 32727
rect -49386 32693 -49353 32727
rect -49295 32693 -49262 32727
rect -49228 32693 -49195 32727
rect -49137 32693 -49104 32727
rect -49070 32693 -49037 32727
rect -48979 32693 -48946 32727
rect -48912 32693 -48879 32727
rect -50942 32602 -50588 32618
rect -50447 32640 -50413 32659
rect -50447 32572 -50413 32574
rect -50447 32536 -50413 32538
rect -50447 32451 -50413 32470
rect -50289 32640 -50255 32659
rect -50289 32572 -50255 32574
rect -50289 32536 -50255 32538
rect -50289 32451 -50255 32470
rect -50131 32640 -50097 32659
rect -50131 32572 -50097 32574
rect -50131 32536 -50097 32538
rect -50131 32451 -50097 32470
rect -49973 32640 -49939 32659
rect -49973 32572 -49939 32574
rect -49973 32536 -49939 32538
rect -49973 32451 -49939 32470
rect -49815 32640 -49781 32659
rect -49815 32572 -49781 32574
rect -49815 32536 -49781 32538
rect -49815 32451 -49781 32470
rect -49657 32640 -49623 32659
rect -49657 32572 -49623 32574
rect -49657 32536 -49623 32538
rect -49657 32451 -49623 32470
rect -49499 32640 -49465 32659
rect -49499 32572 -49465 32574
rect -49499 32536 -49465 32538
rect -49499 32451 -49465 32470
rect -49341 32640 -49307 32659
rect -49341 32572 -49307 32574
rect -49341 32536 -49307 32538
rect -49341 32451 -49307 32470
rect -49183 32640 -49149 32659
rect -49183 32572 -49149 32574
rect -49183 32536 -49149 32538
rect -49183 32451 -49149 32470
rect -49025 32640 -48991 32659
rect -49025 32572 -48991 32574
rect -49025 32536 -48991 32538
rect -49025 32451 -48991 32470
rect -48867 32640 -48833 32659
rect -48867 32572 -48833 32574
rect -48867 32536 -48833 32538
rect -48867 32451 -48833 32470
rect 2023 32635 2119 32669
rect 2153 32635 2187 32669
rect 2221 32635 2317 32669
rect 2023 32573 2057 32635
rect 2283 32573 2317 32635
rect 2405 32618 2421 32940
rect 2743 32831 2759 32940
rect 2900 32908 2934 32925
rect 3058 33299 3092 33316
rect 3058 33231 3092 33239
rect 3058 33163 3092 33167
rect 3058 33057 3092 33061
rect 3058 32985 3092 32993
rect 3058 32908 3092 32925
rect 3216 33299 3250 33316
rect 3216 33231 3250 33239
rect 3216 33163 3250 33167
rect 3216 33057 3250 33061
rect 3216 32985 3250 32993
rect 3216 32908 3250 32925
rect 3374 33299 3408 33316
rect 3374 33231 3408 33239
rect 3374 33163 3408 33167
rect 3374 33057 3408 33061
rect 3374 32985 3408 32993
rect 3374 32908 3408 32925
rect 3532 33299 3566 33316
rect 3532 33231 3566 33239
rect 3532 33163 3566 33167
rect 3532 33057 3566 33061
rect 3532 32985 3566 32993
rect 3532 32908 3566 32925
rect 3690 33299 3724 33316
rect 3690 33231 3724 33239
rect 3690 33163 3724 33167
rect 3690 33057 3724 33061
rect 3690 32985 3724 32993
rect 3690 32908 3724 32925
rect 3848 33299 3882 33316
rect 3848 33231 3882 33239
rect 3848 33163 3882 33167
rect 3848 33057 3882 33061
rect 3848 32985 3882 32993
rect 3848 32908 3882 32925
rect 4006 33299 4040 33316
rect 4006 33231 4040 33239
rect 4006 33163 4040 33167
rect 4006 33057 4040 33061
rect 4006 32985 4040 32993
rect 4006 32908 4040 32925
rect 4164 33299 4198 33316
rect 4164 33231 4198 33239
rect 4164 33163 4198 33167
rect 4164 33057 4198 33061
rect 4164 32985 4198 32993
rect 4164 32908 4198 32925
rect 4322 33299 4356 33316
rect 4322 33231 4356 33239
rect 4322 33163 4356 33167
rect 4322 33057 4356 33061
rect 4322 32985 4356 32993
rect 4322 32908 4356 32925
rect 4480 33299 4514 33316
rect 4480 33231 4514 33239
rect 4480 33163 4514 33167
rect 4480 33057 4514 33061
rect 4480 32985 4514 32993
rect 4480 32908 4514 32925
rect 2946 32831 2979 32865
rect 3013 32831 3046 32865
rect 3104 32831 3137 32865
rect 3171 32831 3204 32865
rect 3262 32831 3295 32865
rect 3329 32831 3362 32865
rect 3420 32831 3453 32865
rect 3487 32831 3520 32865
rect 3578 32831 3611 32865
rect 3645 32831 3678 32865
rect 3736 32831 3769 32865
rect 3803 32831 3836 32865
rect 3894 32831 3927 32865
rect 3961 32831 3994 32865
rect 4052 32831 4085 32865
rect 4119 32831 4152 32865
rect 4210 32831 4243 32865
rect 4277 32831 4310 32865
rect 4368 32831 4401 32865
rect 4435 32831 4468 32865
rect 2743 32727 4468 32831
rect 2743 32618 2759 32727
rect 2946 32693 2979 32727
rect 3013 32693 3046 32727
rect 3104 32693 3137 32727
rect 3171 32693 3204 32727
rect 3262 32693 3295 32727
rect 3329 32693 3362 32727
rect 3420 32693 3453 32727
rect 3487 32693 3520 32727
rect 3578 32693 3611 32727
rect 3645 32693 3678 32727
rect 3736 32693 3769 32727
rect 3803 32693 3836 32727
rect 3894 32693 3927 32727
rect 3961 32693 3994 32727
rect 4052 32693 4085 32727
rect 4119 32693 4152 32727
rect 4210 32693 4243 32727
rect 4277 32693 4310 32727
rect 4368 32693 4401 32727
rect 4435 32693 4468 32727
rect 2405 32602 2759 32618
rect 2900 32640 2934 32659
rect 2023 32505 2057 32539
rect 2137 32539 2203 32571
rect 2137 32505 2153 32539
rect 2187 32505 2203 32539
rect 2137 32473 2203 32505
rect 2283 32505 2317 32539
rect 2023 32409 2057 32471
rect 2283 32409 2317 32471
rect 2900 32572 2934 32574
rect 2900 32536 2934 32538
rect 2900 32451 2934 32470
rect 3058 32640 3092 32659
rect 3058 32572 3092 32574
rect 3058 32536 3092 32538
rect 3058 32451 3092 32470
rect 3216 32640 3250 32659
rect 3216 32572 3250 32574
rect 3216 32536 3250 32538
rect 3216 32451 3250 32470
rect 3374 32640 3408 32659
rect 3374 32572 3408 32574
rect 3374 32536 3408 32538
rect 3374 32451 3408 32470
rect 3532 32640 3566 32659
rect 3532 32572 3566 32574
rect 3532 32536 3566 32538
rect 3532 32451 3566 32470
rect 3690 32640 3724 32659
rect 3690 32572 3724 32574
rect 3690 32536 3724 32538
rect 3690 32451 3724 32470
rect 3848 32640 3882 32659
rect 3848 32572 3882 32574
rect 3848 32536 3882 32538
rect 3848 32451 3882 32470
rect 4006 32640 4040 32659
rect 4006 32572 4040 32574
rect 4006 32536 4040 32538
rect 4006 32451 4040 32470
rect 4164 32640 4198 32659
rect 4164 32572 4198 32574
rect 4164 32536 4198 32538
rect 4164 32451 4198 32470
rect 4322 32640 4356 32659
rect 4322 32572 4356 32574
rect 4322 32536 4356 32538
rect 4322 32451 4356 32470
rect 4480 32640 4514 32659
rect 4480 32572 4514 32574
rect 4480 32536 4514 32538
rect 4480 32451 4514 32470
rect 2023 32375 2119 32409
rect 2153 32375 2187 32409
rect 2221 32375 2317 32409
rect -50465 32349 -48815 32365
rect -50465 32243 -50449 32349
rect -48831 32243 -48815 32349
rect -50465 32227 -48815 32243
rect 1963 32359 2317 32375
rect 1963 32253 1979 32359
rect 2301 32253 2317 32359
rect 1963 32237 2317 32253
rect 2882 32349 4532 32365
rect 2882 32243 2898 32349
rect 4516 32243 4532 32349
rect 2882 32227 4532 32243
rect -50899 32131 -50803 32165
rect -50769 32131 -50735 32165
rect -50701 32149 -50467 32165
rect -50701 32131 -50589 32149
rect -50899 32069 -50865 32131
rect -50639 32069 -50589 32131
rect -50899 32001 -50865 32035
rect -50801 32035 -50703 32051
rect -50801 32001 -50769 32035
rect -50735 32001 -50703 32035
rect -50801 31985 -50703 32001
rect -50605 32035 -50589 32069
rect -50639 32001 -50589 32035
rect -50899 31905 -50865 31967
rect -50605 31967 -50589 32001
rect -50639 31905 -50589 31967
rect -50899 31871 -50803 31905
rect -50769 31871 -50735 31905
rect -50701 31871 -50589 31905
rect -50605 31827 -50589 31871
rect -50483 31827 -50467 32149
rect -50605 31811 -50467 31827
rect -47362 24973 -47284 24984
rect -47362 24954 -47340 24973
rect -47306 24954 -47284 24973
rect -47362 24712 -47356 24954
rect -47286 24712 -47284 24954
rect -42524 5414 -42490 5441
rect -42524 5342 -42490 5360
rect -42524 5270 -42490 5292
rect -42524 5198 -42490 5224
rect -42524 5126 -42490 5156
rect -42524 5054 -42490 5088
rect -42524 4986 -42490 5020
rect -42524 4918 -42490 4948
rect -42524 4850 -42490 4876
rect -42524 4782 -42490 4804
rect -42524 4714 -42490 4732
rect -42524 4633 -42490 4660
rect -42428 5414 -42394 5441
rect -42428 5342 -42394 5360
rect -42428 5270 -42394 5292
rect -42428 5198 -42394 5224
rect -42428 5126 -42394 5156
rect -42428 5054 -42394 5088
rect -42428 4986 -42394 5020
rect -42428 4918 -42394 4948
rect -42428 4850 -42394 4876
rect -42428 4782 -42394 4804
rect -42428 4714 -42394 4732
rect -42428 4633 -42394 4660
rect -42332 5414 -42298 5441
rect -42332 5342 -42298 5360
rect -42332 5270 -42298 5292
rect -42332 5198 -42298 5224
rect -42332 5126 -42298 5156
rect -42332 5054 -42298 5088
rect -42332 4986 -42298 5020
rect -42332 4918 -42298 4948
rect -42332 4850 -42298 4876
rect -42332 4782 -42298 4804
rect -42332 4714 -42298 4732
rect -42332 4633 -42298 4660
rect -42236 5414 -42202 5441
rect -42236 5342 -42202 5360
rect -42236 5270 -42202 5292
rect -42236 5198 -42202 5224
rect -42236 5126 -42202 5156
rect -42236 5054 -42202 5088
rect -42236 4986 -42202 5020
rect -42236 4918 -42202 4948
rect -42236 4850 -42202 4876
rect -42236 4782 -42202 4804
rect -42236 4714 -42202 4732
rect -42236 4633 -42202 4660
rect -42140 5414 -42106 5441
rect -42140 5342 -42106 5360
rect -42140 5270 -42106 5292
rect -42140 5198 -42106 5224
rect -42140 5126 -42106 5156
rect -42140 5054 -42106 5088
rect -42140 4986 -42106 5020
rect -42140 4918 -42106 4948
rect -42140 4850 -42106 4876
rect -42140 4782 -42106 4804
rect -42140 4714 -42106 4732
rect -42140 4633 -42106 4660
rect -42044 5414 -42010 5441
rect -42044 5342 -42010 5360
rect -42044 5270 -42010 5292
rect -42044 5198 -42010 5224
rect -42044 5126 -42010 5156
rect -42044 5054 -42010 5088
rect -42044 4986 -42010 5020
rect -42044 4918 -42010 4948
rect -42044 4850 -42010 4876
rect -42044 4782 -42010 4804
rect -42044 4714 -42010 4732
rect -42044 4633 -42010 4660
rect -41948 5414 -41914 5441
rect -41948 5342 -41914 5360
rect -41948 5270 -41914 5292
rect -41948 5198 -41914 5224
rect -41948 5126 -41914 5156
rect -41948 5054 -41914 5088
rect -41948 4986 -41914 5020
rect -41948 4918 -41914 4948
rect -41948 4850 -41914 4876
rect -41948 4782 -41914 4804
rect -41948 4714 -41914 4732
rect -41948 4633 -41914 4660
rect -41852 5414 -41818 5441
rect -41852 5342 -41818 5360
rect -41852 5270 -41818 5292
rect -41852 5198 -41818 5224
rect -41852 5126 -41818 5156
rect -41852 5054 -41818 5088
rect -41852 4986 -41818 5020
rect -41852 4918 -41818 4948
rect -41852 4850 -41818 4876
rect -41852 4782 -41818 4804
rect -41852 4714 -41818 4732
rect -41852 4633 -41818 4660
rect -41756 5414 -41722 5441
rect -41756 5342 -41722 5360
rect -41756 5270 -41722 5292
rect -41756 5198 -41722 5224
rect -41756 5126 -41722 5156
rect -41756 5054 -41722 5088
rect -41756 4986 -41722 5020
rect -41756 4918 -41722 4948
rect -41756 4850 -41722 4876
rect -41756 4782 -41722 4804
rect -41756 4714 -41722 4732
rect -41756 4633 -41722 4660
rect -41660 5414 -41626 5441
rect -41660 5342 -41626 5360
rect -41660 5270 -41626 5292
rect -41660 5198 -41626 5224
rect -41660 5126 -41626 5156
rect -41660 5054 -41626 5088
rect -41660 4986 -41626 5020
rect -41660 4918 -41626 4948
rect -41660 4850 -41626 4876
rect -41660 4782 -41626 4804
rect -41660 4714 -41626 4732
rect -41660 4633 -41626 4660
rect -41564 5414 -41530 5441
rect -41564 5342 -41530 5360
rect -41564 5270 -41530 5292
rect -41564 5198 -41530 5224
rect -41564 5126 -41530 5156
rect -41564 5054 -41530 5088
rect -41564 4986 -41530 5020
rect -41564 4918 -41530 4948
rect -41564 4850 -41530 4876
rect -41564 4782 -41530 4804
rect -41564 4714 -41530 4732
rect -41564 4633 -41530 4660
rect -41468 5414 -41434 5441
rect -41468 5342 -41434 5360
rect -41468 5270 -41434 5292
rect -41468 5198 -41434 5224
rect -41468 5126 -41434 5156
rect -41468 5054 -41434 5088
rect -41468 4986 -41434 5020
rect -41468 4918 -41434 4948
rect -41468 4850 -41434 4876
rect -41468 4782 -41434 4804
rect -41468 4714 -41434 4732
rect -41468 4633 -41434 4660
rect -41372 5414 -41338 5441
rect -41372 5342 -41338 5360
rect -41372 5270 -41338 5292
rect -41372 5198 -41338 5224
rect -41372 5126 -41338 5156
rect -41372 5054 -41338 5088
rect -41372 4986 -41338 5020
rect -41372 4918 -41338 4948
rect -41372 4850 -41338 4876
rect -41372 4782 -41338 4804
rect -41372 4714 -41338 4732
rect -41372 4633 -41338 4660
rect -41276 5414 -41242 5441
rect -41276 5342 -41242 5360
rect -41276 5270 -41242 5292
rect -41276 5198 -41242 5224
rect -41276 5126 -41242 5156
rect -41276 5054 -41242 5088
rect -41276 4986 -41242 5020
rect -41276 4918 -41242 4948
rect -41276 4850 -41242 4876
rect -41276 4782 -41242 4804
rect -41276 4714 -41242 4732
rect -41276 4633 -41242 4660
rect -41180 5414 -41146 5441
rect -41180 5342 -41146 5360
rect -41180 5270 -41146 5292
rect -41180 5198 -41146 5224
rect -41180 5126 -41146 5156
rect -41180 5054 -41146 5088
rect -41180 4986 -41146 5020
rect -41180 4918 -41146 4948
rect -41180 4850 -41146 4876
rect -41180 4782 -41146 4804
rect -41180 4714 -41146 4732
rect -41180 4633 -41146 4660
rect -41084 5414 -41050 5441
rect -41084 5342 -41050 5360
rect -41084 5270 -41050 5292
rect -41084 5198 -41050 5224
rect -41084 5126 -41050 5156
rect -41084 5054 -41050 5088
rect -41084 4986 -41050 5020
rect -41084 4918 -41050 4948
rect -41084 4850 -41050 4876
rect -41084 4782 -41050 4804
rect -41084 4714 -41050 4732
rect -41084 4633 -41050 4660
rect -40988 5414 -40954 5441
rect -40988 5342 -40954 5360
rect -40988 5270 -40954 5292
rect -40988 5198 -40954 5224
rect -40988 5126 -40954 5156
rect -40988 5054 -40954 5088
rect -40988 4986 -40954 5020
rect -40988 4918 -40954 4948
rect -40988 4850 -40954 4876
rect -40988 4782 -40954 4804
rect -40988 4714 -40954 4732
rect -40988 4633 -40954 4660
rect -40892 5414 -40858 5441
rect -40892 5342 -40858 5360
rect -40892 5270 -40858 5292
rect -40892 5198 -40858 5224
rect -40892 5126 -40858 5156
rect -40892 5054 -40858 5088
rect -40892 4986 -40858 5020
rect -40892 4918 -40858 4948
rect -40892 4850 -40858 4876
rect -40892 4782 -40858 4804
rect -40892 4714 -40858 4732
rect -40892 4633 -40858 4660
rect -40796 5414 -40762 5441
rect -40796 5342 -40762 5360
rect -40796 5270 -40762 5292
rect -40796 5198 -40762 5224
rect -40796 5126 -40762 5156
rect -40796 5054 -40762 5088
rect -40796 4986 -40762 5020
rect -40796 4918 -40762 4948
rect -40796 4850 -40762 4876
rect -40796 4782 -40762 4804
rect -40796 4714 -40762 4732
rect -40796 4633 -40762 4660
rect -40700 5414 -40666 5441
rect -40700 5342 -40666 5360
rect -40700 5270 -40666 5292
rect -40700 5198 -40666 5224
rect -40700 5126 -40666 5156
rect -40700 5054 -40666 5088
rect -40700 4986 -40666 5020
rect -40700 4918 -40666 4948
rect -40700 4850 -40666 4876
rect -40700 4782 -40666 4804
rect -40700 4714 -40666 4732
rect -40700 4633 -40666 4660
rect 104 5402 138 5429
rect 104 5330 138 5348
rect 104 5258 138 5280
rect 104 5186 138 5212
rect 104 5114 138 5144
rect 104 5042 138 5076
rect 104 4974 138 5008
rect 104 4906 138 4936
rect 104 4838 138 4864
rect 104 4770 138 4792
rect 104 4702 138 4720
rect 104 4621 138 4648
rect 200 5402 234 5429
rect 200 5330 234 5348
rect 200 5258 234 5280
rect 200 5186 234 5212
rect 200 5114 234 5144
rect 200 5042 234 5076
rect 200 4974 234 5008
rect 200 4906 234 4936
rect 200 4838 234 4864
rect 200 4770 234 4792
rect 200 4702 234 4720
rect 200 4621 234 4648
rect 296 5402 330 5429
rect 296 5330 330 5348
rect 296 5258 330 5280
rect 296 5186 330 5212
rect 296 5114 330 5144
rect 296 5042 330 5076
rect 296 4974 330 5008
rect 296 4906 330 4936
rect 296 4838 330 4864
rect 296 4770 330 4792
rect 296 4702 330 4720
rect 296 4621 330 4648
rect 392 5402 426 5429
rect 392 5330 426 5348
rect 392 5258 426 5280
rect 392 5186 426 5212
rect 392 5114 426 5144
rect 392 5042 426 5076
rect 392 4974 426 5008
rect 392 4906 426 4936
rect 392 4838 426 4864
rect 392 4770 426 4792
rect 392 4702 426 4720
rect 392 4621 426 4648
rect 488 5402 522 5429
rect 488 5330 522 5348
rect 488 5258 522 5280
rect 488 5186 522 5212
rect 488 5114 522 5144
rect 488 5042 522 5076
rect 488 4974 522 5008
rect 488 4906 522 4936
rect 488 4838 522 4864
rect 488 4770 522 4792
rect 488 4702 522 4720
rect 488 4621 522 4648
rect 584 5402 618 5429
rect 584 5330 618 5348
rect 584 5258 618 5280
rect 584 5186 618 5212
rect 584 5114 618 5144
rect 584 5042 618 5076
rect 584 4974 618 5008
rect 584 4906 618 4936
rect 584 4838 618 4864
rect 584 4770 618 4792
rect 584 4702 618 4720
rect 584 4621 618 4648
rect 680 5402 714 5429
rect 680 5330 714 5348
rect 680 5258 714 5280
rect 680 5186 714 5212
rect 680 5114 714 5144
rect 680 5042 714 5076
rect 680 4974 714 5008
rect 680 4906 714 4936
rect 680 4838 714 4864
rect 680 4770 714 4792
rect 680 4702 714 4720
rect 680 4621 714 4648
rect 776 5402 810 5429
rect 776 5330 810 5348
rect 776 5258 810 5280
rect 776 5186 810 5212
rect 776 5114 810 5144
rect 776 5042 810 5076
rect 776 4974 810 5008
rect 776 4906 810 4936
rect 776 4838 810 4864
rect 776 4770 810 4792
rect 776 4702 810 4720
rect 776 4621 810 4648
rect 872 5402 906 5429
rect 872 5330 906 5348
rect 872 5258 906 5280
rect 872 5186 906 5212
rect 872 5114 906 5144
rect 872 5042 906 5076
rect 872 4974 906 5008
rect 872 4906 906 4936
rect 872 4838 906 4864
rect 872 4770 906 4792
rect 872 4702 906 4720
rect 872 4621 906 4648
rect 968 5402 1002 5429
rect 968 5330 1002 5348
rect 968 5258 1002 5280
rect 968 5186 1002 5212
rect 968 5114 1002 5144
rect 968 5042 1002 5076
rect 968 4974 1002 5008
rect 968 4906 1002 4936
rect 968 4838 1002 4864
rect 968 4770 1002 4792
rect 968 4702 1002 4720
rect 968 4621 1002 4648
rect 1064 5402 1098 5429
rect 1064 5330 1098 5348
rect 1064 5258 1098 5280
rect 1064 5186 1098 5212
rect 1064 5114 1098 5144
rect 1064 5042 1098 5076
rect 1064 4974 1098 5008
rect 1064 4906 1098 4936
rect 1064 4838 1098 4864
rect 1064 4770 1098 4792
rect 1064 4702 1098 4720
rect 1064 4621 1098 4648
rect 1160 5402 1194 5429
rect 1160 5330 1194 5348
rect 1160 5258 1194 5280
rect 1160 5186 1194 5212
rect 1160 5114 1194 5144
rect 1160 5042 1194 5076
rect 1160 4974 1194 5008
rect 1160 4906 1194 4936
rect 1160 4838 1194 4864
rect 1160 4770 1194 4792
rect 1160 4702 1194 4720
rect 1160 4621 1194 4648
rect 1256 5402 1290 5429
rect 1256 5330 1290 5348
rect 1256 5258 1290 5280
rect 1256 5186 1290 5212
rect 1256 5114 1290 5144
rect 1256 5042 1290 5076
rect 1256 4974 1290 5008
rect 1256 4906 1290 4936
rect 1256 4838 1290 4864
rect 1256 4770 1290 4792
rect 1256 4702 1290 4720
rect 1256 4621 1290 4648
rect 1352 5402 1386 5429
rect 1352 5330 1386 5348
rect 1352 5258 1386 5280
rect 1352 5186 1386 5212
rect 1352 5114 1386 5144
rect 1352 5042 1386 5076
rect 1352 4974 1386 5008
rect 1352 4906 1386 4936
rect 1352 4838 1386 4864
rect 1352 4770 1386 4792
rect 1352 4702 1386 4720
rect 1352 4621 1386 4648
rect 1448 5402 1482 5429
rect 1448 5330 1482 5348
rect 1448 5258 1482 5280
rect 1448 5186 1482 5212
rect 1448 5114 1482 5144
rect 1448 5042 1482 5076
rect 1448 4974 1482 5008
rect 1448 4906 1482 4936
rect 1448 4838 1482 4864
rect 1448 4770 1482 4792
rect 1448 4702 1482 4720
rect 1448 4621 1482 4648
rect 1544 5402 1578 5429
rect 1544 5330 1578 5348
rect 1544 5258 1578 5280
rect 1544 5186 1578 5212
rect 1544 5114 1578 5144
rect 1544 5042 1578 5076
rect 1544 4974 1578 5008
rect 1544 4906 1578 4936
rect 1544 4838 1578 4864
rect 1544 4770 1578 4792
rect 1544 4702 1578 4720
rect 1544 4621 1578 4648
rect 1640 5402 1674 5429
rect 1640 5330 1674 5348
rect 1640 5258 1674 5280
rect 1640 5186 1674 5212
rect 1640 5114 1674 5144
rect 1640 5042 1674 5076
rect 1640 4974 1674 5008
rect 1640 4906 1674 4936
rect 1640 4838 1674 4864
rect 1640 4770 1674 4792
rect 1640 4702 1674 4720
rect 1640 4621 1674 4648
rect 1736 5402 1770 5429
rect 1736 5330 1770 5348
rect 1736 5258 1770 5280
rect 1736 5186 1770 5212
rect 1736 5114 1770 5144
rect 1736 5042 1770 5076
rect 1736 4974 1770 5008
rect 1736 4906 1770 4936
rect 1736 4838 1770 4864
rect 1736 4770 1770 4792
rect 1736 4702 1770 4720
rect 1736 4621 1770 4648
rect 1832 5402 1866 5429
rect 1832 5330 1866 5348
rect 1832 5258 1866 5280
rect 1832 5186 1866 5212
rect 1832 5114 1866 5144
rect 1832 5042 1866 5076
rect 1832 4974 1866 5008
rect 1832 4906 1866 4936
rect 1832 4838 1866 4864
rect 1832 4770 1866 4792
rect 1832 4702 1866 4720
rect 1832 4621 1866 4648
rect 1928 5402 1962 5429
rect 1928 5330 1962 5348
rect 1928 5258 1962 5280
rect 1928 5186 1962 5212
rect 1928 5114 1962 5144
rect 1928 5042 1962 5076
rect 1928 4974 1962 5008
rect 1928 4906 1962 4936
rect 1928 4838 1962 4864
rect 1928 4770 1962 4792
rect 1928 4702 1962 4720
rect 1928 4621 1962 4648
rect -42834 4567 -40734 4583
rect -42834 4533 -42440 4567
rect -42406 4533 -42368 4567
rect -42334 4533 -42296 4567
rect -42262 4533 -42224 4567
rect -42190 4533 -42152 4567
rect -42118 4533 -42080 4567
rect -42046 4533 -42008 4567
rect -41974 4533 -41936 4567
rect -41902 4533 -41864 4567
rect -41830 4533 -41792 4567
rect -41758 4533 -41720 4567
rect -41686 4533 -41648 4567
rect -41614 4533 -41576 4567
rect -41542 4533 -41504 4567
rect -41470 4533 -41432 4567
rect -41398 4533 -41360 4567
rect -41326 4533 -41288 4567
rect -41254 4533 -41216 4567
rect -41182 4533 -41144 4567
rect -41110 4533 -41072 4567
rect -41038 4533 -41000 4567
rect -40966 4533 -40928 4567
rect -40894 4533 -40856 4567
rect -40822 4533 -40784 4567
rect -40750 4533 -40734 4567
rect -42834 4495 -40734 4533
rect -42834 4461 -42440 4495
rect -42406 4461 -42368 4495
rect -42334 4461 -42296 4495
rect -42262 4461 -42224 4495
rect -42190 4461 -42152 4495
rect -42118 4461 -42080 4495
rect -42046 4461 -42008 4495
rect -41974 4461 -41936 4495
rect -41902 4461 -41864 4495
rect -41830 4461 -41792 4495
rect -41758 4461 -41720 4495
rect -41686 4461 -41648 4495
rect -41614 4461 -41576 4495
rect -41542 4461 -41504 4495
rect -41470 4461 -41432 4495
rect -41398 4461 -41360 4495
rect -41326 4461 -41288 4495
rect -41254 4461 -41216 4495
rect -41182 4461 -41144 4495
rect -41110 4461 -41072 4495
rect -41038 4461 -41000 4495
rect -40966 4461 -40928 4495
rect -40894 4461 -40856 4495
rect -40822 4461 -40784 4495
rect -40750 4461 -40734 4495
rect -42834 4445 -40734 4461
rect 172 4560 2404 4576
rect 172 4526 188 4560
rect 222 4526 260 4560
rect 294 4526 332 4560
rect 366 4526 404 4560
rect 438 4526 476 4560
rect 510 4526 548 4560
rect 582 4526 620 4560
rect 654 4526 692 4560
rect 726 4526 764 4560
rect 798 4526 836 4560
rect 870 4526 908 4560
rect 942 4526 980 4560
rect 1014 4526 1052 4560
rect 1086 4526 1124 4560
rect 1158 4526 1196 4560
rect 1230 4526 1268 4560
rect 1302 4526 1340 4560
rect 1374 4526 1412 4560
rect 1446 4526 1484 4560
rect 1518 4526 1556 4560
rect 1590 4526 1628 4560
rect 1662 4526 1700 4560
rect 1734 4526 1772 4560
rect 1806 4526 1844 4560
rect 1878 4526 2404 4560
rect 172 4488 2404 4526
rect 172 4454 188 4488
rect 222 4454 260 4488
rect 294 4454 332 4488
rect 366 4454 404 4488
rect 438 4454 476 4488
rect 510 4454 548 4488
rect 582 4454 620 4488
rect 654 4454 692 4488
rect 726 4454 764 4488
rect 798 4454 836 4488
rect 870 4454 908 4488
rect 942 4454 980 4488
rect 1014 4454 1052 4488
rect 1086 4454 1124 4488
rect 1158 4454 1196 4488
rect 1230 4454 1268 4488
rect 1302 4454 1340 4488
rect 1374 4454 1412 4488
rect 1446 4454 1484 4488
rect 1518 4454 1556 4488
rect 1590 4454 1628 4488
rect 1662 4454 1700 4488
rect 1734 4454 1772 4488
rect 1806 4454 1844 4488
rect 1878 4454 2404 4488
rect 172 4438 2404 4454
rect -42525 -4760 -42491 -4733
rect -42525 -4832 -42491 -4814
rect -42525 -4904 -42491 -4882
rect -42525 -4976 -42491 -4950
rect -42525 -5048 -42491 -5018
rect -42525 -5120 -42491 -5086
rect -42525 -5188 -42491 -5154
rect -42525 -5256 -42491 -5226
rect -42525 -5324 -42491 -5298
rect -42525 -5392 -42491 -5370
rect -42525 -5460 -42491 -5442
rect -42525 -5541 -42491 -5514
rect -42429 -4760 -42395 -4733
rect -42429 -4832 -42395 -4814
rect -42429 -4904 -42395 -4882
rect -42429 -4976 -42395 -4950
rect -42429 -5048 -42395 -5018
rect -42429 -5120 -42395 -5086
rect -42429 -5188 -42395 -5154
rect -42429 -5256 -42395 -5226
rect -42429 -5324 -42395 -5298
rect -42429 -5392 -42395 -5370
rect -42429 -5460 -42395 -5442
rect -42429 -5541 -42395 -5514
rect -42333 -4760 -42299 -4733
rect -42333 -4832 -42299 -4814
rect -42333 -4904 -42299 -4882
rect -42333 -4976 -42299 -4950
rect -42333 -5048 -42299 -5018
rect -42333 -5120 -42299 -5086
rect -42333 -5188 -42299 -5154
rect -42333 -5256 -42299 -5226
rect -42333 -5324 -42299 -5298
rect -42333 -5392 -42299 -5370
rect -42333 -5460 -42299 -5442
rect -42333 -5541 -42299 -5514
rect -42237 -4760 -42203 -4733
rect -42237 -4832 -42203 -4814
rect -42237 -4904 -42203 -4882
rect -42237 -4976 -42203 -4950
rect -42237 -5048 -42203 -5018
rect -42237 -5120 -42203 -5086
rect -42237 -5188 -42203 -5154
rect -42237 -5256 -42203 -5226
rect -42237 -5324 -42203 -5298
rect -42237 -5392 -42203 -5370
rect -42237 -5460 -42203 -5442
rect -42237 -5541 -42203 -5514
rect -42141 -4760 -42107 -4733
rect -42141 -4832 -42107 -4814
rect -42141 -4904 -42107 -4882
rect -42141 -4976 -42107 -4950
rect -42141 -5048 -42107 -5018
rect -42141 -5120 -42107 -5086
rect -42141 -5188 -42107 -5154
rect -42141 -5256 -42107 -5226
rect -42141 -5324 -42107 -5298
rect -42141 -5392 -42107 -5370
rect -42141 -5460 -42107 -5442
rect -42141 -5541 -42107 -5514
rect -42045 -4760 -42011 -4733
rect -42045 -4832 -42011 -4814
rect -42045 -4904 -42011 -4882
rect -42045 -4976 -42011 -4950
rect -42045 -5048 -42011 -5018
rect -42045 -5120 -42011 -5086
rect -42045 -5188 -42011 -5154
rect -42045 -5256 -42011 -5226
rect -42045 -5324 -42011 -5298
rect -42045 -5392 -42011 -5370
rect -42045 -5460 -42011 -5442
rect -42045 -5541 -42011 -5514
rect -41949 -4760 -41915 -4733
rect -41949 -4832 -41915 -4814
rect -41949 -4904 -41915 -4882
rect -41949 -4976 -41915 -4950
rect -41949 -5048 -41915 -5018
rect -41949 -5120 -41915 -5086
rect -41949 -5188 -41915 -5154
rect -41949 -5256 -41915 -5226
rect -41949 -5324 -41915 -5298
rect -41949 -5392 -41915 -5370
rect -41949 -5460 -41915 -5442
rect -41949 -5541 -41915 -5514
rect -41853 -4760 -41819 -4733
rect -41853 -4832 -41819 -4814
rect -41853 -4904 -41819 -4882
rect -41853 -4976 -41819 -4950
rect -41853 -5048 -41819 -5018
rect -41853 -5120 -41819 -5086
rect -41853 -5188 -41819 -5154
rect -41853 -5256 -41819 -5226
rect -41853 -5324 -41819 -5298
rect -41853 -5392 -41819 -5370
rect -41853 -5460 -41819 -5442
rect -41853 -5541 -41819 -5514
rect -41757 -4760 -41723 -4733
rect -41757 -4832 -41723 -4814
rect -41757 -4904 -41723 -4882
rect -41757 -4976 -41723 -4950
rect -41757 -5048 -41723 -5018
rect -41757 -5120 -41723 -5086
rect -41757 -5188 -41723 -5154
rect -41757 -5256 -41723 -5226
rect -41757 -5324 -41723 -5298
rect -41757 -5392 -41723 -5370
rect -41757 -5460 -41723 -5442
rect -41757 -5541 -41723 -5514
rect -41661 -4760 -41627 -4733
rect -41661 -4832 -41627 -4814
rect -41661 -4904 -41627 -4882
rect -41661 -4976 -41627 -4950
rect -41661 -5048 -41627 -5018
rect -41661 -5120 -41627 -5086
rect -41661 -5188 -41627 -5154
rect -41661 -5256 -41627 -5226
rect -41661 -5324 -41627 -5298
rect -41661 -5392 -41627 -5370
rect -41661 -5460 -41627 -5442
rect -41661 -5541 -41627 -5514
rect -41565 -4760 -41531 -4733
rect -41565 -4832 -41531 -4814
rect -41565 -4904 -41531 -4882
rect -41565 -4976 -41531 -4950
rect -41565 -5048 -41531 -5018
rect -41565 -5120 -41531 -5086
rect -41565 -5188 -41531 -5154
rect -41565 -5256 -41531 -5226
rect -41565 -5324 -41531 -5298
rect -41565 -5392 -41531 -5370
rect -41565 -5460 -41531 -5442
rect -41565 -5541 -41531 -5514
rect -41469 -4760 -41435 -4733
rect -41469 -4832 -41435 -4814
rect -41469 -4904 -41435 -4882
rect -41469 -4976 -41435 -4950
rect -41469 -5048 -41435 -5018
rect -41469 -5120 -41435 -5086
rect -41469 -5188 -41435 -5154
rect -41469 -5256 -41435 -5226
rect -41469 -5324 -41435 -5298
rect -41469 -5392 -41435 -5370
rect -41469 -5460 -41435 -5442
rect -41469 -5541 -41435 -5514
rect -41373 -4760 -41339 -4733
rect -41373 -4832 -41339 -4814
rect -41373 -4904 -41339 -4882
rect -41373 -4976 -41339 -4950
rect -41373 -5048 -41339 -5018
rect -41373 -5120 -41339 -5086
rect -41373 -5188 -41339 -5154
rect -41373 -5256 -41339 -5226
rect -41373 -5324 -41339 -5298
rect -41373 -5392 -41339 -5370
rect -41373 -5460 -41339 -5442
rect -41373 -5541 -41339 -5514
rect -41277 -4760 -41243 -4733
rect -41277 -4832 -41243 -4814
rect -41277 -4904 -41243 -4882
rect -41277 -4976 -41243 -4950
rect -41277 -5048 -41243 -5018
rect -41277 -5120 -41243 -5086
rect -41277 -5188 -41243 -5154
rect -41277 -5256 -41243 -5226
rect -41277 -5324 -41243 -5298
rect -41277 -5392 -41243 -5370
rect -41277 -5460 -41243 -5442
rect -41277 -5541 -41243 -5514
rect -41181 -4760 -41147 -4733
rect -41181 -4832 -41147 -4814
rect -41181 -4904 -41147 -4882
rect -41181 -4976 -41147 -4950
rect -41181 -5048 -41147 -5018
rect -41181 -5120 -41147 -5086
rect -41181 -5188 -41147 -5154
rect -41181 -5256 -41147 -5226
rect -41181 -5324 -41147 -5298
rect -41181 -5392 -41147 -5370
rect -41181 -5460 -41147 -5442
rect -41181 -5541 -41147 -5514
rect -41085 -4760 -41051 -4733
rect -41085 -4832 -41051 -4814
rect -41085 -4904 -41051 -4882
rect -41085 -4976 -41051 -4950
rect -41085 -5048 -41051 -5018
rect -41085 -5120 -41051 -5086
rect -41085 -5188 -41051 -5154
rect -41085 -5256 -41051 -5226
rect -41085 -5324 -41051 -5298
rect -41085 -5392 -41051 -5370
rect -41085 -5460 -41051 -5442
rect -41085 -5541 -41051 -5514
rect -40989 -4760 -40955 -4733
rect -40989 -4832 -40955 -4814
rect -40989 -4904 -40955 -4882
rect -40989 -4976 -40955 -4950
rect -40989 -5048 -40955 -5018
rect -40989 -5120 -40955 -5086
rect -40989 -5188 -40955 -5154
rect -40989 -5256 -40955 -5226
rect -40989 -5324 -40955 -5298
rect -40989 -5392 -40955 -5370
rect -40989 -5460 -40955 -5442
rect -40989 -5541 -40955 -5514
rect -40893 -4760 -40859 -4733
rect -40893 -4832 -40859 -4814
rect -40893 -4904 -40859 -4882
rect -40893 -4976 -40859 -4950
rect -40893 -5048 -40859 -5018
rect -40893 -5120 -40859 -5086
rect -40893 -5188 -40859 -5154
rect -40893 -5256 -40859 -5226
rect -40893 -5324 -40859 -5298
rect -40893 -5392 -40859 -5370
rect -40893 -5460 -40859 -5442
rect -40893 -5541 -40859 -5514
rect -40797 -4760 -40763 -4733
rect -40797 -4832 -40763 -4814
rect -40797 -4904 -40763 -4882
rect -40797 -4976 -40763 -4950
rect -40797 -5048 -40763 -5018
rect -40797 -5120 -40763 -5086
rect -40797 -5188 -40763 -5154
rect -40797 -5256 -40763 -5226
rect -40797 -5324 -40763 -5298
rect -40797 -5392 -40763 -5370
rect -40797 -5460 -40763 -5442
rect -40797 -5541 -40763 -5514
rect -40701 -4760 -40667 -4733
rect -40701 -4832 -40667 -4814
rect -40701 -4904 -40667 -4882
rect -40701 -4976 -40667 -4950
rect -40701 -5048 -40667 -5018
rect -40701 -5120 -40667 -5086
rect -40701 -5188 -40667 -5154
rect -40701 -5256 -40667 -5226
rect -40701 -5324 -40667 -5298
rect -40701 -5392 -40667 -5370
rect -40701 -5460 -40667 -5442
rect -40701 -5541 -40667 -5514
rect 116 -4786 150 -4759
rect 116 -4858 150 -4840
rect 116 -4930 150 -4908
rect 116 -5002 150 -4976
rect 116 -5074 150 -5044
rect 116 -5146 150 -5112
rect 116 -5214 150 -5180
rect 116 -5282 150 -5252
rect 116 -5350 150 -5324
rect 116 -5418 150 -5396
rect 116 -5486 150 -5468
rect 116 -5567 150 -5540
rect 212 -4786 246 -4759
rect 212 -4858 246 -4840
rect 212 -4930 246 -4908
rect 212 -5002 246 -4976
rect 212 -5074 246 -5044
rect 212 -5146 246 -5112
rect 212 -5214 246 -5180
rect 212 -5282 246 -5252
rect 212 -5350 246 -5324
rect 212 -5418 246 -5396
rect 212 -5486 246 -5468
rect 212 -5567 246 -5540
rect 308 -4786 342 -4759
rect 308 -4858 342 -4840
rect 308 -4930 342 -4908
rect 308 -5002 342 -4976
rect 308 -5074 342 -5044
rect 308 -5146 342 -5112
rect 308 -5214 342 -5180
rect 308 -5282 342 -5252
rect 308 -5350 342 -5324
rect 308 -5418 342 -5396
rect 308 -5486 342 -5468
rect 308 -5567 342 -5540
rect 404 -4786 438 -4759
rect 404 -4858 438 -4840
rect 404 -4930 438 -4908
rect 404 -5002 438 -4976
rect 404 -5074 438 -5044
rect 404 -5146 438 -5112
rect 404 -5214 438 -5180
rect 404 -5282 438 -5252
rect 404 -5350 438 -5324
rect 404 -5418 438 -5396
rect 404 -5486 438 -5468
rect 404 -5567 438 -5540
rect 500 -4786 534 -4759
rect 500 -4858 534 -4840
rect 500 -4930 534 -4908
rect 500 -5002 534 -4976
rect 500 -5074 534 -5044
rect 500 -5146 534 -5112
rect 500 -5214 534 -5180
rect 500 -5282 534 -5252
rect 500 -5350 534 -5324
rect 500 -5418 534 -5396
rect 500 -5486 534 -5468
rect 500 -5567 534 -5540
rect 596 -4786 630 -4759
rect 596 -4858 630 -4840
rect 596 -4930 630 -4908
rect 596 -5002 630 -4976
rect 596 -5074 630 -5044
rect 596 -5146 630 -5112
rect 596 -5214 630 -5180
rect 596 -5282 630 -5252
rect 596 -5350 630 -5324
rect 596 -5418 630 -5396
rect 596 -5486 630 -5468
rect 596 -5567 630 -5540
rect 692 -4786 726 -4759
rect 692 -4858 726 -4840
rect 692 -4930 726 -4908
rect 692 -5002 726 -4976
rect 692 -5074 726 -5044
rect 692 -5146 726 -5112
rect 692 -5214 726 -5180
rect 692 -5282 726 -5252
rect 692 -5350 726 -5324
rect 692 -5418 726 -5396
rect 692 -5486 726 -5468
rect 692 -5567 726 -5540
rect 788 -4786 822 -4759
rect 788 -4858 822 -4840
rect 788 -4930 822 -4908
rect 788 -5002 822 -4976
rect 788 -5074 822 -5044
rect 788 -5146 822 -5112
rect 788 -5214 822 -5180
rect 788 -5282 822 -5252
rect 788 -5350 822 -5324
rect 788 -5418 822 -5396
rect 788 -5486 822 -5468
rect 788 -5567 822 -5540
rect 884 -4786 918 -4759
rect 884 -4858 918 -4840
rect 884 -4930 918 -4908
rect 884 -5002 918 -4976
rect 884 -5074 918 -5044
rect 884 -5146 918 -5112
rect 884 -5214 918 -5180
rect 884 -5282 918 -5252
rect 884 -5350 918 -5324
rect 884 -5418 918 -5396
rect 884 -5486 918 -5468
rect 884 -5567 918 -5540
rect 980 -4786 1014 -4759
rect 980 -4858 1014 -4840
rect 980 -4930 1014 -4908
rect 980 -5002 1014 -4976
rect 980 -5074 1014 -5044
rect 980 -5146 1014 -5112
rect 980 -5214 1014 -5180
rect 980 -5282 1014 -5252
rect 980 -5350 1014 -5324
rect 980 -5418 1014 -5396
rect 980 -5486 1014 -5468
rect 980 -5567 1014 -5540
rect 1076 -4786 1110 -4759
rect 1076 -4858 1110 -4840
rect 1076 -4930 1110 -4908
rect 1076 -5002 1110 -4976
rect 1076 -5074 1110 -5044
rect 1076 -5146 1110 -5112
rect 1076 -5214 1110 -5180
rect 1076 -5282 1110 -5252
rect 1076 -5350 1110 -5324
rect 1076 -5418 1110 -5396
rect 1076 -5486 1110 -5468
rect 1076 -5567 1110 -5540
rect 1172 -4786 1206 -4759
rect 1172 -4858 1206 -4840
rect 1172 -4930 1206 -4908
rect 1172 -5002 1206 -4976
rect 1172 -5074 1206 -5044
rect 1172 -5146 1206 -5112
rect 1172 -5214 1206 -5180
rect 1172 -5282 1206 -5252
rect 1172 -5350 1206 -5324
rect 1172 -5418 1206 -5396
rect 1172 -5486 1206 -5468
rect 1172 -5567 1206 -5540
rect 1268 -4786 1302 -4759
rect 1268 -4858 1302 -4840
rect 1268 -4930 1302 -4908
rect 1268 -5002 1302 -4976
rect 1268 -5074 1302 -5044
rect 1268 -5146 1302 -5112
rect 1268 -5214 1302 -5180
rect 1268 -5282 1302 -5252
rect 1268 -5350 1302 -5324
rect 1268 -5418 1302 -5396
rect 1268 -5486 1302 -5468
rect 1268 -5567 1302 -5540
rect 1364 -4786 1398 -4759
rect 1364 -4858 1398 -4840
rect 1364 -4930 1398 -4908
rect 1364 -5002 1398 -4976
rect 1364 -5074 1398 -5044
rect 1364 -5146 1398 -5112
rect 1364 -5214 1398 -5180
rect 1364 -5282 1398 -5252
rect 1364 -5350 1398 -5324
rect 1364 -5418 1398 -5396
rect 1364 -5486 1398 -5468
rect 1364 -5567 1398 -5540
rect 1460 -4786 1494 -4759
rect 1460 -4858 1494 -4840
rect 1460 -4930 1494 -4908
rect 1460 -5002 1494 -4976
rect 1460 -5074 1494 -5044
rect 1460 -5146 1494 -5112
rect 1460 -5214 1494 -5180
rect 1460 -5282 1494 -5252
rect 1460 -5350 1494 -5324
rect 1460 -5418 1494 -5396
rect 1460 -5486 1494 -5468
rect 1460 -5567 1494 -5540
rect 1556 -4786 1590 -4759
rect 1556 -4858 1590 -4840
rect 1556 -4930 1590 -4908
rect 1556 -5002 1590 -4976
rect 1556 -5074 1590 -5044
rect 1556 -5146 1590 -5112
rect 1556 -5214 1590 -5180
rect 1556 -5282 1590 -5252
rect 1556 -5350 1590 -5324
rect 1556 -5418 1590 -5396
rect 1556 -5486 1590 -5468
rect 1556 -5567 1590 -5540
rect 1652 -4786 1686 -4759
rect 1652 -4858 1686 -4840
rect 1652 -4930 1686 -4908
rect 1652 -5002 1686 -4976
rect 1652 -5074 1686 -5044
rect 1652 -5146 1686 -5112
rect 1652 -5214 1686 -5180
rect 1652 -5282 1686 -5252
rect 1652 -5350 1686 -5324
rect 1652 -5418 1686 -5396
rect 1652 -5486 1686 -5468
rect 1652 -5567 1686 -5540
rect 1748 -4786 1782 -4759
rect 1748 -4858 1782 -4840
rect 1748 -4930 1782 -4908
rect 1748 -5002 1782 -4976
rect 1748 -5074 1782 -5044
rect 1748 -5146 1782 -5112
rect 1748 -5214 1782 -5180
rect 1748 -5282 1782 -5252
rect 1748 -5350 1782 -5324
rect 1748 -5418 1782 -5396
rect 1748 -5486 1782 -5468
rect 1748 -5567 1782 -5540
rect 1844 -4786 1878 -4759
rect 1844 -4858 1878 -4840
rect 1844 -4930 1878 -4908
rect 1844 -5002 1878 -4976
rect 1844 -5074 1878 -5044
rect 1844 -5146 1878 -5112
rect 1844 -5214 1878 -5180
rect 1844 -5282 1878 -5252
rect 1844 -5350 1878 -5324
rect 1844 -5418 1878 -5396
rect 1844 -5486 1878 -5468
rect 1844 -5567 1878 -5540
rect 1940 -4786 1974 -4759
rect 1940 -4858 1974 -4840
rect 1940 -4930 1974 -4908
rect 1940 -5002 1974 -4976
rect 1940 -5074 1974 -5044
rect 1940 -5146 1974 -5112
rect 1940 -5214 1974 -5180
rect 1940 -5282 1974 -5252
rect 1940 -5350 1974 -5324
rect 1940 -5418 1974 -5396
rect 1940 -5486 1974 -5468
rect 1940 -5567 1974 -5540
rect -42834 -5603 -40735 -5591
rect -42902 -5607 -40735 -5603
rect -42902 -5641 -42441 -5607
rect -42407 -5641 -42369 -5607
rect -42335 -5641 -42297 -5607
rect -42263 -5641 -42225 -5607
rect -42191 -5641 -42153 -5607
rect -42119 -5641 -42081 -5607
rect -42047 -5641 -42009 -5607
rect -41975 -5641 -41937 -5607
rect -41903 -5641 -41865 -5607
rect -41831 -5641 -41793 -5607
rect -41759 -5641 -41721 -5607
rect -41687 -5641 -41649 -5607
rect -41615 -5641 -41577 -5607
rect -41543 -5641 -41505 -5607
rect -41471 -5641 -41433 -5607
rect -41399 -5641 -41361 -5607
rect -41327 -5641 -41289 -5607
rect -41255 -5641 -41217 -5607
rect -41183 -5641 -41145 -5607
rect -41111 -5641 -41073 -5607
rect -41039 -5641 -41001 -5607
rect -40967 -5641 -40929 -5607
rect -40895 -5641 -40857 -5607
rect -40823 -5641 -40785 -5607
rect -40751 -5641 -40735 -5607
rect -42902 -5679 -40735 -5641
rect -42902 -5713 -42441 -5679
rect -42407 -5713 -42369 -5679
rect -42335 -5713 -42297 -5679
rect -42263 -5713 -42225 -5679
rect -42191 -5713 -42153 -5679
rect -42119 -5713 -42081 -5679
rect -42047 -5713 -42009 -5679
rect -41975 -5713 -41937 -5679
rect -41903 -5713 -41865 -5679
rect -41831 -5713 -41793 -5679
rect -41759 -5713 -41721 -5679
rect -41687 -5713 -41649 -5679
rect -41615 -5713 -41577 -5679
rect -41543 -5713 -41505 -5679
rect -41471 -5713 -41433 -5679
rect -41399 -5713 -41361 -5679
rect -41327 -5713 -41289 -5679
rect -41255 -5713 -41217 -5679
rect -41183 -5713 -41145 -5679
rect -41111 -5713 -41073 -5679
rect -41039 -5713 -41001 -5679
rect -40967 -5713 -40929 -5679
rect -40895 -5713 -40857 -5679
rect -40823 -5713 -40785 -5679
rect -40751 -5713 -40735 -5679
rect -42902 -5729 -40735 -5713
rect 184 -5623 2404 -5617
rect 184 -5633 2472 -5623
rect 184 -5667 200 -5633
rect 234 -5667 272 -5633
rect 306 -5667 344 -5633
rect 378 -5667 416 -5633
rect 450 -5667 488 -5633
rect 522 -5667 560 -5633
rect 594 -5667 632 -5633
rect 666 -5667 704 -5633
rect 738 -5667 776 -5633
rect 810 -5667 848 -5633
rect 882 -5667 920 -5633
rect 954 -5667 992 -5633
rect 1026 -5667 1064 -5633
rect 1098 -5667 1136 -5633
rect 1170 -5667 1208 -5633
rect 1242 -5667 1280 -5633
rect 1314 -5667 1352 -5633
rect 1386 -5667 1424 -5633
rect 1458 -5667 1496 -5633
rect 1530 -5667 1568 -5633
rect 1602 -5667 1640 -5633
rect 1674 -5667 1712 -5633
rect 1746 -5667 1784 -5633
rect 1818 -5667 1856 -5633
rect 1890 -5667 2472 -5633
rect 184 -5705 2472 -5667
rect 184 -5739 200 -5705
rect 234 -5739 272 -5705
rect 306 -5739 344 -5705
rect 378 -5739 416 -5705
rect 450 -5739 488 -5705
rect 522 -5739 560 -5705
rect 594 -5739 632 -5705
rect 666 -5739 704 -5705
rect 738 -5739 776 -5705
rect 810 -5739 848 -5705
rect 882 -5739 920 -5705
rect 954 -5739 992 -5705
rect 1026 -5739 1064 -5705
rect 1098 -5739 1136 -5705
rect 1170 -5739 1208 -5705
rect 1242 -5739 1280 -5705
rect 1314 -5739 1352 -5705
rect 1386 -5739 1424 -5705
rect 1458 -5739 1496 -5705
rect 1530 -5739 1568 -5705
rect 1602 -5739 1640 -5705
rect 1674 -5739 1712 -5705
rect 1746 -5739 1784 -5705
rect 1818 -5739 1856 -5705
rect 1890 -5739 2472 -5705
rect 184 -5755 2472 -5739
<< viali >>
rect -50449 33490 -50415 33524
rect -50415 33490 -50377 33524
rect -50377 33490 -50343 33524
rect -50343 33490 -50305 33524
rect -50305 33490 -50271 33524
rect -50271 33490 -50233 33524
rect -50233 33490 -50199 33524
rect -50199 33490 -50161 33524
rect -50161 33490 -50127 33524
rect -50127 33490 -50089 33524
rect -50089 33490 -50055 33524
rect -50055 33490 -50017 33524
rect -50017 33490 -49983 33524
rect -49983 33490 -49945 33524
rect -49945 33490 -49911 33524
rect -49911 33490 -49873 33524
rect -49873 33490 -49839 33524
rect -49839 33490 -49801 33524
rect -49801 33490 -49767 33524
rect -49767 33490 -49729 33524
rect -49729 33490 -49695 33524
rect -49695 33490 -49657 33524
rect -49657 33490 -49623 33524
rect -49623 33490 -49585 33524
rect -49585 33490 -49551 33524
rect -49551 33490 -49513 33524
rect -49513 33490 -49479 33524
rect -49479 33490 -49441 33524
rect -49441 33490 -49407 33524
rect -49407 33490 -49369 33524
rect -49369 33490 -49335 33524
rect -49335 33490 -49297 33524
rect -49297 33490 -49263 33524
rect -49263 33490 -49225 33524
rect -49225 33490 -49191 33524
rect -49191 33490 -49153 33524
rect -49153 33490 -49119 33524
rect -49119 33490 -49081 33524
rect -49081 33490 -49047 33524
rect -49047 33490 -49009 33524
rect -49009 33490 -48975 33524
rect -48975 33490 -48937 33524
rect -48937 33490 -48903 33524
rect -48903 33490 -48865 33524
rect -48865 33490 -48831 33524
rect -50449 33452 -48831 33490
rect -50449 33418 -50415 33452
rect -50415 33418 -50377 33452
rect -50377 33418 -50343 33452
rect -50343 33418 -50305 33452
rect -50305 33418 -50271 33452
rect -50271 33418 -50233 33452
rect -50233 33418 -50199 33452
rect -50199 33418 -50161 33452
rect -50161 33418 -50127 33452
rect -50127 33418 -50089 33452
rect -50089 33418 -50055 33452
rect -50055 33418 -50017 33452
rect -50017 33418 -49983 33452
rect -49983 33418 -49945 33452
rect -49945 33418 -49911 33452
rect -49911 33418 -49873 33452
rect -49873 33418 -49839 33452
rect -49839 33418 -49801 33452
rect -49801 33418 -49767 33452
rect -49767 33418 -49729 33452
rect -49729 33418 -49695 33452
rect -49695 33418 -49657 33452
rect -49657 33418 -49623 33452
rect -49623 33418 -49585 33452
rect -49585 33418 -49551 33452
rect -49551 33418 -49513 33452
rect -49513 33418 -49479 33452
rect -49479 33418 -49441 33452
rect -49441 33418 -49407 33452
rect -49407 33418 -49369 33452
rect -49369 33418 -49335 33452
rect -49335 33418 -49297 33452
rect -49297 33418 -49263 33452
rect -49263 33418 -49225 33452
rect -49225 33418 -49191 33452
rect -49191 33418 -49153 33452
rect -49153 33418 -49119 33452
rect -49119 33418 -49081 33452
rect -49081 33418 -49047 33452
rect -49047 33418 -49009 33452
rect -49009 33418 -48975 33452
rect -48975 33418 -48937 33452
rect -48937 33418 -48903 33452
rect -48903 33418 -48865 33452
rect -48865 33418 -48831 33452
rect 2898 33490 2932 33524
rect 2932 33490 2970 33524
rect 2970 33490 3004 33524
rect 3004 33490 3042 33524
rect 3042 33490 3076 33524
rect 3076 33490 3114 33524
rect 3114 33490 3148 33524
rect 3148 33490 3186 33524
rect 3186 33490 3220 33524
rect 3220 33490 3258 33524
rect 3258 33490 3292 33524
rect 3292 33490 3330 33524
rect 3330 33490 3364 33524
rect 3364 33490 3402 33524
rect 3402 33490 3436 33524
rect 3436 33490 3474 33524
rect 3474 33490 3508 33524
rect 3508 33490 3546 33524
rect 3546 33490 3580 33524
rect 3580 33490 3618 33524
rect 3618 33490 3652 33524
rect 3652 33490 3690 33524
rect 3690 33490 3724 33524
rect 3724 33490 3762 33524
rect 3762 33490 3796 33524
rect 3796 33490 3834 33524
rect 3834 33490 3868 33524
rect 3868 33490 3906 33524
rect 3906 33490 3940 33524
rect 3940 33490 3978 33524
rect 3978 33490 4012 33524
rect 4012 33490 4050 33524
rect 4050 33490 4084 33524
rect 4084 33490 4122 33524
rect 4122 33490 4156 33524
rect 4156 33490 4194 33524
rect 4194 33490 4228 33524
rect 4228 33490 4266 33524
rect 4266 33490 4300 33524
rect 4300 33490 4338 33524
rect 4338 33490 4372 33524
rect 4372 33490 4410 33524
rect 4410 33490 4444 33524
rect 4444 33490 4482 33524
rect 4482 33490 4516 33524
rect 2898 33452 4516 33490
rect 2898 33418 2932 33452
rect 2932 33418 2970 33452
rect 2970 33418 3004 33452
rect 3004 33418 3042 33452
rect 3042 33418 3076 33452
rect 3076 33418 3114 33452
rect 3114 33418 3148 33452
rect 3148 33418 3186 33452
rect 3186 33418 3220 33452
rect 3220 33418 3258 33452
rect 3258 33418 3292 33452
rect 3292 33418 3330 33452
rect 3330 33418 3364 33452
rect 3364 33418 3402 33452
rect 3402 33418 3436 33452
rect 3436 33418 3474 33452
rect 3474 33418 3508 33452
rect 3508 33418 3546 33452
rect 3546 33418 3580 33452
rect 3580 33418 3618 33452
rect 3618 33418 3652 33452
rect 3652 33418 3690 33452
rect 3690 33418 3724 33452
rect 3724 33418 3762 33452
rect 3762 33418 3796 33452
rect 3796 33418 3834 33452
rect 3834 33418 3868 33452
rect 3868 33418 3906 33452
rect 3906 33418 3940 33452
rect 3940 33418 3978 33452
rect 3978 33418 4012 33452
rect 4012 33418 4050 33452
rect 4050 33418 4084 33452
rect 4084 33418 4122 33452
rect 4122 33418 4156 33452
rect 4156 33418 4194 33452
rect 4194 33418 4228 33452
rect 4228 33418 4266 33452
rect 4266 33418 4300 33452
rect 4300 33418 4338 33452
rect 4338 33418 4372 33452
rect 4372 33418 4410 33452
rect 4410 33418 4444 33452
rect 4444 33418 4482 33452
rect 4482 33418 4516 33452
rect -50447 33265 -50413 33273
rect -50447 33239 -50413 33265
rect -50447 33197 -50413 33201
rect -50447 33167 -50413 33197
rect -50447 33095 -50413 33129
rect -50447 33027 -50413 33057
rect -50447 33023 -50413 33027
rect -50447 32959 -50413 32985
rect -50926 32618 -50604 32940
rect -50447 32951 -50413 32959
rect -50289 33265 -50255 33273
rect -50289 33239 -50255 33265
rect -50289 33197 -50255 33201
rect -50289 33167 -50255 33197
rect -50289 33095 -50255 33129
rect -50289 33027 -50255 33057
rect -50289 33023 -50255 33027
rect -50289 32959 -50255 32985
rect -50289 32951 -50255 32959
rect -50131 33265 -50097 33273
rect -50131 33239 -50097 33265
rect -50131 33197 -50097 33201
rect -50131 33167 -50097 33197
rect -50131 33095 -50097 33129
rect -50131 33027 -50097 33057
rect -50131 33023 -50097 33027
rect -50131 32959 -50097 32985
rect -50131 32951 -50097 32959
rect -49973 33265 -49939 33273
rect -49973 33239 -49939 33265
rect -49973 33197 -49939 33201
rect -49973 33167 -49939 33197
rect -49973 33095 -49939 33129
rect -49973 33027 -49939 33057
rect -49973 33023 -49939 33027
rect -49973 32959 -49939 32985
rect -49973 32951 -49939 32959
rect -49815 33265 -49781 33273
rect -49815 33239 -49781 33265
rect -49815 33197 -49781 33201
rect -49815 33167 -49781 33197
rect -49815 33095 -49781 33129
rect -49815 33027 -49781 33057
rect -49815 33023 -49781 33027
rect -49815 32959 -49781 32985
rect -49815 32951 -49781 32959
rect -49657 33265 -49623 33273
rect -49657 33239 -49623 33265
rect -49657 33197 -49623 33201
rect -49657 33167 -49623 33197
rect -49657 33095 -49623 33129
rect -49657 33027 -49623 33057
rect -49657 33023 -49623 33027
rect -49657 32959 -49623 32985
rect -49657 32951 -49623 32959
rect -49499 33265 -49465 33273
rect -49499 33239 -49465 33265
rect -49499 33197 -49465 33201
rect -49499 33167 -49465 33197
rect -49499 33095 -49465 33129
rect -49499 33027 -49465 33057
rect -49499 33023 -49465 33027
rect -49499 32959 -49465 32985
rect -49499 32951 -49465 32959
rect -49341 33265 -49307 33273
rect -49341 33239 -49307 33265
rect -49341 33197 -49307 33201
rect -49341 33167 -49307 33197
rect -49341 33095 -49307 33129
rect -49341 33027 -49307 33057
rect -49341 33023 -49307 33027
rect -49341 32959 -49307 32985
rect -49341 32951 -49307 32959
rect -49183 33265 -49149 33273
rect -49183 33239 -49149 33265
rect -49183 33197 -49149 33201
rect -49183 33167 -49149 33197
rect -49183 33095 -49149 33129
rect -49183 33027 -49149 33057
rect -49183 33023 -49149 33027
rect -49183 32959 -49149 32985
rect -49183 32951 -49149 32959
rect -49025 33265 -48991 33273
rect -49025 33239 -48991 33265
rect -49025 33197 -48991 33201
rect -49025 33167 -48991 33197
rect -49025 33095 -48991 33129
rect -49025 33027 -48991 33057
rect -49025 33023 -48991 33027
rect -49025 32959 -48991 32985
rect -49025 32951 -48991 32959
rect -48867 33265 -48833 33273
rect -48867 33239 -48833 33265
rect -48867 33197 -48833 33201
rect -48867 33167 -48833 33197
rect -48867 33095 -48833 33129
rect -48867 33027 -48833 33057
rect -48867 33023 -48833 33027
rect -48867 32959 -48833 32985
rect -48867 32951 -48833 32959
rect 2900 33265 2934 33273
rect 2900 33239 2934 33265
rect 2900 33197 2934 33201
rect 2900 33167 2934 33197
rect 2900 33095 2934 33129
rect 2900 33027 2934 33057
rect 2900 33023 2934 33027
rect 2900 32959 2934 32985
rect -50368 32831 -50334 32865
rect -50210 32831 -50176 32865
rect -50052 32831 -50018 32865
rect -49894 32831 -49860 32865
rect -49736 32831 -49702 32865
rect -49578 32831 -49544 32865
rect -49420 32831 -49386 32865
rect -49262 32831 -49228 32865
rect -49104 32831 -49070 32865
rect -48946 32831 -48912 32865
rect -50368 32693 -50334 32727
rect -50210 32693 -50176 32727
rect -50052 32693 -50018 32727
rect -49894 32693 -49860 32727
rect -49736 32693 -49702 32727
rect -49578 32693 -49544 32727
rect -49420 32693 -49386 32727
rect -49262 32693 -49228 32727
rect -49104 32693 -49070 32727
rect -48946 32693 -48912 32727
rect -50447 32606 -50413 32608
rect -50447 32574 -50413 32606
rect -50447 32504 -50413 32536
rect -50447 32502 -50413 32504
rect -50289 32606 -50255 32608
rect -50289 32574 -50255 32606
rect -50289 32504 -50255 32536
rect -50289 32502 -50255 32504
rect -50131 32606 -50097 32608
rect -50131 32574 -50097 32606
rect -50131 32504 -50097 32536
rect -50131 32502 -50097 32504
rect -49973 32606 -49939 32608
rect -49973 32574 -49939 32606
rect -49973 32504 -49939 32536
rect -49973 32502 -49939 32504
rect -49815 32606 -49781 32608
rect -49815 32574 -49781 32606
rect -49815 32504 -49781 32536
rect -49815 32502 -49781 32504
rect -49657 32606 -49623 32608
rect -49657 32574 -49623 32606
rect -49657 32504 -49623 32536
rect -49657 32502 -49623 32504
rect -49499 32606 -49465 32608
rect -49499 32574 -49465 32606
rect -49499 32504 -49465 32536
rect -49499 32502 -49465 32504
rect -49341 32606 -49307 32608
rect -49341 32574 -49307 32606
rect -49341 32504 -49307 32536
rect -49341 32502 -49307 32504
rect -49183 32606 -49149 32608
rect -49183 32574 -49149 32606
rect -49183 32504 -49149 32536
rect -49183 32502 -49149 32504
rect -49025 32606 -48991 32608
rect -49025 32574 -48991 32606
rect -49025 32504 -48991 32536
rect -49025 32502 -48991 32504
rect -48867 32606 -48833 32608
rect -48867 32574 -48833 32606
rect -48867 32504 -48833 32536
rect -48867 32502 -48833 32504
rect 2421 32618 2743 32940
rect 2900 32951 2934 32959
rect 3058 33265 3092 33273
rect 3058 33239 3092 33265
rect 3058 33197 3092 33201
rect 3058 33167 3092 33197
rect 3058 33095 3092 33129
rect 3058 33027 3092 33057
rect 3058 33023 3092 33027
rect 3058 32959 3092 32985
rect 3058 32951 3092 32959
rect 3216 33265 3250 33273
rect 3216 33239 3250 33265
rect 3216 33197 3250 33201
rect 3216 33167 3250 33197
rect 3216 33095 3250 33129
rect 3216 33027 3250 33057
rect 3216 33023 3250 33027
rect 3216 32959 3250 32985
rect 3216 32951 3250 32959
rect 3374 33265 3408 33273
rect 3374 33239 3408 33265
rect 3374 33197 3408 33201
rect 3374 33167 3408 33197
rect 3374 33095 3408 33129
rect 3374 33027 3408 33057
rect 3374 33023 3408 33027
rect 3374 32959 3408 32985
rect 3374 32951 3408 32959
rect 3532 33265 3566 33273
rect 3532 33239 3566 33265
rect 3532 33197 3566 33201
rect 3532 33167 3566 33197
rect 3532 33095 3566 33129
rect 3532 33027 3566 33057
rect 3532 33023 3566 33027
rect 3532 32959 3566 32985
rect 3532 32951 3566 32959
rect 3690 33265 3724 33273
rect 3690 33239 3724 33265
rect 3690 33197 3724 33201
rect 3690 33167 3724 33197
rect 3690 33095 3724 33129
rect 3690 33027 3724 33057
rect 3690 33023 3724 33027
rect 3690 32959 3724 32985
rect 3690 32951 3724 32959
rect 3848 33265 3882 33273
rect 3848 33239 3882 33265
rect 3848 33197 3882 33201
rect 3848 33167 3882 33197
rect 3848 33095 3882 33129
rect 3848 33027 3882 33057
rect 3848 33023 3882 33027
rect 3848 32959 3882 32985
rect 3848 32951 3882 32959
rect 4006 33265 4040 33273
rect 4006 33239 4040 33265
rect 4006 33197 4040 33201
rect 4006 33167 4040 33197
rect 4006 33095 4040 33129
rect 4006 33027 4040 33057
rect 4006 33023 4040 33027
rect 4006 32959 4040 32985
rect 4006 32951 4040 32959
rect 4164 33265 4198 33273
rect 4164 33239 4198 33265
rect 4164 33197 4198 33201
rect 4164 33167 4198 33197
rect 4164 33095 4198 33129
rect 4164 33027 4198 33057
rect 4164 33023 4198 33027
rect 4164 32959 4198 32985
rect 4164 32951 4198 32959
rect 4322 33265 4356 33273
rect 4322 33239 4356 33265
rect 4322 33197 4356 33201
rect 4322 33167 4356 33197
rect 4322 33095 4356 33129
rect 4322 33027 4356 33057
rect 4322 33023 4356 33027
rect 4322 32959 4356 32985
rect 4322 32951 4356 32959
rect 4480 33265 4514 33273
rect 4480 33239 4514 33265
rect 4480 33197 4514 33201
rect 4480 33167 4514 33197
rect 4480 33095 4514 33129
rect 4480 33027 4514 33057
rect 4480 33023 4514 33027
rect 4480 32959 4514 32985
rect 4480 32951 4514 32959
rect 2979 32831 3013 32865
rect 3137 32831 3171 32865
rect 3295 32831 3329 32865
rect 3453 32831 3487 32865
rect 3611 32831 3645 32865
rect 3769 32831 3803 32865
rect 3927 32831 3961 32865
rect 4085 32831 4119 32865
rect 4243 32831 4277 32865
rect 4401 32831 4435 32865
rect 2979 32693 3013 32727
rect 3137 32693 3171 32727
rect 3295 32693 3329 32727
rect 3453 32693 3487 32727
rect 3611 32693 3645 32727
rect 3769 32693 3803 32727
rect 3927 32693 3961 32727
rect 4085 32693 4119 32727
rect 4243 32693 4277 32727
rect 4401 32693 4435 32727
rect 2900 32606 2934 32608
rect 2153 32505 2187 32539
rect 2900 32574 2934 32606
rect 2900 32504 2934 32536
rect 2900 32502 2934 32504
rect 3058 32606 3092 32608
rect 3058 32574 3092 32606
rect 3058 32504 3092 32536
rect 3058 32502 3092 32504
rect 3216 32606 3250 32608
rect 3216 32574 3250 32606
rect 3216 32504 3250 32536
rect 3216 32502 3250 32504
rect 3374 32606 3408 32608
rect 3374 32574 3408 32606
rect 3374 32504 3408 32536
rect 3374 32502 3408 32504
rect 3532 32606 3566 32608
rect 3532 32574 3566 32606
rect 3532 32504 3566 32536
rect 3532 32502 3566 32504
rect 3690 32606 3724 32608
rect 3690 32574 3724 32606
rect 3690 32504 3724 32536
rect 3690 32502 3724 32504
rect 3848 32606 3882 32608
rect 3848 32574 3882 32606
rect 3848 32504 3882 32536
rect 3848 32502 3882 32504
rect 4006 32606 4040 32608
rect 4006 32574 4040 32606
rect 4006 32504 4040 32536
rect 4006 32502 4040 32504
rect 4164 32606 4198 32608
rect 4164 32574 4198 32606
rect 4164 32504 4198 32536
rect 4164 32502 4198 32504
rect 4322 32606 4356 32608
rect 4322 32574 4356 32606
rect 4322 32504 4356 32536
rect 4322 32502 4356 32504
rect 4480 32606 4514 32608
rect 4480 32574 4514 32606
rect 4480 32504 4514 32536
rect 4480 32502 4514 32504
rect -50449 32315 -50415 32349
rect -50415 32315 -50377 32349
rect -50377 32315 -50343 32349
rect -50343 32315 -50305 32349
rect -50305 32315 -50271 32349
rect -50271 32315 -50233 32349
rect -50233 32315 -50199 32349
rect -50199 32315 -50161 32349
rect -50161 32315 -50127 32349
rect -50127 32315 -50089 32349
rect -50089 32315 -50055 32349
rect -50055 32315 -50017 32349
rect -50017 32315 -49983 32349
rect -49983 32315 -49945 32349
rect -49945 32315 -49911 32349
rect -49911 32315 -49873 32349
rect -49873 32315 -49839 32349
rect -49839 32315 -49801 32349
rect -49801 32315 -49767 32349
rect -49767 32315 -49729 32349
rect -49729 32315 -49695 32349
rect -49695 32315 -49657 32349
rect -49657 32315 -49623 32349
rect -49623 32315 -49585 32349
rect -49585 32315 -49551 32349
rect -49551 32315 -49513 32349
rect -49513 32315 -49479 32349
rect -49479 32315 -49441 32349
rect -49441 32315 -49407 32349
rect -49407 32315 -49369 32349
rect -49369 32315 -49335 32349
rect -49335 32315 -49297 32349
rect -49297 32315 -49263 32349
rect -49263 32315 -49225 32349
rect -49225 32315 -49191 32349
rect -49191 32315 -49153 32349
rect -49153 32315 -49119 32349
rect -49119 32315 -49081 32349
rect -49081 32315 -49047 32349
rect -49047 32315 -49009 32349
rect -49009 32315 -48975 32349
rect -48975 32315 -48937 32349
rect -48937 32315 -48903 32349
rect -48903 32315 -48865 32349
rect -48865 32315 -48831 32349
rect -50449 32277 -48831 32315
rect -50449 32243 -50415 32277
rect -50415 32243 -50377 32277
rect -50377 32243 -50343 32277
rect -50343 32243 -50305 32277
rect -50305 32243 -50271 32277
rect -50271 32243 -50233 32277
rect -50233 32243 -50199 32277
rect -50199 32243 -50161 32277
rect -50161 32243 -50127 32277
rect -50127 32243 -50089 32277
rect -50089 32243 -50055 32277
rect -50055 32243 -50017 32277
rect -50017 32243 -49983 32277
rect -49983 32243 -49945 32277
rect -49945 32243 -49911 32277
rect -49911 32243 -49873 32277
rect -49873 32243 -49839 32277
rect -49839 32243 -49801 32277
rect -49801 32243 -49767 32277
rect -49767 32243 -49729 32277
rect -49729 32243 -49695 32277
rect -49695 32243 -49657 32277
rect -49657 32243 -49623 32277
rect -49623 32243 -49585 32277
rect -49585 32243 -49551 32277
rect -49551 32243 -49513 32277
rect -49513 32243 -49479 32277
rect -49479 32243 -49441 32277
rect -49441 32243 -49407 32277
rect -49407 32243 -49369 32277
rect -49369 32243 -49335 32277
rect -49335 32243 -49297 32277
rect -49297 32243 -49263 32277
rect -49263 32243 -49225 32277
rect -49225 32243 -49191 32277
rect -49191 32243 -49153 32277
rect -49153 32243 -49119 32277
rect -49119 32243 -49081 32277
rect -49081 32243 -49047 32277
rect -49047 32243 -49009 32277
rect -49009 32243 -48975 32277
rect -48975 32243 -48937 32277
rect -48937 32243 -48903 32277
rect -48903 32243 -48865 32277
rect -48865 32243 -48831 32277
rect 1979 32253 2301 32359
rect 2898 32315 2932 32349
rect 2932 32315 2970 32349
rect 2970 32315 3004 32349
rect 3004 32315 3042 32349
rect 3042 32315 3076 32349
rect 3076 32315 3114 32349
rect 3114 32315 3148 32349
rect 3148 32315 3186 32349
rect 3186 32315 3220 32349
rect 3220 32315 3258 32349
rect 3258 32315 3292 32349
rect 3292 32315 3330 32349
rect 3330 32315 3364 32349
rect 3364 32315 3402 32349
rect 3402 32315 3436 32349
rect 3436 32315 3474 32349
rect 3474 32315 3508 32349
rect 3508 32315 3546 32349
rect 3546 32315 3580 32349
rect 3580 32315 3618 32349
rect 3618 32315 3652 32349
rect 3652 32315 3690 32349
rect 3690 32315 3724 32349
rect 3724 32315 3762 32349
rect 3762 32315 3796 32349
rect 3796 32315 3834 32349
rect 3834 32315 3868 32349
rect 3868 32315 3906 32349
rect 3906 32315 3940 32349
rect 3940 32315 3978 32349
rect 3978 32315 4012 32349
rect 4012 32315 4050 32349
rect 4050 32315 4084 32349
rect 4084 32315 4122 32349
rect 4122 32315 4156 32349
rect 4156 32315 4194 32349
rect 4194 32315 4228 32349
rect 4228 32315 4266 32349
rect 4266 32315 4300 32349
rect 4300 32315 4338 32349
rect 4338 32315 4372 32349
rect 4372 32315 4410 32349
rect 4410 32315 4444 32349
rect 4444 32315 4482 32349
rect 4482 32315 4516 32349
rect 2898 32277 4516 32315
rect 2898 32243 2932 32277
rect 2932 32243 2970 32277
rect 2970 32243 3004 32277
rect 3004 32243 3042 32277
rect 3042 32243 3076 32277
rect 3076 32243 3114 32277
rect 3114 32243 3148 32277
rect 3148 32243 3186 32277
rect 3186 32243 3220 32277
rect 3220 32243 3258 32277
rect 3258 32243 3292 32277
rect 3292 32243 3330 32277
rect 3330 32243 3364 32277
rect 3364 32243 3402 32277
rect 3402 32243 3436 32277
rect 3436 32243 3474 32277
rect 3474 32243 3508 32277
rect 3508 32243 3546 32277
rect 3546 32243 3580 32277
rect 3580 32243 3618 32277
rect 3618 32243 3652 32277
rect 3652 32243 3690 32277
rect 3690 32243 3724 32277
rect 3724 32243 3762 32277
rect 3762 32243 3796 32277
rect 3796 32243 3834 32277
rect 3834 32243 3868 32277
rect 3868 32243 3906 32277
rect 3906 32243 3940 32277
rect 3940 32243 3978 32277
rect 3978 32243 4012 32277
rect 4012 32243 4050 32277
rect 4050 32243 4084 32277
rect 4084 32243 4122 32277
rect 4122 32243 4156 32277
rect 4156 32243 4194 32277
rect 4194 32243 4228 32277
rect 4228 32243 4266 32277
rect 4266 32243 4300 32277
rect 4300 32243 4338 32277
rect 4338 32243 4372 32277
rect 4372 32243 4410 32277
rect 4410 32243 4444 32277
rect 4444 32243 4482 32277
rect 4482 32243 4516 32277
rect -50769 32001 -50735 32035
rect -50589 31827 -50483 32149
rect -47340 24954 -47306 24973
rect -47340 24939 -47306 24954
rect -47340 24867 -47306 24901
rect -47340 24795 -47306 24829
rect -47340 24723 -47306 24757
rect 6874 24919 6908 24953
rect 6874 24847 6908 24881
rect 6874 24775 6908 24809
rect 6874 24703 6908 24737
rect -42524 5394 -42490 5414
rect -42524 5380 -42490 5394
rect -42524 5326 -42490 5342
rect -42524 5308 -42490 5326
rect -42524 5258 -42490 5270
rect -42524 5236 -42490 5258
rect -42524 5190 -42490 5198
rect -42524 5164 -42490 5190
rect -42524 5122 -42490 5126
rect -42524 5092 -42490 5122
rect -42524 5020 -42490 5054
rect -42524 4952 -42490 4982
rect -42524 4948 -42490 4952
rect -42524 4884 -42490 4910
rect -42524 4876 -42490 4884
rect -42524 4816 -42490 4838
rect -42524 4804 -42490 4816
rect -42524 4748 -42490 4766
rect -42524 4732 -42490 4748
rect -42524 4680 -42490 4694
rect -42524 4660 -42490 4680
rect -42428 5394 -42394 5414
rect -42428 5380 -42394 5394
rect -42428 5326 -42394 5342
rect -42428 5308 -42394 5326
rect -42428 5258 -42394 5270
rect -42428 5236 -42394 5258
rect -42428 5190 -42394 5198
rect -42428 5164 -42394 5190
rect -42428 5122 -42394 5126
rect -42428 5092 -42394 5122
rect -42428 5020 -42394 5054
rect -42428 4952 -42394 4982
rect -42428 4948 -42394 4952
rect -42428 4884 -42394 4910
rect -42428 4876 -42394 4884
rect -42428 4816 -42394 4838
rect -42428 4804 -42394 4816
rect -42428 4748 -42394 4766
rect -42428 4732 -42394 4748
rect -42428 4680 -42394 4694
rect -42428 4660 -42394 4680
rect -42332 5394 -42298 5414
rect -42332 5380 -42298 5394
rect -42332 5326 -42298 5342
rect -42332 5308 -42298 5326
rect -42332 5258 -42298 5270
rect -42332 5236 -42298 5258
rect -42332 5190 -42298 5198
rect -42332 5164 -42298 5190
rect -42332 5122 -42298 5126
rect -42332 5092 -42298 5122
rect -42332 5020 -42298 5054
rect -42332 4952 -42298 4982
rect -42332 4948 -42298 4952
rect -42332 4884 -42298 4910
rect -42332 4876 -42298 4884
rect -42332 4816 -42298 4838
rect -42332 4804 -42298 4816
rect -42332 4748 -42298 4766
rect -42332 4732 -42298 4748
rect -42332 4680 -42298 4694
rect -42332 4660 -42298 4680
rect -42236 5394 -42202 5414
rect -42236 5380 -42202 5394
rect -42236 5326 -42202 5342
rect -42236 5308 -42202 5326
rect -42236 5258 -42202 5270
rect -42236 5236 -42202 5258
rect -42236 5190 -42202 5198
rect -42236 5164 -42202 5190
rect -42236 5122 -42202 5126
rect -42236 5092 -42202 5122
rect -42236 5020 -42202 5054
rect -42236 4952 -42202 4982
rect -42236 4948 -42202 4952
rect -42236 4884 -42202 4910
rect -42236 4876 -42202 4884
rect -42236 4816 -42202 4838
rect -42236 4804 -42202 4816
rect -42236 4748 -42202 4766
rect -42236 4732 -42202 4748
rect -42236 4680 -42202 4694
rect -42236 4660 -42202 4680
rect -42140 5394 -42106 5414
rect -42140 5380 -42106 5394
rect -42140 5326 -42106 5342
rect -42140 5308 -42106 5326
rect -42140 5258 -42106 5270
rect -42140 5236 -42106 5258
rect -42140 5190 -42106 5198
rect -42140 5164 -42106 5190
rect -42140 5122 -42106 5126
rect -42140 5092 -42106 5122
rect -42140 5020 -42106 5054
rect -42140 4952 -42106 4982
rect -42140 4948 -42106 4952
rect -42140 4884 -42106 4910
rect -42140 4876 -42106 4884
rect -42140 4816 -42106 4838
rect -42140 4804 -42106 4816
rect -42140 4748 -42106 4766
rect -42140 4732 -42106 4748
rect -42140 4680 -42106 4694
rect -42140 4660 -42106 4680
rect -42044 5394 -42010 5414
rect -42044 5380 -42010 5394
rect -42044 5326 -42010 5342
rect -42044 5308 -42010 5326
rect -42044 5258 -42010 5270
rect -42044 5236 -42010 5258
rect -42044 5190 -42010 5198
rect -42044 5164 -42010 5190
rect -42044 5122 -42010 5126
rect -42044 5092 -42010 5122
rect -42044 5020 -42010 5054
rect -42044 4952 -42010 4982
rect -42044 4948 -42010 4952
rect -42044 4884 -42010 4910
rect -42044 4876 -42010 4884
rect -42044 4816 -42010 4838
rect -42044 4804 -42010 4816
rect -42044 4748 -42010 4766
rect -42044 4732 -42010 4748
rect -42044 4680 -42010 4694
rect -42044 4660 -42010 4680
rect -41948 5394 -41914 5414
rect -41948 5380 -41914 5394
rect -41948 5326 -41914 5342
rect -41948 5308 -41914 5326
rect -41948 5258 -41914 5270
rect -41948 5236 -41914 5258
rect -41948 5190 -41914 5198
rect -41948 5164 -41914 5190
rect -41948 5122 -41914 5126
rect -41948 5092 -41914 5122
rect -41948 5020 -41914 5054
rect -41948 4952 -41914 4982
rect -41948 4948 -41914 4952
rect -41948 4884 -41914 4910
rect -41948 4876 -41914 4884
rect -41948 4816 -41914 4838
rect -41948 4804 -41914 4816
rect -41948 4748 -41914 4766
rect -41948 4732 -41914 4748
rect -41948 4680 -41914 4694
rect -41948 4660 -41914 4680
rect -41852 5394 -41818 5414
rect -41852 5380 -41818 5394
rect -41852 5326 -41818 5342
rect -41852 5308 -41818 5326
rect -41852 5258 -41818 5270
rect -41852 5236 -41818 5258
rect -41852 5190 -41818 5198
rect -41852 5164 -41818 5190
rect -41852 5122 -41818 5126
rect -41852 5092 -41818 5122
rect -41852 5020 -41818 5054
rect -41852 4952 -41818 4982
rect -41852 4948 -41818 4952
rect -41852 4884 -41818 4910
rect -41852 4876 -41818 4884
rect -41852 4816 -41818 4838
rect -41852 4804 -41818 4816
rect -41852 4748 -41818 4766
rect -41852 4732 -41818 4748
rect -41852 4680 -41818 4694
rect -41852 4660 -41818 4680
rect -41756 5394 -41722 5414
rect -41756 5380 -41722 5394
rect -41756 5326 -41722 5342
rect -41756 5308 -41722 5326
rect -41756 5258 -41722 5270
rect -41756 5236 -41722 5258
rect -41756 5190 -41722 5198
rect -41756 5164 -41722 5190
rect -41756 5122 -41722 5126
rect -41756 5092 -41722 5122
rect -41756 5020 -41722 5054
rect -41756 4952 -41722 4982
rect -41756 4948 -41722 4952
rect -41756 4884 -41722 4910
rect -41756 4876 -41722 4884
rect -41756 4816 -41722 4838
rect -41756 4804 -41722 4816
rect -41756 4748 -41722 4766
rect -41756 4732 -41722 4748
rect -41756 4680 -41722 4694
rect -41756 4660 -41722 4680
rect -41660 5394 -41626 5414
rect -41660 5380 -41626 5394
rect -41660 5326 -41626 5342
rect -41660 5308 -41626 5326
rect -41660 5258 -41626 5270
rect -41660 5236 -41626 5258
rect -41660 5190 -41626 5198
rect -41660 5164 -41626 5190
rect -41660 5122 -41626 5126
rect -41660 5092 -41626 5122
rect -41660 5020 -41626 5054
rect -41660 4952 -41626 4982
rect -41660 4948 -41626 4952
rect -41660 4884 -41626 4910
rect -41660 4876 -41626 4884
rect -41660 4816 -41626 4838
rect -41660 4804 -41626 4816
rect -41660 4748 -41626 4766
rect -41660 4732 -41626 4748
rect -41660 4680 -41626 4694
rect -41660 4660 -41626 4680
rect -41564 5394 -41530 5414
rect -41564 5380 -41530 5394
rect -41564 5326 -41530 5342
rect -41564 5308 -41530 5326
rect -41564 5258 -41530 5270
rect -41564 5236 -41530 5258
rect -41564 5190 -41530 5198
rect -41564 5164 -41530 5190
rect -41564 5122 -41530 5126
rect -41564 5092 -41530 5122
rect -41564 5020 -41530 5054
rect -41564 4952 -41530 4982
rect -41564 4948 -41530 4952
rect -41564 4884 -41530 4910
rect -41564 4876 -41530 4884
rect -41564 4816 -41530 4838
rect -41564 4804 -41530 4816
rect -41564 4748 -41530 4766
rect -41564 4732 -41530 4748
rect -41564 4680 -41530 4694
rect -41564 4660 -41530 4680
rect -41468 5394 -41434 5414
rect -41468 5380 -41434 5394
rect -41468 5326 -41434 5342
rect -41468 5308 -41434 5326
rect -41468 5258 -41434 5270
rect -41468 5236 -41434 5258
rect -41468 5190 -41434 5198
rect -41468 5164 -41434 5190
rect -41468 5122 -41434 5126
rect -41468 5092 -41434 5122
rect -41468 5020 -41434 5054
rect -41468 4952 -41434 4982
rect -41468 4948 -41434 4952
rect -41468 4884 -41434 4910
rect -41468 4876 -41434 4884
rect -41468 4816 -41434 4838
rect -41468 4804 -41434 4816
rect -41468 4748 -41434 4766
rect -41468 4732 -41434 4748
rect -41468 4680 -41434 4694
rect -41468 4660 -41434 4680
rect -41372 5394 -41338 5414
rect -41372 5380 -41338 5394
rect -41372 5326 -41338 5342
rect -41372 5308 -41338 5326
rect -41372 5258 -41338 5270
rect -41372 5236 -41338 5258
rect -41372 5190 -41338 5198
rect -41372 5164 -41338 5190
rect -41372 5122 -41338 5126
rect -41372 5092 -41338 5122
rect -41372 5020 -41338 5054
rect -41372 4952 -41338 4982
rect -41372 4948 -41338 4952
rect -41372 4884 -41338 4910
rect -41372 4876 -41338 4884
rect -41372 4816 -41338 4838
rect -41372 4804 -41338 4816
rect -41372 4748 -41338 4766
rect -41372 4732 -41338 4748
rect -41372 4680 -41338 4694
rect -41372 4660 -41338 4680
rect -41276 5394 -41242 5414
rect -41276 5380 -41242 5394
rect -41276 5326 -41242 5342
rect -41276 5308 -41242 5326
rect -41276 5258 -41242 5270
rect -41276 5236 -41242 5258
rect -41276 5190 -41242 5198
rect -41276 5164 -41242 5190
rect -41276 5122 -41242 5126
rect -41276 5092 -41242 5122
rect -41276 5020 -41242 5054
rect -41276 4952 -41242 4982
rect -41276 4948 -41242 4952
rect -41276 4884 -41242 4910
rect -41276 4876 -41242 4884
rect -41276 4816 -41242 4838
rect -41276 4804 -41242 4816
rect -41276 4748 -41242 4766
rect -41276 4732 -41242 4748
rect -41276 4680 -41242 4694
rect -41276 4660 -41242 4680
rect -41180 5394 -41146 5414
rect -41180 5380 -41146 5394
rect -41180 5326 -41146 5342
rect -41180 5308 -41146 5326
rect -41180 5258 -41146 5270
rect -41180 5236 -41146 5258
rect -41180 5190 -41146 5198
rect -41180 5164 -41146 5190
rect -41180 5122 -41146 5126
rect -41180 5092 -41146 5122
rect -41180 5020 -41146 5054
rect -41180 4952 -41146 4982
rect -41180 4948 -41146 4952
rect -41180 4884 -41146 4910
rect -41180 4876 -41146 4884
rect -41180 4816 -41146 4838
rect -41180 4804 -41146 4816
rect -41180 4748 -41146 4766
rect -41180 4732 -41146 4748
rect -41180 4680 -41146 4694
rect -41180 4660 -41146 4680
rect -41084 5394 -41050 5414
rect -41084 5380 -41050 5394
rect -41084 5326 -41050 5342
rect -41084 5308 -41050 5326
rect -41084 5258 -41050 5270
rect -41084 5236 -41050 5258
rect -41084 5190 -41050 5198
rect -41084 5164 -41050 5190
rect -41084 5122 -41050 5126
rect -41084 5092 -41050 5122
rect -41084 5020 -41050 5054
rect -41084 4952 -41050 4982
rect -41084 4948 -41050 4952
rect -41084 4884 -41050 4910
rect -41084 4876 -41050 4884
rect -41084 4816 -41050 4838
rect -41084 4804 -41050 4816
rect -41084 4748 -41050 4766
rect -41084 4732 -41050 4748
rect -41084 4680 -41050 4694
rect -41084 4660 -41050 4680
rect -40988 5394 -40954 5414
rect -40988 5380 -40954 5394
rect -40988 5326 -40954 5342
rect -40988 5308 -40954 5326
rect -40988 5258 -40954 5270
rect -40988 5236 -40954 5258
rect -40988 5190 -40954 5198
rect -40988 5164 -40954 5190
rect -40988 5122 -40954 5126
rect -40988 5092 -40954 5122
rect -40988 5020 -40954 5054
rect -40988 4952 -40954 4982
rect -40988 4948 -40954 4952
rect -40988 4884 -40954 4910
rect -40988 4876 -40954 4884
rect -40988 4816 -40954 4838
rect -40988 4804 -40954 4816
rect -40988 4748 -40954 4766
rect -40988 4732 -40954 4748
rect -40988 4680 -40954 4694
rect -40988 4660 -40954 4680
rect -40892 5394 -40858 5414
rect -40892 5380 -40858 5394
rect -40892 5326 -40858 5342
rect -40892 5308 -40858 5326
rect -40892 5258 -40858 5270
rect -40892 5236 -40858 5258
rect -40892 5190 -40858 5198
rect -40892 5164 -40858 5190
rect -40892 5122 -40858 5126
rect -40892 5092 -40858 5122
rect -40892 5020 -40858 5054
rect -40892 4952 -40858 4982
rect -40892 4948 -40858 4952
rect -40892 4884 -40858 4910
rect -40892 4876 -40858 4884
rect -40892 4816 -40858 4838
rect -40892 4804 -40858 4816
rect -40892 4748 -40858 4766
rect -40892 4732 -40858 4748
rect -40892 4680 -40858 4694
rect -40892 4660 -40858 4680
rect -40796 5394 -40762 5414
rect -40796 5380 -40762 5394
rect -40796 5326 -40762 5342
rect -40796 5308 -40762 5326
rect -40796 5258 -40762 5270
rect -40796 5236 -40762 5258
rect -40796 5190 -40762 5198
rect -40796 5164 -40762 5190
rect -40796 5122 -40762 5126
rect -40796 5092 -40762 5122
rect -40796 5020 -40762 5054
rect -40796 4952 -40762 4982
rect -40796 4948 -40762 4952
rect -40796 4884 -40762 4910
rect -40796 4876 -40762 4884
rect -40796 4816 -40762 4838
rect -40796 4804 -40762 4816
rect -40796 4748 -40762 4766
rect -40796 4732 -40762 4748
rect -40796 4680 -40762 4694
rect -40796 4660 -40762 4680
rect -40700 5394 -40666 5414
rect -40700 5380 -40666 5394
rect -40700 5326 -40666 5342
rect -40700 5308 -40666 5326
rect -40700 5258 -40666 5270
rect -40700 5236 -40666 5258
rect -40700 5190 -40666 5198
rect -40700 5164 -40666 5190
rect -40700 5122 -40666 5126
rect -40700 5092 -40666 5122
rect -40700 5020 -40666 5054
rect -40700 4952 -40666 4982
rect -40700 4948 -40666 4952
rect -40700 4884 -40666 4910
rect -40700 4876 -40666 4884
rect -40700 4816 -40666 4838
rect -40700 4804 -40666 4816
rect -40700 4748 -40666 4766
rect -40700 4732 -40666 4748
rect -40700 4680 -40666 4694
rect -40700 4660 -40666 4680
rect 104 5382 138 5402
rect 104 5368 138 5382
rect 104 5314 138 5330
rect 104 5296 138 5314
rect 104 5246 138 5258
rect 104 5224 138 5246
rect 104 5178 138 5186
rect 104 5152 138 5178
rect 104 5110 138 5114
rect 104 5080 138 5110
rect 104 5008 138 5042
rect 104 4940 138 4970
rect 104 4936 138 4940
rect 104 4872 138 4898
rect 104 4864 138 4872
rect 104 4804 138 4826
rect 104 4792 138 4804
rect 104 4736 138 4754
rect 104 4720 138 4736
rect 104 4668 138 4682
rect 104 4648 138 4668
rect 200 5382 234 5402
rect 200 5368 234 5382
rect 200 5314 234 5330
rect 200 5296 234 5314
rect 200 5246 234 5258
rect 200 5224 234 5246
rect 200 5178 234 5186
rect 200 5152 234 5178
rect 200 5110 234 5114
rect 200 5080 234 5110
rect 200 5008 234 5042
rect 200 4940 234 4970
rect 200 4936 234 4940
rect 200 4872 234 4898
rect 200 4864 234 4872
rect 200 4804 234 4826
rect 200 4792 234 4804
rect 200 4736 234 4754
rect 200 4720 234 4736
rect 200 4668 234 4682
rect 200 4648 234 4668
rect 296 5382 330 5402
rect 296 5368 330 5382
rect 296 5314 330 5330
rect 296 5296 330 5314
rect 296 5246 330 5258
rect 296 5224 330 5246
rect 296 5178 330 5186
rect 296 5152 330 5178
rect 296 5110 330 5114
rect 296 5080 330 5110
rect 296 5008 330 5042
rect 296 4940 330 4970
rect 296 4936 330 4940
rect 296 4872 330 4898
rect 296 4864 330 4872
rect 296 4804 330 4826
rect 296 4792 330 4804
rect 296 4736 330 4754
rect 296 4720 330 4736
rect 296 4668 330 4682
rect 296 4648 330 4668
rect 392 5382 426 5402
rect 392 5368 426 5382
rect 392 5314 426 5330
rect 392 5296 426 5314
rect 392 5246 426 5258
rect 392 5224 426 5246
rect 392 5178 426 5186
rect 392 5152 426 5178
rect 392 5110 426 5114
rect 392 5080 426 5110
rect 392 5008 426 5042
rect 392 4940 426 4970
rect 392 4936 426 4940
rect 392 4872 426 4898
rect 392 4864 426 4872
rect 392 4804 426 4826
rect 392 4792 426 4804
rect 392 4736 426 4754
rect 392 4720 426 4736
rect 392 4668 426 4682
rect 392 4648 426 4668
rect 488 5382 522 5402
rect 488 5368 522 5382
rect 488 5314 522 5330
rect 488 5296 522 5314
rect 488 5246 522 5258
rect 488 5224 522 5246
rect 488 5178 522 5186
rect 488 5152 522 5178
rect 488 5110 522 5114
rect 488 5080 522 5110
rect 488 5008 522 5042
rect 488 4940 522 4970
rect 488 4936 522 4940
rect 488 4872 522 4898
rect 488 4864 522 4872
rect 488 4804 522 4826
rect 488 4792 522 4804
rect 488 4736 522 4754
rect 488 4720 522 4736
rect 488 4668 522 4682
rect 488 4648 522 4668
rect 584 5382 618 5402
rect 584 5368 618 5382
rect 584 5314 618 5330
rect 584 5296 618 5314
rect 584 5246 618 5258
rect 584 5224 618 5246
rect 584 5178 618 5186
rect 584 5152 618 5178
rect 584 5110 618 5114
rect 584 5080 618 5110
rect 584 5008 618 5042
rect 584 4940 618 4970
rect 584 4936 618 4940
rect 584 4872 618 4898
rect 584 4864 618 4872
rect 584 4804 618 4826
rect 584 4792 618 4804
rect 584 4736 618 4754
rect 584 4720 618 4736
rect 584 4668 618 4682
rect 584 4648 618 4668
rect 680 5382 714 5402
rect 680 5368 714 5382
rect 680 5314 714 5330
rect 680 5296 714 5314
rect 680 5246 714 5258
rect 680 5224 714 5246
rect 680 5178 714 5186
rect 680 5152 714 5178
rect 680 5110 714 5114
rect 680 5080 714 5110
rect 680 5008 714 5042
rect 680 4940 714 4970
rect 680 4936 714 4940
rect 680 4872 714 4898
rect 680 4864 714 4872
rect 680 4804 714 4826
rect 680 4792 714 4804
rect 680 4736 714 4754
rect 680 4720 714 4736
rect 680 4668 714 4682
rect 680 4648 714 4668
rect 776 5382 810 5402
rect 776 5368 810 5382
rect 776 5314 810 5330
rect 776 5296 810 5314
rect 776 5246 810 5258
rect 776 5224 810 5246
rect 776 5178 810 5186
rect 776 5152 810 5178
rect 776 5110 810 5114
rect 776 5080 810 5110
rect 776 5008 810 5042
rect 776 4940 810 4970
rect 776 4936 810 4940
rect 776 4872 810 4898
rect 776 4864 810 4872
rect 776 4804 810 4826
rect 776 4792 810 4804
rect 776 4736 810 4754
rect 776 4720 810 4736
rect 776 4668 810 4682
rect 776 4648 810 4668
rect 872 5382 906 5402
rect 872 5368 906 5382
rect 872 5314 906 5330
rect 872 5296 906 5314
rect 872 5246 906 5258
rect 872 5224 906 5246
rect 872 5178 906 5186
rect 872 5152 906 5178
rect 872 5110 906 5114
rect 872 5080 906 5110
rect 872 5008 906 5042
rect 872 4940 906 4970
rect 872 4936 906 4940
rect 872 4872 906 4898
rect 872 4864 906 4872
rect 872 4804 906 4826
rect 872 4792 906 4804
rect 872 4736 906 4754
rect 872 4720 906 4736
rect 872 4668 906 4682
rect 872 4648 906 4668
rect 968 5382 1002 5402
rect 968 5368 1002 5382
rect 968 5314 1002 5330
rect 968 5296 1002 5314
rect 968 5246 1002 5258
rect 968 5224 1002 5246
rect 968 5178 1002 5186
rect 968 5152 1002 5178
rect 968 5110 1002 5114
rect 968 5080 1002 5110
rect 968 5008 1002 5042
rect 968 4940 1002 4970
rect 968 4936 1002 4940
rect 968 4872 1002 4898
rect 968 4864 1002 4872
rect 968 4804 1002 4826
rect 968 4792 1002 4804
rect 968 4736 1002 4754
rect 968 4720 1002 4736
rect 968 4668 1002 4682
rect 968 4648 1002 4668
rect 1064 5382 1098 5402
rect 1064 5368 1098 5382
rect 1064 5314 1098 5330
rect 1064 5296 1098 5314
rect 1064 5246 1098 5258
rect 1064 5224 1098 5246
rect 1064 5178 1098 5186
rect 1064 5152 1098 5178
rect 1064 5110 1098 5114
rect 1064 5080 1098 5110
rect 1064 5008 1098 5042
rect 1064 4940 1098 4970
rect 1064 4936 1098 4940
rect 1064 4872 1098 4898
rect 1064 4864 1098 4872
rect 1064 4804 1098 4826
rect 1064 4792 1098 4804
rect 1064 4736 1098 4754
rect 1064 4720 1098 4736
rect 1064 4668 1098 4682
rect 1064 4648 1098 4668
rect 1160 5382 1194 5402
rect 1160 5368 1194 5382
rect 1160 5314 1194 5330
rect 1160 5296 1194 5314
rect 1160 5246 1194 5258
rect 1160 5224 1194 5246
rect 1160 5178 1194 5186
rect 1160 5152 1194 5178
rect 1160 5110 1194 5114
rect 1160 5080 1194 5110
rect 1160 5008 1194 5042
rect 1160 4940 1194 4970
rect 1160 4936 1194 4940
rect 1160 4872 1194 4898
rect 1160 4864 1194 4872
rect 1160 4804 1194 4826
rect 1160 4792 1194 4804
rect 1160 4736 1194 4754
rect 1160 4720 1194 4736
rect 1160 4668 1194 4682
rect 1160 4648 1194 4668
rect 1256 5382 1290 5402
rect 1256 5368 1290 5382
rect 1256 5314 1290 5330
rect 1256 5296 1290 5314
rect 1256 5246 1290 5258
rect 1256 5224 1290 5246
rect 1256 5178 1290 5186
rect 1256 5152 1290 5178
rect 1256 5110 1290 5114
rect 1256 5080 1290 5110
rect 1256 5008 1290 5042
rect 1256 4940 1290 4970
rect 1256 4936 1290 4940
rect 1256 4872 1290 4898
rect 1256 4864 1290 4872
rect 1256 4804 1290 4826
rect 1256 4792 1290 4804
rect 1256 4736 1290 4754
rect 1256 4720 1290 4736
rect 1256 4668 1290 4682
rect 1256 4648 1290 4668
rect 1352 5382 1386 5402
rect 1352 5368 1386 5382
rect 1352 5314 1386 5330
rect 1352 5296 1386 5314
rect 1352 5246 1386 5258
rect 1352 5224 1386 5246
rect 1352 5178 1386 5186
rect 1352 5152 1386 5178
rect 1352 5110 1386 5114
rect 1352 5080 1386 5110
rect 1352 5008 1386 5042
rect 1352 4940 1386 4970
rect 1352 4936 1386 4940
rect 1352 4872 1386 4898
rect 1352 4864 1386 4872
rect 1352 4804 1386 4826
rect 1352 4792 1386 4804
rect 1352 4736 1386 4754
rect 1352 4720 1386 4736
rect 1352 4668 1386 4682
rect 1352 4648 1386 4668
rect 1448 5382 1482 5402
rect 1448 5368 1482 5382
rect 1448 5314 1482 5330
rect 1448 5296 1482 5314
rect 1448 5246 1482 5258
rect 1448 5224 1482 5246
rect 1448 5178 1482 5186
rect 1448 5152 1482 5178
rect 1448 5110 1482 5114
rect 1448 5080 1482 5110
rect 1448 5008 1482 5042
rect 1448 4940 1482 4970
rect 1448 4936 1482 4940
rect 1448 4872 1482 4898
rect 1448 4864 1482 4872
rect 1448 4804 1482 4826
rect 1448 4792 1482 4804
rect 1448 4736 1482 4754
rect 1448 4720 1482 4736
rect 1448 4668 1482 4682
rect 1448 4648 1482 4668
rect 1544 5382 1578 5402
rect 1544 5368 1578 5382
rect 1544 5314 1578 5330
rect 1544 5296 1578 5314
rect 1544 5246 1578 5258
rect 1544 5224 1578 5246
rect 1544 5178 1578 5186
rect 1544 5152 1578 5178
rect 1544 5110 1578 5114
rect 1544 5080 1578 5110
rect 1544 5008 1578 5042
rect 1544 4940 1578 4970
rect 1544 4936 1578 4940
rect 1544 4872 1578 4898
rect 1544 4864 1578 4872
rect 1544 4804 1578 4826
rect 1544 4792 1578 4804
rect 1544 4736 1578 4754
rect 1544 4720 1578 4736
rect 1544 4668 1578 4682
rect 1544 4648 1578 4668
rect 1640 5382 1674 5402
rect 1640 5368 1674 5382
rect 1640 5314 1674 5330
rect 1640 5296 1674 5314
rect 1640 5246 1674 5258
rect 1640 5224 1674 5246
rect 1640 5178 1674 5186
rect 1640 5152 1674 5178
rect 1640 5110 1674 5114
rect 1640 5080 1674 5110
rect 1640 5008 1674 5042
rect 1640 4940 1674 4970
rect 1640 4936 1674 4940
rect 1640 4872 1674 4898
rect 1640 4864 1674 4872
rect 1640 4804 1674 4826
rect 1640 4792 1674 4804
rect 1640 4736 1674 4754
rect 1640 4720 1674 4736
rect 1640 4668 1674 4682
rect 1640 4648 1674 4668
rect 1736 5382 1770 5402
rect 1736 5368 1770 5382
rect 1736 5314 1770 5330
rect 1736 5296 1770 5314
rect 1736 5246 1770 5258
rect 1736 5224 1770 5246
rect 1736 5178 1770 5186
rect 1736 5152 1770 5178
rect 1736 5110 1770 5114
rect 1736 5080 1770 5110
rect 1736 5008 1770 5042
rect 1736 4940 1770 4970
rect 1736 4936 1770 4940
rect 1736 4872 1770 4898
rect 1736 4864 1770 4872
rect 1736 4804 1770 4826
rect 1736 4792 1770 4804
rect 1736 4736 1770 4754
rect 1736 4720 1770 4736
rect 1736 4668 1770 4682
rect 1736 4648 1770 4668
rect 1832 5382 1866 5402
rect 1832 5368 1866 5382
rect 1832 5314 1866 5330
rect 1832 5296 1866 5314
rect 1832 5246 1866 5258
rect 1832 5224 1866 5246
rect 1832 5178 1866 5186
rect 1832 5152 1866 5178
rect 1832 5110 1866 5114
rect 1832 5080 1866 5110
rect 1832 5008 1866 5042
rect 1832 4940 1866 4970
rect 1832 4936 1866 4940
rect 1832 4872 1866 4898
rect 1832 4864 1866 4872
rect 1832 4804 1866 4826
rect 1832 4792 1866 4804
rect 1832 4736 1866 4754
rect 1832 4720 1866 4736
rect 1832 4668 1866 4682
rect 1832 4648 1866 4668
rect 1928 5382 1962 5402
rect 1928 5368 1962 5382
rect 1928 5314 1962 5330
rect 1928 5296 1962 5314
rect 1928 5246 1962 5258
rect 1928 5224 1962 5246
rect 1928 5178 1962 5186
rect 1928 5152 1962 5178
rect 1928 5110 1962 5114
rect 1928 5080 1962 5110
rect 1928 5008 1962 5042
rect 1928 4940 1962 4970
rect 1928 4936 1962 4940
rect 1928 4872 1962 4898
rect 1928 4864 1962 4872
rect 1928 4804 1962 4826
rect 1928 4792 1962 4804
rect 1928 4736 1962 4754
rect 1928 4720 1962 4736
rect 1928 4668 1962 4682
rect 1928 4648 1962 4668
rect -42525 -4780 -42491 -4760
rect -42525 -4794 -42491 -4780
rect -42525 -4848 -42491 -4832
rect -42525 -4866 -42491 -4848
rect -42525 -4916 -42491 -4904
rect -42525 -4938 -42491 -4916
rect -42525 -4984 -42491 -4976
rect -42525 -5010 -42491 -4984
rect -42525 -5052 -42491 -5048
rect -42525 -5082 -42491 -5052
rect -42525 -5154 -42491 -5120
rect -42525 -5222 -42491 -5192
rect -42525 -5226 -42491 -5222
rect -42525 -5290 -42491 -5264
rect -42525 -5298 -42491 -5290
rect -42525 -5358 -42491 -5336
rect -42525 -5370 -42491 -5358
rect -42525 -5426 -42491 -5408
rect -42525 -5442 -42491 -5426
rect -42525 -5494 -42491 -5480
rect -42525 -5514 -42491 -5494
rect -42429 -4780 -42395 -4760
rect -42429 -4794 -42395 -4780
rect -42429 -4848 -42395 -4832
rect -42429 -4866 -42395 -4848
rect -42429 -4916 -42395 -4904
rect -42429 -4938 -42395 -4916
rect -42429 -4984 -42395 -4976
rect -42429 -5010 -42395 -4984
rect -42429 -5052 -42395 -5048
rect -42429 -5082 -42395 -5052
rect -42429 -5154 -42395 -5120
rect -42429 -5222 -42395 -5192
rect -42429 -5226 -42395 -5222
rect -42429 -5290 -42395 -5264
rect -42429 -5298 -42395 -5290
rect -42429 -5358 -42395 -5336
rect -42429 -5370 -42395 -5358
rect -42429 -5426 -42395 -5408
rect -42429 -5442 -42395 -5426
rect -42429 -5494 -42395 -5480
rect -42429 -5514 -42395 -5494
rect -42333 -4780 -42299 -4760
rect -42333 -4794 -42299 -4780
rect -42333 -4848 -42299 -4832
rect -42333 -4866 -42299 -4848
rect -42333 -4916 -42299 -4904
rect -42333 -4938 -42299 -4916
rect -42333 -4984 -42299 -4976
rect -42333 -5010 -42299 -4984
rect -42333 -5052 -42299 -5048
rect -42333 -5082 -42299 -5052
rect -42333 -5154 -42299 -5120
rect -42333 -5222 -42299 -5192
rect -42333 -5226 -42299 -5222
rect -42333 -5290 -42299 -5264
rect -42333 -5298 -42299 -5290
rect -42333 -5358 -42299 -5336
rect -42333 -5370 -42299 -5358
rect -42333 -5426 -42299 -5408
rect -42333 -5442 -42299 -5426
rect -42333 -5494 -42299 -5480
rect -42333 -5514 -42299 -5494
rect -42237 -4780 -42203 -4760
rect -42237 -4794 -42203 -4780
rect -42237 -4848 -42203 -4832
rect -42237 -4866 -42203 -4848
rect -42237 -4916 -42203 -4904
rect -42237 -4938 -42203 -4916
rect -42237 -4984 -42203 -4976
rect -42237 -5010 -42203 -4984
rect -42237 -5052 -42203 -5048
rect -42237 -5082 -42203 -5052
rect -42237 -5154 -42203 -5120
rect -42237 -5222 -42203 -5192
rect -42237 -5226 -42203 -5222
rect -42237 -5290 -42203 -5264
rect -42237 -5298 -42203 -5290
rect -42237 -5358 -42203 -5336
rect -42237 -5370 -42203 -5358
rect -42237 -5426 -42203 -5408
rect -42237 -5442 -42203 -5426
rect -42237 -5494 -42203 -5480
rect -42237 -5514 -42203 -5494
rect -42141 -4780 -42107 -4760
rect -42141 -4794 -42107 -4780
rect -42141 -4848 -42107 -4832
rect -42141 -4866 -42107 -4848
rect -42141 -4916 -42107 -4904
rect -42141 -4938 -42107 -4916
rect -42141 -4984 -42107 -4976
rect -42141 -5010 -42107 -4984
rect -42141 -5052 -42107 -5048
rect -42141 -5082 -42107 -5052
rect -42141 -5154 -42107 -5120
rect -42141 -5222 -42107 -5192
rect -42141 -5226 -42107 -5222
rect -42141 -5290 -42107 -5264
rect -42141 -5298 -42107 -5290
rect -42141 -5358 -42107 -5336
rect -42141 -5370 -42107 -5358
rect -42141 -5426 -42107 -5408
rect -42141 -5442 -42107 -5426
rect -42141 -5494 -42107 -5480
rect -42141 -5514 -42107 -5494
rect -42045 -4780 -42011 -4760
rect -42045 -4794 -42011 -4780
rect -42045 -4848 -42011 -4832
rect -42045 -4866 -42011 -4848
rect -42045 -4916 -42011 -4904
rect -42045 -4938 -42011 -4916
rect -42045 -4984 -42011 -4976
rect -42045 -5010 -42011 -4984
rect -42045 -5052 -42011 -5048
rect -42045 -5082 -42011 -5052
rect -42045 -5154 -42011 -5120
rect -42045 -5222 -42011 -5192
rect -42045 -5226 -42011 -5222
rect -42045 -5290 -42011 -5264
rect -42045 -5298 -42011 -5290
rect -42045 -5358 -42011 -5336
rect -42045 -5370 -42011 -5358
rect -42045 -5426 -42011 -5408
rect -42045 -5442 -42011 -5426
rect -42045 -5494 -42011 -5480
rect -42045 -5514 -42011 -5494
rect -41949 -4780 -41915 -4760
rect -41949 -4794 -41915 -4780
rect -41949 -4848 -41915 -4832
rect -41949 -4866 -41915 -4848
rect -41949 -4916 -41915 -4904
rect -41949 -4938 -41915 -4916
rect -41949 -4984 -41915 -4976
rect -41949 -5010 -41915 -4984
rect -41949 -5052 -41915 -5048
rect -41949 -5082 -41915 -5052
rect -41949 -5154 -41915 -5120
rect -41949 -5222 -41915 -5192
rect -41949 -5226 -41915 -5222
rect -41949 -5290 -41915 -5264
rect -41949 -5298 -41915 -5290
rect -41949 -5358 -41915 -5336
rect -41949 -5370 -41915 -5358
rect -41949 -5426 -41915 -5408
rect -41949 -5442 -41915 -5426
rect -41949 -5494 -41915 -5480
rect -41949 -5514 -41915 -5494
rect -41853 -4780 -41819 -4760
rect -41853 -4794 -41819 -4780
rect -41853 -4848 -41819 -4832
rect -41853 -4866 -41819 -4848
rect -41853 -4916 -41819 -4904
rect -41853 -4938 -41819 -4916
rect -41853 -4984 -41819 -4976
rect -41853 -5010 -41819 -4984
rect -41853 -5052 -41819 -5048
rect -41853 -5082 -41819 -5052
rect -41853 -5154 -41819 -5120
rect -41853 -5222 -41819 -5192
rect -41853 -5226 -41819 -5222
rect -41853 -5290 -41819 -5264
rect -41853 -5298 -41819 -5290
rect -41853 -5358 -41819 -5336
rect -41853 -5370 -41819 -5358
rect -41853 -5426 -41819 -5408
rect -41853 -5442 -41819 -5426
rect -41853 -5494 -41819 -5480
rect -41853 -5514 -41819 -5494
rect -41757 -4780 -41723 -4760
rect -41757 -4794 -41723 -4780
rect -41757 -4848 -41723 -4832
rect -41757 -4866 -41723 -4848
rect -41757 -4916 -41723 -4904
rect -41757 -4938 -41723 -4916
rect -41757 -4984 -41723 -4976
rect -41757 -5010 -41723 -4984
rect -41757 -5052 -41723 -5048
rect -41757 -5082 -41723 -5052
rect -41757 -5154 -41723 -5120
rect -41757 -5222 -41723 -5192
rect -41757 -5226 -41723 -5222
rect -41757 -5290 -41723 -5264
rect -41757 -5298 -41723 -5290
rect -41757 -5358 -41723 -5336
rect -41757 -5370 -41723 -5358
rect -41757 -5426 -41723 -5408
rect -41757 -5442 -41723 -5426
rect -41757 -5494 -41723 -5480
rect -41757 -5514 -41723 -5494
rect -41661 -4780 -41627 -4760
rect -41661 -4794 -41627 -4780
rect -41661 -4848 -41627 -4832
rect -41661 -4866 -41627 -4848
rect -41661 -4916 -41627 -4904
rect -41661 -4938 -41627 -4916
rect -41661 -4984 -41627 -4976
rect -41661 -5010 -41627 -4984
rect -41661 -5052 -41627 -5048
rect -41661 -5082 -41627 -5052
rect -41661 -5154 -41627 -5120
rect -41661 -5222 -41627 -5192
rect -41661 -5226 -41627 -5222
rect -41661 -5290 -41627 -5264
rect -41661 -5298 -41627 -5290
rect -41661 -5358 -41627 -5336
rect -41661 -5370 -41627 -5358
rect -41661 -5426 -41627 -5408
rect -41661 -5442 -41627 -5426
rect -41661 -5494 -41627 -5480
rect -41661 -5514 -41627 -5494
rect -41565 -4780 -41531 -4760
rect -41565 -4794 -41531 -4780
rect -41565 -4848 -41531 -4832
rect -41565 -4866 -41531 -4848
rect -41565 -4916 -41531 -4904
rect -41565 -4938 -41531 -4916
rect -41565 -4984 -41531 -4976
rect -41565 -5010 -41531 -4984
rect -41565 -5052 -41531 -5048
rect -41565 -5082 -41531 -5052
rect -41565 -5154 -41531 -5120
rect -41565 -5222 -41531 -5192
rect -41565 -5226 -41531 -5222
rect -41565 -5290 -41531 -5264
rect -41565 -5298 -41531 -5290
rect -41565 -5358 -41531 -5336
rect -41565 -5370 -41531 -5358
rect -41565 -5426 -41531 -5408
rect -41565 -5442 -41531 -5426
rect -41565 -5494 -41531 -5480
rect -41565 -5514 -41531 -5494
rect -41469 -4780 -41435 -4760
rect -41469 -4794 -41435 -4780
rect -41469 -4848 -41435 -4832
rect -41469 -4866 -41435 -4848
rect -41469 -4916 -41435 -4904
rect -41469 -4938 -41435 -4916
rect -41469 -4984 -41435 -4976
rect -41469 -5010 -41435 -4984
rect -41469 -5052 -41435 -5048
rect -41469 -5082 -41435 -5052
rect -41469 -5154 -41435 -5120
rect -41469 -5222 -41435 -5192
rect -41469 -5226 -41435 -5222
rect -41469 -5290 -41435 -5264
rect -41469 -5298 -41435 -5290
rect -41469 -5358 -41435 -5336
rect -41469 -5370 -41435 -5358
rect -41469 -5426 -41435 -5408
rect -41469 -5442 -41435 -5426
rect -41469 -5494 -41435 -5480
rect -41469 -5514 -41435 -5494
rect -41373 -4780 -41339 -4760
rect -41373 -4794 -41339 -4780
rect -41373 -4848 -41339 -4832
rect -41373 -4866 -41339 -4848
rect -41373 -4916 -41339 -4904
rect -41373 -4938 -41339 -4916
rect -41373 -4984 -41339 -4976
rect -41373 -5010 -41339 -4984
rect -41373 -5052 -41339 -5048
rect -41373 -5082 -41339 -5052
rect -41373 -5154 -41339 -5120
rect -41373 -5222 -41339 -5192
rect -41373 -5226 -41339 -5222
rect -41373 -5290 -41339 -5264
rect -41373 -5298 -41339 -5290
rect -41373 -5358 -41339 -5336
rect -41373 -5370 -41339 -5358
rect -41373 -5426 -41339 -5408
rect -41373 -5442 -41339 -5426
rect -41373 -5494 -41339 -5480
rect -41373 -5514 -41339 -5494
rect -41277 -4780 -41243 -4760
rect -41277 -4794 -41243 -4780
rect -41277 -4848 -41243 -4832
rect -41277 -4866 -41243 -4848
rect -41277 -4916 -41243 -4904
rect -41277 -4938 -41243 -4916
rect -41277 -4984 -41243 -4976
rect -41277 -5010 -41243 -4984
rect -41277 -5052 -41243 -5048
rect -41277 -5082 -41243 -5052
rect -41277 -5154 -41243 -5120
rect -41277 -5222 -41243 -5192
rect -41277 -5226 -41243 -5222
rect -41277 -5290 -41243 -5264
rect -41277 -5298 -41243 -5290
rect -41277 -5358 -41243 -5336
rect -41277 -5370 -41243 -5358
rect -41277 -5426 -41243 -5408
rect -41277 -5442 -41243 -5426
rect -41277 -5494 -41243 -5480
rect -41277 -5514 -41243 -5494
rect -41181 -4780 -41147 -4760
rect -41181 -4794 -41147 -4780
rect -41181 -4848 -41147 -4832
rect -41181 -4866 -41147 -4848
rect -41181 -4916 -41147 -4904
rect -41181 -4938 -41147 -4916
rect -41181 -4984 -41147 -4976
rect -41181 -5010 -41147 -4984
rect -41181 -5052 -41147 -5048
rect -41181 -5082 -41147 -5052
rect -41181 -5154 -41147 -5120
rect -41181 -5222 -41147 -5192
rect -41181 -5226 -41147 -5222
rect -41181 -5290 -41147 -5264
rect -41181 -5298 -41147 -5290
rect -41181 -5358 -41147 -5336
rect -41181 -5370 -41147 -5358
rect -41181 -5426 -41147 -5408
rect -41181 -5442 -41147 -5426
rect -41181 -5494 -41147 -5480
rect -41181 -5514 -41147 -5494
rect -41085 -4780 -41051 -4760
rect -41085 -4794 -41051 -4780
rect -41085 -4848 -41051 -4832
rect -41085 -4866 -41051 -4848
rect -41085 -4916 -41051 -4904
rect -41085 -4938 -41051 -4916
rect -41085 -4984 -41051 -4976
rect -41085 -5010 -41051 -4984
rect -41085 -5052 -41051 -5048
rect -41085 -5082 -41051 -5052
rect -41085 -5154 -41051 -5120
rect -41085 -5222 -41051 -5192
rect -41085 -5226 -41051 -5222
rect -41085 -5290 -41051 -5264
rect -41085 -5298 -41051 -5290
rect -41085 -5358 -41051 -5336
rect -41085 -5370 -41051 -5358
rect -41085 -5426 -41051 -5408
rect -41085 -5442 -41051 -5426
rect -41085 -5494 -41051 -5480
rect -41085 -5514 -41051 -5494
rect -40989 -4780 -40955 -4760
rect -40989 -4794 -40955 -4780
rect -40989 -4848 -40955 -4832
rect -40989 -4866 -40955 -4848
rect -40989 -4916 -40955 -4904
rect -40989 -4938 -40955 -4916
rect -40989 -4984 -40955 -4976
rect -40989 -5010 -40955 -4984
rect -40989 -5052 -40955 -5048
rect -40989 -5082 -40955 -5052
rect -40989 -5154 -40955 -5120
rect -40989 -5222 -40955 -5192
rect -40989 -5226 -40955 -5222
rect -40989 -5290 -40955 -5264
rect -40989 -5298 -40955 -5290
rect -40989 -5358 -40955 -5336
rect -40989 -5370 -40955 -5358
rect -40989 -5426 -40955 -5408
rect -40989 -5442 -40955 -5426
rect -40989 -5494 -40955 -5480
rect -40989 -5514 -40955 -5494
rect -40893 -4780 -40859 -4760
rect -40893 -4794 -40859 -4780
rect -40893 -4848 -40859 -4832
rect -40893 -4866 -40859 -4848
rect -40893 -4916 -40859 -4904
rect -40893 -4938 -40859 -4916
rect -40893 -4984 -40859 -4976
rect -40893 -5010 -40859 -4984
rect -40893 -5052 -40859 -5048
rect -40893 -5082 -40859 -5052
rect -40893 -5154 -40859 -5120
rect -40893 -5222 -40859 -5192
rect -40893 -5226 -40859 -5222
rect -40893 -5290 -40859 -5264
rect -40893 -5298 -40859 -5290
rect -40893 -5358 -40859 -5336
rect -40893 -5370 -40859 -5358
rect -40893 -5426 -40859 -5408
rect -40893 -5442 -40859 -5426
rect -40893 -5494 -40859 -5480
rect -40893 -5514 -40859 -5494
rect -40797 -4780 -40763 -4760
rect -40797 -4794 -40763 -4780
rect -40797 -4848 -40763 -4832
rect -40797 -4866 -40763 -4848
rect -40797 -4916 -40763 -4904
rect -40797 -4938 -40763 -4916
rect -40797 -4984 -40763 -4976
rect -40797 -5010 -40763 -4984
rect -40797 -5052 -40763 -5048
rect -40797 -5082 -40763 -5052
rect -40797 -5154 -40763 -5120
rect -40797 -5222 -40763 -5192
rect -40797 -5226 -40763 -5222
rect -40797 -5290 -40763 -5264
rect -40797 -5298 -40763 -5290
rect -40797 -5358 -40763 -5336
rect -40797 -5370 -40763 -5358
rect -40797 -5426 -40763 -5408
rect -40797 -5442 -40763 -5426
rect -40797 -5494 -40763 -5480
rect -40797 -5514 -40763 -5494
rect -40701 -4780 -40667 -4760
rect -40701 -4794 -40667 -4780
rect -40701 -4848 -40667 -4832
rect -40701 -4866 -40667 -4848
rect -40701 -4916 -40667 -4904
rect -40701 -4938 -40667 -4916
rect -40701 -4984 -40667 -4976
rect -40701 -5010 -40667 -4984
rect -40701 -5052 -40667 -5048
rect -40701 -5082 -40667 -5052
rect -40701 -5154 -40667 -5120
rect -40701 -5222 -40667 -5192
rect -40701 -5226 -40667 -5222
rect -40701 -5290 -40667 -5264
rect -40701 -5298 -40667 -5290
rect -40701 -5358 -40667 -5336
rect -40701 -5370 -40667 -5358
rect -40701 -5426 -40667 -5408
rect -40701 -5442 -40667 -5426
rect -40701 -5494 -40667 -5480
rect -40701 -5514 -40667 -5494
rect 116 -4806 150 -4786
rect 116 -4820 150 -4806
rect 116 -4874 150 -4858
rect 116 -4892 150 -4874
rect 116 -4942 150 -4930
rect 116 -4964 150 -4942
rect 116 -5010 150 -5002
rect 116 -5036 150 -5010
rect 116 -5078 150 -5074
rect 116 -5108 150 -5078
rect 116 -5180 150 -5146
rect 116 -5248 150 -5218
rect 116 -5252 150 -5248
rect 116 -5316 150 -5290
rect 116 -5324 150 -5316
rect 116 -5384 150 -5362
rect 116 -5396 150 -5384
rect 116 -5452 150 -5434
rect 116 -5468 150 -5452
rect 116 -5520 150 -5506
rect 116 -5540 150 -5520
rect 212 -4806 246 -4786
rect 212 -4820 246 -4806
rect 212 -4874 246 -4858
rect 212 -4892 246 -4874
rect 212 -4942 246 -4930
rect 212 -4964 246 -4942
rect 212 -5010 246 -5002
rect 212 -5036 246 -5010
rect 212 -5078 246 -5074
rect 212 -5108 246 -5078
rect 212 -5180 246 -5146
rect 212 -5248 246 -5218
rect 212 -5252 246 -5248
rect 212 -5316 246 -5290
rect 212 -5324 246 -5316
rect 212 -5384 246 -5362
rect 212 -5396 246 -5384
rect 212 -5452 246 -5434
rect 212 -5468 246 -5452
rect 212 -5520 246 -5506
rect 212 -5540 246 -5520
rect 308 -4806 342 -4786
rect 308 -4820 342 -4806
rect 308 -4874 342 -4858
rect 308 -4892 342 -4874
rect 308 -4942 342 -4930
rect 308 -4964 342 -4942
rect 308 -5010 342 -5002
rect 308 -5036 342 -5010
rect 308 -5078 342 -5074
rect 308 -5108 342 -5078
rect 308 -5180 342 -5146
rect 308 -5248 342 -5218
rect 308 -5252 342 -5248
rect 308 -5316 342 -5290
rect 308 -5324 342 -5316
rect 308 -5384 342 -5362
rect 308 -5396 342 -5384
rect 308 -5452 342 -5434
rect 308 -5468 342 -5452
rect 308 -5520 342 -5506
rect 308 -5540 342 -5520
rect 404 -4806 438 -4786
rect 404 -4820 438 -4806
rect 404 -4874 438 -4858
rect 404 -4892 438 -4874
rect 404 -4942 438 -4930
rect 404 -4964 438 -4942
rect 404 -5010 438 -5002
rect 404 -5036 438 -5010
rect 404 -5078 438 -5074
rect 404 -5108 438 -5078
rect 404 -5180 438 -5146
rect 404 -5248 438 -5218
rect 404 -5252 438 -5248
rect 404 -5316 438 -5290
rect 404 -5324 438 -5316
rect 404 -5384 438 -5362
rect 404 -5396 438 -5384
rect 404 -5452 438 -5434
rect 404 -5468 438 -5452
rect 404 -5520 438 -5506
rect 404 -5540 438 -5520
rect 500 -4806 534 -4786
rect 500 -4820 534 -4806
rect 500 -4874 534 -4858
rect 500 -4892 534 -4874
rect 500 -4942 534 -4930
rect 500 -4964 534 -4942
rect 500 -5010 534 -5002
rect 500 -5036 534 -5010
rect 500 -5078 534 -5074
rect 500 -5108 534 -5078
rect 500 -5180 534 -5146
rect 500 -5248 534 -5218
rect 500 -5252 534 -5248
rect 500 -5316 534 -5290
rect 500 -5324 534 -5316
rect 500 -5384 534 -5362
rect 500 -5396 534 -5384
rect 500 -5452 534 -5434
rect 500 -5468 534 -5452
rect 500 -5520 534 -5506
rect 500 -5540 534 -5520
rect 596 -4806 630 -4786
rect 596 -4820 630 -4806
rect 596 -4874 630 -4858
rect 596 -4892 630 -4874
rect 596 -4942 630 -4930
rect 596 -4964 630 -4942
rect 596 -5010 630 -5002
rect 596 -5036 630 -5010
rect 596 -5078 630 -5074
rect 596 -5108 630 -5078
rect 596 -5180 630 -5146
rect 596 -5248 630 -5218
rect 596 -5252 630 -5248
rect 596 -5316 630 -5290
rect 596 -5324 630 -5316
rect 596 -5384 630 -5362
rect 596 -5396 630 -5384
rect 596 -5452 630 -5434
rect 596 -5468 630 -5452
rect 596 -5520 630 -5506
rect 596 -5540 630 -5520
rect 692 -4806 726 -4786
rect 692 -4820 726 -4806
rect 692 -4874 726 -4858
rect 692 -4892 726 -4874
rect 692 -4942 726 -4930
rect 692 -4964 726 -4942
rect 692 -5010 726 -5002
rect 692 -5036 726 -5010
rect 692 -5078 726 -5074
rect 692 -5108 726 -5078
rect 692 -5180 726 -5146
rect 692 -5248 726 -5218
rect 692 -5252 726 -5248
rect 692 -5316 726 -5290
rect 692 -5324 726 -5316
rect 692 -5384 726 -5362
rect 692 -5396 726 -5384
rect 692 -5452 726 -5434
rect 692 -5468 726 -5452
rect 692 -5520 726 -5506
rect 692 -5540 726 -5520
rect 788 -4806 822 -4786
rect 788 -4820 822 -4806
rect 788 -4874 822 -4858
rect 788 -4892 822 -4874
rect 788 -4942 822 -4930
rect 788 -4964 822 -4942
rect 788 -5010 822 -5002
rect 788 -5036 822 -5010
rect 788 -5078 822 -5074
rect 788 -5108 822 -5078
rect 788 -5180 822 -5146
rect 788 -5248 822 -5218
rect 788 -5252 822 -5248
rect 788 -5316 822 -5290
rect 788 -5324 822 -5316
rect 788 -5384 822 -5362
rect 788 -5396 822 -5384
rect 788 -5452 822 -5434
rect 788 -5468 822 -5452
rect 788 -5520 822 -5506
rect 788 -5540 822 -5520
rect 884 -4806 918 -4786
rect 884 -4820 918 -4806
rect 884 -4874 918 -4858
rect 884 -4892 918 -4874
rect 884 -4942 918 -4930
rect 884 -4964 918 -4942
rect 884 -5010 918 -5002
rect 884 -5036 918 -5010
rect 884 -5078 918 -5074
rect 884 -5108 918 -5078
rect 884 -5180 918 -5146
rect 884 -5248 918 -5218
rect 884 -5252 918 -5248
rect 884 -5316 918 -5290
rect 884 -5324 918 -5316
rect 884 -5384 918 -5362
rect 884 -5396 918 -5384
rect 884 -5452 918 -5434
rect 884 -5468 918 -5452
rect 884 -5520 918 -5506
rect 884 -5540 918 -5520
rect 980 -4806 1014 -4786
rect 980 -4820 1014 -4806
rect 980 -4874 1014 -4858
rect 980 -4892 1014 -4874
rect 980 -4942 1014 -4930
rect 980 -4964 1014 -4942
rect 980 -5010 1014 -5002
rect 980 -5036 1014 -5010
rect 980 -5078 1014 -5074
rect 980 -5108 1014 -5078
rect 980 -5180 1014 -5146
rect 980 -5248 1014 -5218
rect 980 -5252 1014 -5248
rect 980 -5316 1014 -5290
rect 980 -5324 1014 -5316
rect 980 -5384 1014 -5362
rect 980 -5396 1014 -5384
rect 980 -5452 1014 -5434
rect 980 -5468 1014 -5452
rect 980 -5520 1014 -5506
rect 980 -5540 1014 -5520
rect 1076 -4806 1110 -4786
rect 1076 -4820 1110 -4806
rect 1076 -4874 1110 -4858
rect 1076 -4892 1110 -4874
rect 1076 -4942 1110 -4930
rect 1076 -4964 1110 -4942
rect 1076 -5010 1110 -5002
rect 1076 -5036 1110 -5010
rect 1076 -5078 1110 -5074
rect 1076 -5108 1110 -5078
rect 1076 -5180 1110 -5146
rect 1076 -5248 1110 -5218
rect 1076 -5252 1110 -5248
rect 1076 -5316 1110 -5290
rect 1076 -5324 1110 -5316
rect 1076 -5384 1110 -5362
rect 1076 -5396 1110 -5384
rect 1076 -5452 1110 -5434
rect 1076 -5468 1110 -5452
rect 1076 -5520 1110 -5506
rect 1076 -5540 1110 -5520
rect 1172 -4806 1206 -4786
rect 1172 -4820 1206 -4806
rect 1172 -4874 1206 -4858
rect 1172 -4892 1206 -4874
rect 1172 -4942 1206 -4930
rect 1172 -4964 1206 -4942
rect 1172 -5010 1206 -5002
rect 1172 -5036 1206 -5010
rect 1172 -5078 1206 -5074
rect 1172 -5108 1206 -5078
rect 1172 -5180 1206 -5146
rect 1172 -5248 1206 -5218
rect 1172 -5252 1206 -5248
rect 1172 -5316 1206 -5290
rect 1172 -5324 1206 -5316
rect 1172 -5384 1206 -5362
rect 1172 -5396 1206 -5384
rect 1172 -5452 1206 -5434
rect 1172 -5468 1206 -5452
rect 1172 -5520 1206 -5506
rect 1172 -5540 1206 -5520
rect 1268 -4806 1302 -4786
rect 1268 -4820 1302 -4806
rect 1268 -4874 1302 -4858
rect 1268 -4892 1302 -4874
rect 1268 -4942 1302 -4930
rect 1268 -4964 1302 -4942
rect 1268 -5010 1302 -5002
rect 1268 -5036 1302 -5010
rect 1268 -5078 1302 -5074
rect 1268 -5108 1302 -5078
rect 1268 -5180 1302 -5146
rect 1268 -5248 1302 -5218
rect 1268 -5252 1302 -5248
rect 1268 -5316 1302 -5290
rect 1268 -5324 1302 -5316
rect 1268 -5384 1302 -5362
rect 1268 -5396 1302 -5384
rect 1268 -5452 1302 -5434
rect 1268 -5468 1302 -5452
rect 1268 -5520 1302 -5506
rect 1268 -5540 1302 -5520
rect 1364 -4806 1398 -4786
rect 1364 -4820 1398 -4806
rect 1364 -4874 1398 -4858
rect 1364 -4892 1398 -4874
rect 1364 -4942 1398 -4930
rect 1364 -4964 1398 -4942
rect 1364 -5010 1398 -5002
rect 1364 -5036 1398 -5010
rect 1364 -5078 1398 -5074
rect 1364 -5108 1398 -5078
rect 1364 -5180 1398 -5146
rect 1364 -5248 1398 -5218
rect 1364 -5252 1398 -5248
rect 1364 -5316 1398 -5290
rect 1364 -5324 1398 -5316
rect 1364 -5384 1398 -5362
rect 1364 -5396 1398 -5384
rect 1364 -5452 1398 -5434
rect 1364 -5468 1398 -5452
rect 1364 -5520 1398 -5506
rect 1364 -5540 1398 -5520
rect 1460 -4806 1494 -4786
rect 1460 -4820 1494 -4806
rect 1460 -4874 1494 -4858
rect 1460 -4892 1494 -4874
rect 1460 -4942 1494 -4930
rect 1460 -4964 1494 -4942
rect 1460 -5010 1494 -5002
rect 1460 -5036 1494 -5010
rect 1460 -5078 1494 -5074
rect 1460 -5108 1494 -5078
rect 1460 -5180 1494 -5146
rect 1460 -5248 1494 -5218
rect 1460 -5252 1494 -5248
rect 1460 -5316 1494 -5290
rect 1460 -5324 1494 -5316
rect 1460 -5384 1494 -5362
rect 1460 -5396 1494 -5384
rect 1460 -5452 1494 -5434
rect 1460 -5468 1494 -5452
rect 1460 -5520 1494 -5506
rect 1460 -5540 1494 -5520
rect 1556 -4806 1590 -4786
rect 1556 -4820 1590 -4806
rect 1556 -4874 1590 -4858
rect 1556 -4892 1590 -4874
rect 1556 -4942 1590 -4930
rect 1556 -4964 1590 -4942
rect 1556 -5010 1590 -5002
rect 1556 -5036 1590 -5010
rect 1556 -5078 1590 -5074
rect 1556 -5108 1590 -5078
rect 1556 -5180 1590 -5146
rect 1556 -5248 1590 -5218
rect 1556 -5252 1590 -5248
rect 1556 -5316 1590 -5290
rect 1556 -5324 1590 -5316
rect 1556 -5384 1590 -5362
rect 1556 -5396 1590 -5384
rect 1556 -5452 1590 -5434
rect 1556 -5468 1590 -5452
rect 1556 -5520 1590 -5506
rect 1556 -5540 1590 -5520
rect 1652 -4806 1686 -4786
rect 1652 -4820 1686 -4806
rect 1652 -4874 1686 -4858
rect 1652 -4892 1686 -4874
rect 1652 -4942 1686 -4930
rect 1652 -4964 1686 -4942
rect 1652 -5010 1686 -5002
rect 1652 -5036 1686 -5010
rect 1652 -5078 1686 -5074
rect 1652 -5108 1686 -5078
rect 1652 -5180 1686 -5146
rect 1652 -5248 1686 -5218
rect 1652 -5252 1686 -5248
rect 1652 -5316 1686 -5290
rect 1652 -5324 1686 -5316
rect 1652 -5384 1686 -5362
rect 1652 -5396 1686 -5384
rect 1652 -5452 1686 -5434
rect 1652 -5468 1686 -5452
rect 1652 -5520 1686 -5506
rect 1652 -5540 1686 -5520
rect 1748 -4806 1782 -4786
rect 1748 -4820 1782 -4806
rect 1748 -4874 1782 -4858
rect 1748 -4892 1782 -4874
rect 1748 -4942 1782 -4930
rect 1748 -4964 1782 -4942
rect 1748 -5010 1782 -5002
rect 1748 -5036 1782 -5010
rect 1748 -5078 1782 -5074
rect 1748 -5108 1782 -5078
rect 1748 -5180 1782 -5146
rect 1748 -5248 1782 -5218
rect 1748 -5252 1782 -5248
rect 1748 -5316 1782 -5290
rect 1748 -5324 1782 -5316
rect 1748 -5384 1782 -5362
rect 1748 -5396 1782 -5384
rect 1748 -5452 1782 -5434
rect 1748 -5468 1782 -5452
rect 1748 -5520 1782 -5506
rect 1748 -5540 1782 -5520
rect 1844 -4806 1878 -4786
rect 1844 -4820 1878 -4806
rect 1844 -4874 1878 -4858
rect 1844 -4892 1878 -4874
rect 1844 -4942 1878 -4930
rect 1844 -4964 1878 -4942
rect 1844 -5010 1878 -5002
rect 1844 -5036 1878 -5010
rect 1844 -5078 1878 -5074
rect 1844 -5108 1878 -5078
rect 1844 -5180 1878 -5146
rect 1844 -5248 1878 -5218
rect 1844 -5252 1878 -5248
rect 1844 -5316 1878 -5290
rect 1844 -5324 1878 -5316
rect 1844 -5384 1878 -5362
rect 1844 -5396 1878 -5384
rect 1844 -5452 1878 -5434
rect 1844 -5468 1878 -5452
rect 1844 -5520 1878 -5506
rect 1844 -5540 1878 -5520
rect 1940 -4806 1974 -4786
rect 1940 -4820 1974 -4806
rect 1940 -4874 1974 -4858
rect 1940 -4892 1974 -4874
rect 1940 -4942 1974 -4930
rect 1940 -4964 1974 -4942
rect 1940 -5010 1974 -5002
rect 1940 -5036 1974 -5010
rect 1940 -5078 1974 -5074
rect 1940 -5108 1974 -5078
rect 1940 -5180 1974 -5146
rect 1940 -5248 1974 -5218
rect 1940 -5252 1974 -5248
rect 1940 -5316 1974 -5290
rect 1940 -5324 1974 -5316
rect 1940 -5384 1974 -5362
rect 1940 -5396 1974 -5384
rect 1940 -5452 1974 -5434
rect 1940 -5468 1974 -5452
rect 1940 -5520 1974 -5506
rect 1940 -5540 1974 -5520
<< metal1 >>
rect -74485 38544 -74165 38550
rect -74485 38236 -74479 38544
rect -74171 38236 -74165 38544
rect -74485 38210 -74165 38236
rect -73485 38544 -73165 38550
rect -73485 38236 -73479 38544
rect -73171 38236 -73165 38544
rect -73485 38210 -73165 38236
rect -72485 38544 -72165 38550
rect -72485 38236 -72479 38544
rect -72171 38236 -72165 38544
rect -72485 38210 -72165 38236
rect -71485 38544 -71165 38550
rect -71485 38236 -71479 38544
rect -71171 38236 -71165 38544
rect -71485 38210 -71165 38236
rect -70485 38544 -70165 38550
rect -70485 38236 -70479 38544
rect -70171 38236 -70165 38544
rect -70485 38210 -70165 38236
rect -69485 38544 -69165 38550
rect -69485 38236 -69479 38544
rect -69171 38236 -69165 38544
rect -69485 38210 -69165 38236
rect -68485 38544 -68165 38550
rect -68485 38236 -68479 38544
rect -68171 38236 -68165 38544
rect -68485 38210 -68165 38236
rect -67485 38544 -67165 38550
rect -67485 38236 -67479 38544
rect -67171 38236 -67165 38544
rect -67485 38210 -67165 38236
rect -66485 38544 -66165 38550
rect -66485 38236 -66479 38544
rect -66171 38236 -66165 38544
rect -66485 38210 -66165 38236
rect -65485 38544 -65165 38550
rect -65485 38236 -65479 38544
rect -65171 38236 -65165 38544
rect -65485 38210 -65165 38236
rect -64485 38544 -64165 38550
rect -64485 38236 -64479 38544
rect -64171 38236 -64165 38544
rect -64485 38210 -64165 38236
rect -63485 38544 -63165 38550
rect -63485 38236 -63479 38544
rect -63171 38236 -63165 38544
rect -63485 38210 -63165 38236
rect -62485 38544 -62165 38550
rect -62485 38236 -62479 38544
rect -62171 38236 -62165 38544
rect -62485 38210 -62165 38236
rect -61485 38544 -61165 38550
rect -61485 38236 -61479 38544
rect -61171 38236 -61165 38544
rect -61485 38210 -61165 38236
rect -60485 38544 -60165 38550
rect -60485 38236 -60479 38544
rect -60171 38236 -60165 38544
rect -60485 38210 -60165 38236
rect -59485 38544 -59165 38550
rect -59485 38236 -59479 38544
rect -59171 38236 -59165 38544
rect -59485 38210 -59165 38236
rect 9994 38544 10314 38550
rect 9994 38236 10000 38544
rect 10308 38236 10314 38544
rect 9994 38210 10314 38236
rect 10994 38544 11314 38550
rect 10994 38236 11000 38544
rect 11308 38236 11314 38544
rect 10994 38210 11314 38236
rect 11994 38544 12314 38550
rect 11994 38236 12000 38544
rect 12308 38236 12314 38544
rect 11994 38210 12314 38236
rect 12994 38544 13314 38550
rect 12994 38236 13000 38544
rect 13308 38236 13314 38544
rect 12994 38210 13314 38236
rect 13994 38544 14314 38550
rect 13994 38236 14000 38544
rect 14308 38236 14314 38544
rect 13994 38210 14314 38236
rect 14994 38544 15314 38550
rect 14994 38236 15000 38544
rect 15308 38236 15314 38544
rect 14994 38210 15314 38236
rect 15994 38544 16314 38550
rect 15994 38236 16000 38544
rect 16308 38236 16314 38544
rect 15994 38210 16314 38236
rect 16994 38544 17314 38550
rect 16994 38236 17000 38544
rect 17308 38236 17314 38544
rect 16994 38210 17314 38236
rect 17994 38544 18314 38550
rect 17994 38236 18000 38544
rect 18308 38236 18314 38544
rect 17994 38210 18314 38236
rect 18994 38544 19314 38550
rect 18994 38236 19000 38544
rect 19308 38236 19314 38544
rect 18994 38210 19314 38236
rect 19994 38544 20314 38550
rect 19994 38236 20000 38544
rect 20308 38236 20314 38544
rect 19994 38210 20314 38236
rect 20994 38544 21314 38550
rect 20994 38236 21000 38544
rect 21308 38236 21314 38544
rect 20994 38210 21314 38236
rect 21994 38544 22314 38550
rect 21994 38236 22000 38544
rect 22308 38236 22314 38544
rect 21994 38210 22314 38236
rect 22994 38544 23314 38550
rect 22994 38236 23000 38544
rect 23308 38236 23314 38544
rect 22994 38210 23314 38236
rect 23994 38544 24314 38550
rect 23994 38236 24000 38544
rect 24308 38236 24314 38544
rect 23994 38210 24314 38236
rect 24994 38544 25314 38550
rect 24994 38236 25000 38544
rect 25308 38236 25314 38544
rect 24994 38210 25314 38236
rect 25994 38544 26314 38550
rect 25994 38236 26000 38544
rect 26308 38236 26314 38544
rect 25994 38210 26314 38236
rect 26994 38544 27314 38550
rect 26994 38236 27000 38544
rect 27308 38236 27314 38544
rect 26994 38210 27314 38236
rect 27994 38544 28314 38550
rect 27994 38236 28000 38544
rect 28308 38236 28314 38544
rect 27994 38210 28314 38236
rect 28994 38544 29314 38550
rect 28994 38236 29000 38544
rect 29308 38236 29314 38544
rect 28994 38210 29314 38236
rect 29994 38544 30314 38550
rect 29994 38236 30000 38544
rect 30308 38236 30314 38544
rect 29994 38210 30314 38236
rect 30994 38544 31314 38550
rect 30994 38236 31000 38544
rect 31308 38236 31314 38544
rect 30994 38210 31314 38236
rect 31994 38544 32314 38550
rect 31994 38236 32000 38544
rect 32308 38236 32314 38544
rect 31994 38210 32314 38236
rect 32994 38544 33314 38550
rect 32994 38236 33000 38544
rect 33308 38236 33314 38544
rect 32994 38210 33314 38236
rect 33994 38544 34314 38550
rect 33994 38236 34000 38544
rect 34308 38236 34314 38544
rect 33994 38210 34314 38236
rect -74825 38204 -58825 38210
rect -74825 37896 -74819 38204
rect -74511 38172 -74139 38204
rect -74511 37928 -74447 38172
rect -74203 37928 -74139 38172
rect -74511 37896 -74139 37928
rect -73511 38172 -73139 38204
rect -73511 37928 -73447 38172
rect -73203 37928 -73139 38172
rect -73511 37896 -73139 37928
rect -72511 38172 -72139 38204
rect -72511 37928 -72447 38172
rect -72203 37928 -72139 38172
rect -72511 37896 -72139 37928
rect -71511 38172 -71139 38204
rect -71511 37928 -71447 38172
rect -71203 37928 -71139 38172
rect -71511 37896 -71139 37928
rect -70511 38172 -70139 38204
rect -70511 37928 -70447 38172
rect -70203 37928 -70139 38172
rect -70511 37896 -70139 37928
rect -69511 38172 -69139 38204
rect -69511 37928 -69447 38172
rect -69203 37928 -69139 38172
rect -69511 37896 -69139 37928
rect -68511 38172 -68139 38204
rect -68511 37928 -68447 38172
rect -68203 37928 -68139 38172
rect -68511 37896 -68139 37928
rect -67511 38172 -67139 38204
rect -67511 37928 -67447 38172
rect -67203 37928 -67139 38172
rect -67511 37896 -67139 37928
rect -66511 38172 -66139 38204
rect -66511 37928 -66447 38172
rect -66203 37928 -66139 38172
rect -66511 37896 -66139 37928
rect -65511 38172 -65139 38204
rect -65511 37928 -65447 38172
rect -65203 37928 -65139 38172
rect -65511 37896 -65139 37928
rect -64511 38172 -64139 38204
rect -64511 37928 -64447 38172
rect -64203 37928 -64139 38172
rect -64511 37896 -64139 37928
rect -63511 38172 -63139 38204
rect -63511 37928 -63447 38172
rect -63203 37928 -63139 38172
rect -63511 37896 -63139 37928
rect -62511 38172 -62139 38204
rect -62511 37928 -62447 38172
rect -62203 37928 -62139 38172
rect -62511 37896 -62139 37928
rect -61511 38172 -61139 38204
rect -61511 37928 -61447 38172
rect -61203 37928 -61139 38172
rect -61511 37896 -61139 37928
rect -60511 38172 -60139 38204
rect -60511 37928 -60447 38172
rect -60203 37928 -60139 38172
rect -60511 37896 -60139 37928
rect -59511 38172 -59139 38204
rect -59511 37928 -59447 38172
rect -59203 37928 -59139 38172
rect -59511 37896 -59139 37928
rect -58831 37896 -58825 38204
rect -74825 37890 -58825 37896
rect 9654 38204 34654 38210
rect 9654 37896 9660 38204
rect 9968 38172 10340 38204
rect 9968 37928 10032 38172
rect 10276 37928 10340 38172
rect 9968 37896 10340 37928
rect 10968 38172 11340 38204
rect 10968 37928 11032 38172
rect 11276 37928 11340 38172
rect 10968 37896 11340 37928
rect 11968 38172 12340 38204
rect 11968 37928 12032 38172
rect 12276 37928 12340 38172
rect 11968 37896 12340 37928
rect 12968 38172 13340 38204
rect 12968 37928 13032 38172
rect 13276 37928 13340 38172
rect 12968 37896 13340 37928
rect 13968 38172 14340 38204
rect 13968 37928 14032 38172
rect 14276 37928 14340 38172
rect 13968 37896 14340 37928
rect 14968 38172 15340 38204
rect 14968 37928 15032 38172
rect 15276 37928 15340 38172
rect 14968 37896 15340 37928
rect 15968 38172 16340 38204
rect 15968 37928 16032 38172
rect 16276 37928 16340 38172
rect 15968 37896 16340 37928
rect 16968 38172 17340 38204
rect 16968 37928 17032 38172
rect 17276 37928 17340 38172
rect 16968 37896 17340 37928
rect 17968 38172 18340 38204
rect 17968 37928 18032 38172
rect 18276 37928 18340 38172
rect 17968 37896 18340 37928
rect 18968 38172 19340 38204
rect 18968 37928 19032 38172
rect 19276 37928 19340 38172
rect 18968 37896 19340 37928
rect 19968 38172 20340 38204
rect 19968 37928 20032 38172
rect 20276 37928 20340 38172
rect 19968 37896 20340 37928
rect 20968 38172 21340 38204
rect 20968 37928 21032 38172
rect 21276 37928 21340 38172
rect 20968 37896 21340 37928
rect 21968 38172 22340 38204
rect 21968 37928 22032 38172
rect 22276 37928 22340 38172
rect 21968 37896 22340 37928
rect 22968 38172 23340 38204
rect 22968 37928 23032 38172
rect 23276 37928 23340 38172
rect 22968 37896 23340 37928
rect 23968 38172 24340 38204
rect 23968 37928 24032 38172
rect 24276 37928 24340 38172
rect 23968 37896 24340 37928
rect 24968 38172 25340 38204
rect 24968 37928 25032 38172
rect 25276 37928 25340 38172
rect 24968 37896 25340 37928
rect 25968 38172 26340 38204
rect 25968 37928 26032 38172
rect 26276 37928 26340 38172
rect 25968 37896 26340 37928
rect 26968 38172 27340 38204
rect 26968 37928 27032 38172
rect 27276 37928 27340 38172
rect 26968 37896 27340 37928
rect 27968 38172 28340 38204
rect 27968 37928 28032 38172
rect 28276 37928 28340 38172
rect 27968 37896 28340 37928
rect 28968 38172 29340 38204
rect 28968 37928 29032 38172
rect 29276 37928 29340 38172
rect 28968 37896 29340 37928
rect 29968 38172 30340 38204
rect 29968 37928 30032 38172
rect 30276 37928 30340 38172
rect 29968 37896 30340 37928
rect 30968 38172 31340 38204
rect 30968 37928 31032 38172
rect 31276 37928 31340 38172
rect 30968 37896 31340 37928
rect 31968 38172 32340 38204
rect 31968 37928 32032 38172
rect 32276 37928 32340 38172
rect 31968 37896 32340 37928
rect 32968 38172 33340 38204
rect 32968 37928 33032 38172
rect 33276 37928 33340 38172
rect 32968 37896 33340 37928
rect 33968 38172 34340 38204
rect 33968 37928 34032 38172
rect 34276 37928 34340 38172
rect 33968 37896 34340 37928
rect 34648 37896 34654 38204
rect 9654 37890 34654 37896
rect -74485 37864 -74165 37890
rect -74485 37236 -74479 37864
rect -74171 37236 -74165 37864
rect -74485 37210 -74165 37236
rect -73485 37864 -73165 37890
rect -73485 37236 -73479 37864
rect -73171 37236 -73165 37864
rect -73485 37210 -73165 37236
rect -72485 37864 -72165 37890
rect -72485 37236 -72479 37864
rect -72171 37236 -72165 37864
rect -72485 37210 -72165 37236
rect -71485 37864 -71165 37890
rect -71485 37236 -71479 37864
rect -71171 37236 -71165 37864
rect -71485 37210 -71165 37236
rect -70485 37864 -70165 37890
rect -70485 37236 -70479 37864
rect -70171 37236 -70165 37864
rect -70485 37210 -70165 37236
rect -69485 37864 -69165 37890
rect -69485 37236 -69479 37864
rect -69171 37236 -69165 37864
rect -69485 37210 -69165 37236
rect -68485 37864 -68165 37890
rect -68485 37236 -68479 37864
rect -68171 37236 -68165 37864
rect -68485 37210 -68165 37236
rect -67485 37864 -67165 37890
rect -67485 37236 -67479 37864
rect -67171 37236 -67165 37864
rect -67485 37210 -67165 37236
rect -66485 37864 -66165 37890
rect -66485 37236 -66479 37864
rect -66171 37236 -66165 37864
rect -66485 37210 -66165 37236
rect -65485 37864 -65165 37890
rect -65485 37236 -65479 37864
rect -65171 37236 -65165 37864
rect -65485 37210 -65165 37236
rect -64485 37864 -64165 37890
rect -64485 37236 -64479 37864
rect -64171 37236 -64165 37864
rect -64485 37210 -64165 37236
rect -63485 37864 -63165 37890
rect -63485 37236 -63479 37864
rect -63171 37236 -63165 37864
rect -63485 37210 -63165 37236
rect -62485 37864 -62165 37890
rect -62485 37236 -62479 37864
rect -62171 37236 -62165 37864
rect -62485 37210 -62165 37236
rect -61485 37864 -61165 37890
rect -61485 37236 -61479 37864
rect -61171 37236 -61165 37864
rect -61485 37210 -61165 37236
rect -60485 37864 -60165 37890
rect -60485 37236 -60479 37864
rect -60171 37236 -60165 37864
rect -60485 37210 -60165 37236
rect -59485 37864 -59165 37890
rect -59485 37236 -59479 37864
rect -59171 37236 -59165 37864
rect -59485 37210 -59165 37236
rect 9994 37864 10314 37890
rect 9994 37236 10000 37864
rect 10308 37236 10314 37864
rect 9994 37210 10314 37236
rect 10994 37864 11314 37890
rect 10994 37236 11000 37864
rect 11308 37236 11314 37864
rect 10994 37210 11314 37236
rect 11994 37864 12314 37890
rect 11994 37236 12000 37864
rect 12308 37236 12314 37864
rect 11994 37210 12314 37236
rect 12994 37864 13314 37890
rect 12994 37236 13000 37864
rect 13308 37236 13314 37864
rect 12994 37210 13314 37236
rect 13994 37864 14314 37890
rect 13994 37236 14000 37864
rect 14308 37236 14314 37864
rect 13994 37210 14314 37236
rect 14994 37864 15314 37890
rect 14994 37236 15000 37864
rect 15308 37236 15314 37864
rect 14994 37210 15314 37236
rect 15994 37864 16314 37890
rect 15994 37236 16000 37864
rect 16308 37236 16314 37864
rect 15994 37210 16314 37236
rect 16994 37864 17314 37890
rect 16994 37236 17000 37864
rect 17308 37236 17314 37864
rect 16994 37210 17314 37236
rect 17994 37864 18314 37890
rect 17994 37236 18000 37864
rect 18308 37236 18314 37864
rect 17994 37210 18314 37236
rect 18994 37864 19314 37890
rect 18994 37236 19000 37864
rect 19308 37236 19314 37864
rect 18994 37210 19314 37236
rect 19994 37864 20314 37890
rect 19994 37236 20000 37864
rect 20308 37236 20314 37864
rect 19994 37210 20314 37236
rect 20994 37864 21314 37890
rect 20994 37236 21000 37864
rect 21308 37236 21314 37864
rect 20994 37210 21314 37236
rect 21994 37864 22314 37890
rect 21994 37236 22000 37864
rect 22308 37236 22314 37864
rect 21994 37210 22314 37236
rect 22994 37864 23314 37890
rect 22994 37236 23000 37864
rect 23308 37236 23314 37864
rect 22994 37210 23314 37236
rect 23994 37864 24314 37890
rect 23994 37236 24000 37864
rect 24308 37236 24314 37864
rect 23994 37210 24314 37236
rect 24994 37864 25314 37890
rect 24994 37236 25000 37864
rect 25308 37236 25314 37864
rect 24994 37210 25314 37236
rect 25994 37864 26314 37890
rect 25994 37236 26000 37864
rect 26308 37236 26314 37864
rect 25994 37210 26314 37236
rect 26994 37864 27314 37890
rect 26994 37236 27000 37864
rect 27308 37236 27314 37864
rect 26994 37210 27314 37236
rect 27994 37864 28314 37890
rect 27994 37236 28000 37864
rect 28308 37236 28314 37864
rect 27994 37210 28314 37236
rect 28994 37864 29314 37890
rect 28994 37236 29000 37864
rect 29308 37236 29314 37864
rect 28994 37210 29314 37236
rect 29994 37864 30314 37890
rect 29994 37236 30000 37864
rect 30308 37236 30314 37864
rect 29994 37210 30314 37236
rect 30994 37864 31314 37890
rect 30994 37236 31000 37864
rect 31308 37236 31314 37864
rect 30994 37210 31314 37236
rect 31994 37864 32314 37890
rect 31994 37236 32000 37864
rect 32308 37236 32314 37864
rect 31994 37210 32314 37236
rect 32994 37864 33314 37890
rect 32994 37236 33000 37864
rect 33308 37236 33314 37864
rect 32994 37210 33314 37236
rect 33994 37864 34314 37890
rect 33994 37236 34000 37864
rect 34308 37236 34314 37864
rect 33994 37210 34314 37236
rect -74825 37204 -58825 37210
rect -74825 36896 -74819 37204
rect -74511 37172 -74139 37204
rect -74511 36928 -74447 37172
rect -74203 36928 -74139 37172
rect -74511 36896 -74139 36928
rect -73511 37172 -73139 37204
rect -73511 36928 -73447 37172
rect -73203 36928 -73139 37172
rect -73511 36896 -73139 36928
rect -72511 37172 -72139 37204
rect -72511 36928 -72447 37172
rect -72203 36928 -72139 37172
rect -72511 36896 -72139 36928
rect -71511 37172 -71139 37204
rect -71511 36928 -71447 37172
rect -71203 36928 -71139 37172
rect -71511 36896 -71139 36928
rect -70511 37172 -70139 37204
rect -70511 36928 -70447 37172
rect -70203 36928 -70139 37172
rect -70511 36896 -70139 36928
rect -69511 37172 -69139 37204
rect -69511 36928 -69447 37172
rect -69203 36928 -69139 37172
rect -69511 36896 -69139 36928
rect -68511 37172 -68139 37204
rect -68511 36928 -68447 37172
rect -68203 36928 -68139 37172
rect -68511 36896 -68139 36928
rect -67511 37172 -67139 37204
rect -67511 36928 -67447 37172
rect -67203 36928 -67139 37172
rect -67511 36896 -67139 36928
rect -66511 37172 -66139 37204
rect -66511 36928 -66447 37172
rect -66203 36928 -66139 37172
rect -66511 36896 -66139 36928
rect -65511 37172 -65139 37204
rect -65511 36928 -65447 37172
rect -65203 36928 -65139 37172
rect -65511 36896 -65139 36928
rect -64511 37172 -64139 37204
rect -64511 36928 -64447 37172
rect -64203 36928 -64139 37172
rect -64511 36896 -64139 36928
rect -63511 37172 -63139 37204
rect -63511 36928 -63447 37172
rect -63203 36928 -63139 37172
rect -63511 36896 -63139 36928
rect -62511 37172 -62139 37204
rect -62511 36928 -62447 37172
rect -62203 36928 -62139 37172
rect -62511 36896 -62139 36928
rect -61511 37172 -61139 37204
rect -61511 36928 -61447 37172
rect -61203 36928 -61139 37172
rect -61511 36896 -61139 36928
rect -60511 37172 -60139 37204
rect -60511 36928 -60447 37172
rect -60203 36928 -60139 37172
rect -60511 36896 -60139 36928
rect -59511 37172 -59139 37204
rect -59511 36928 -59447 37172
rect -59203 36928 -59139 37172
rect -59511 36896 -59139 36928
rect -58831 36896 -58825 37204
rect -74825 36890 -58825 36896
rect 9654 37204 34654 37210
rect 9654 36896 9660 37204
rect 9968 37172 10340 37204
rect 9968 36928 10032 37172
rect 10276 36928 10340 37172
rect 9968 36896 10340 36928
rect 10968 37172 11340 37204
rect 10968 36928 11032 37172
rect 11276 36928 11340 37172
rect 10968 36896 11340 36928
rect 11968 37172 12340 37204
rect 11968 36928 12032 37172
rect 12276 36928 12340 37172
rect 11968 36896 12340 36928
rect 12968 37172 13340 37204
rect 12968 36928 13032 37172
rect 13276 36928 13340 37172
rect 12968 36896 13340 36928
rect 13968 37172 14340 37204
rect 13968 36928 14032 37172
rect 14276 36928 14340 37172
rect 13968 36896 14340 36928
rect 14968 37172 15340 37204
rect 14968 36928 15032 37172
rect 15276 36928 15340 37172
rect 14968 36896 15340 36928
rect 15968 37172 16340 37204
rect 15968 36928 16032 37172
rect 16276 36928 16340 37172
rect 15968 36896 16340 36928
rect 16968 37172 17340 37204
rect 16968 36928 17032 37172
rect 17276 36928 17340 37172
rect 16968 36896 17340 36928
rect 17968 37172 18340 37204
rect 17968 36928 18032 37172
rect 18276 36928 18340 37172
rect 17968 36896 18340 36928
rect 18968 37172 19340 37204
rect 18968 36928 19032 37172
rect 19276 36928 19340 37172
rect 18968 36896 19340 36928
rect 19968 37172 20340 37204
rect 19968 36928 20032 37172
rect 20276 36928 20340 37172
rect 19968 36896 20340 36928
rect 20968 37172 21340 37204
rect 20968 36928 21032 37172
rect 21276 36928 21340 37172
rect 20968 36896 21340 36928
rect 21968 37172 22340 37204
rect 21968 36928 22032 37172
rect 22276 36928 22340 37172
rect 21968 36896 22340 36928
rect 22968 37172 23340 37204
rect 22968 36928 23032 37172
rect 23276 36928 23340 37172
rect 22968 36896 23340 36928
rect 23968 37172 24340 37204
rect 23968 36928 24032 37172
rect 24276 36928 24340 37172
rect 23968 36896 24340 36928
rect 24968 37172 25340 37204
rect 24968 36928 25032 37172
rect 25276 36928 25340 37172
rect 24968 36896 25340 36928
rect 25968 37172 26340 37204
rect 25968 36928 26032 37172
rect 26276 36928 26340 37172
rect 25968 36896 26340 36928
rect 26968 37172 27340 37204
rect 26968 36928 27032 37172
rect 27276 36928 27340 37172
rect 26968 36896 27340 36928
rect 27968 37172 28340 37204
rect 27968 36928 28032 37172
rect 28276 36928 28340 37172
rect 27968 36896 28340 36928
rect 28968 37172 29340 37204
rect 28968 36928 29032 37172
rect 29276 36928 29340 37172
rect 28968 36896 29340 36928
rect 29968 37172 30340 37204
rect 29968 36928 30032 37172
rect 30276 36928 30340 37172
rect 29968 36896 30340 36928
rect 30968 37172 31340 37204
rect 30968 36928 31032 37172
rect 31276 36928 31340 37172
rect 30968 36896 31340 36928
rect 31968 37172 32340 37204
rect 31968 36928 32032 37172
rect 32276 36928 32340 37172
rect 31968 36896 32340 36928
rect 32968 37172 33340 37204
rect 32968 36928 33032 37172
rect 33276 36928 33340 37172
rect 32968 36896 33340 36928
rect 33968 37172 34340 37204
rect 33968 36928 34032 37172
rect 34276 36928 34340 37172
rect 33968 36896 34340 36928
rect 34648 36896 34654 37204
rect 9654 36890 34654 36896
rect -74485 36864 -74165 36890
rect -74485 36236 -74479 36864
rect -74171 36236 -74165 36864
rect -74485 36210 -74165 36236
rect -73485 36864 -73165 36890
rect -73485 36236 -73479 36864
rect -73171 36236 -73165 36864
rect -73485 36210 -73165 36236
rect -72485 36864 -72165 36890
rect -72485 36236 -72479 36864
rect -72171 36236 -72165 36864
rect -72485 36210 -72165 36236
rect -71485 36864 -71165 36890
rect -71485 36236 -71479 36864
rect -71171 36236 -71165 36864
rect -71485 36210 -71165 36236
rect -70485 36864 -70165 36890
rect -70485 36236 -70479 36864
rect -70171 36236 -70165 36864
rect -70485 36210 -70165 36236
rect -69485 36864 -69165 36890
rect -69485 36236 -69479 36864
rect -69171 36236 -69165 36864
rect -69485 36210 -69165 36236
rect -68485 36864 -68165 36890
rect -68485 36236 -68479 36864
rect -68171 36236 -68165 36864
rect -68485 36210 -68165 36236
rect -67485 36864 -67165 36890
rect -67485 36236 -67479 36864
rect -67171 36236 -67165 36864
rect -67485 36210 -67165 36236
rect -66485 36864 -66165 36890
rect -66485 36236 -66479 36864
rect -66171 36236 -66165 36864
rect -66485 36210 -66165 36236
rect -65485 36864 -65165 36890
rect -65485 36236 -65479 36864
rect -65171 36236 -65165 36864
rect -65485 36210 -65165 36236
rect -64485 36864 -64165 36890
rect -64485 36236 -64479 36864
rect -64171 36236 -64165 36864
rect -64485 36210 -64165 36236
rect -63485 36864 -63165 36890
rect -63485 36236 -63479 36864
rect -63171 36236 -63165 36864
rect -63485 36210 -63165 36236
rect -62485 36864 -62165 36890
rect -62485 36236 -62479 36864
rect -62171 36236 -62165 36864
rect -62485 36210 -62165 36236
rect -61485 36864 -61165 36890
rect -61485 36236 -61479 36864
rect -61171 36236 -61165 36864
rect -61485 36210 -61165 36236
rect -60485 36864 -60165 36890
rect -60485 36236 -60479 36864
rect -60171 36236 -60165 36864
rect -60485 36210 -60165 36236
rect -59485 36864 -59165 36890
rect -59485 36236 -59479 36864
rect -59171 36236 -59165 36864
rect -59485 36210 -59165 36236
rect 9994 36864 10314 36890
rect 9994 36236 10000 36864
rect 10308 36236 10314 36864
rect 9994 36210 10314 36236
rect 10994 36864 11314 36890
rect 10994 36236 11000 36864
rect 11308 36236 11314 36864
rect 10994 36210 11314 36236
rect 11994 36864 12314 36890
rect 11994 36236 12000 36864
rect 12308 36236 12314 36864
rect 11994 36210 12314 36236
rect 12994 36864 13314 36890
rect 12994 36236 13000 36864
rect 13308 36236 13314 36864
rect 12994 36210 13314 36236
rect 13994 36864 14314 36890
rect 13994 36236 14000 36864
rect 14308 36236 14314 36864
rect 13994 36210 14314 36236
rect 14994 36864 15314 36890
rect 14994 36236 15000 36864
rect 15308 36236 15314 36864
rect 14994 36210 15314 36236
rect 15994 36864 16314 36890
rect 15994 36236 16000 36864
rect 16308 36236 16314 36864
rect 15994 36210 16314 36236
rect 16994 36864 17314 36890
rect 16994 36236 17000 36864
rect 17308 36236 17314 36864
rect 16994 36210 17314 36236
rect 17994 36864 18314 36890
rect 17994 36236 18000 36864
rect 18308 36236 18314 36864
rect 17994 36210 18314 36236
rect 18994 36864 19314 36890
rect 18994 36236 19000 36864
rect 19308 36236 19314 36864
rect 18994 36210 19314 36236
rect 19994 36864 20314 36890
rect 19994 36236 20000 36864
rect 20308 36236 20314 36864
rect 19994 36210 20314 36236
rect 20994 36864 21314 36890
rect 20994 36236 21000 36864
rect 21308 36236 21314 36864
rect 20994 36210 21314 36236
rect 21994 36864 22314 36890
rect 21994 36236 22000 36864
rect 22308 36236 22314 36864
rect 21994 36210 22314 36236
rect 22994 36864 23314 36890
rect 22994 36236 23000 36864
rect 23308 36236 23314 36864
rect 22994 36210 23314 36236
rect 23994 36864 24314 36890
rect 23994 36236 24000 36864
rect 24308 36236 24314 36864
rect 23994 36210 24314 36236
rect 24994 36864 25314 36890
rect 24994 36236 25000 36864
rect 25308 36236 25314 36864
rect 24994 36210 25314 36236
rect 25994 36864 26314 36890
rect 25994 36236 26000 36864
rect 26308 36236 26314 36864
rect 25994 36210 26314 36236
rect 26994 36864 27314 36890
rect 26994 36236 27000 36864
rect 27308 36236 27314 36864
rect 26994 36210 27314 36236
rect 27994 36864 28314 36890
rect 27994 36236 28000 36864
rect 28308 36236 28314 36864
rect 27994 36210 28314 36236
rect 28994 36864 29314 36890
rect 28994 36236 29000 36864
rect 29308 36236 29314 36864
rect 28994 36210 29314 36236
rect 29994 36864 30314 36890
rect 29994 36236 30000 36864
rect 30308 36236 30314 36864
rect 29994 36210 30314 36236
rect 30994 36864 31314 36890
rect 30994 36236 31000 36864
rect 31308 36236 31314 36864
rect 30994 36210 31314 36236
rect 31994 36864 32314 36890
rect 31994 36236 32000 36864
rect 32308 36236 32314 36864
rect 31994 36210 32314 36236
rect 32994 36864 33314 36890
rect 32994 36236 33000 36864
rect 33308 36236 33314 36864
rect 32994 36210 33314 36236
rect 33994 36864 34314 36890
rect 33994 36236 34000 36864
rect 34308 36236 34314 36864
rect 33994 36210 34314 36236
rect -74825 36204 -58825 36210
rect -74825 35896 -74819 36204
rect -74511 36172 -74139 36204
rect -74511 35928 -74447 36172
rect -74203 35928 -74139 36172
rect -74511 35896 -74139 35928
rect -73511 36172 -73139 36204
rect -73511 35928 -73447 36172
rect -73203 35928 -73139 36172
rect -73511 35896 -73139 35928
rect -72511 36172 -72139 36204
rect -72511 35928 -72447 36172
rect -72203 35928 -72139 36172
rect -72511 35896 -72139 35928
rect -71511 36172 -71139 36204
rect -71511 35928 -71447 36172
rect -71203 35928 -71139 36172
rect -71511 35896 -71139 35928
rect -70511 36172 -70139 36204
rect -70511 35928 -70447 36172
rect -70203 35928 -70139 36172
rect -70511 35896 -70139 35928
rect -69511 36172 -69139 36204
rect -69511 35928 -69447 36172
rect -69203 35928 -69139 36172
rect -69511 35896 -69139 35928
rect -68511 36172 -68139 36204
rect -68511 35928 -68447 36172
rect -68203 35928 -68139 36172
rect -68511 35896 -68139 35928
rect -67511 36172 -67139 36204
rect -67511 35928 -67447 36172
rect -67203 35928 -67139 36172
rect -67511 35896 -67139 35928
rect -66511 36172 -66139 36204
rect -66511 35928 -66447 36172
rect -66203 35928 -66139 36172
rect -66511 35896 -66139 35928
rect -65511 36172 -65139 36204
rect -65511 35928 -65447 36172
rect -65203 35928 -65139 36172
rect -65511 35896 -65139 35928
rect -64511 36172 -64139 36204
rect -64511 35928 -64447 36172
rect -64203 35928 -64139 36172
rect -64511 35896 -64139 35928
rect -63511 36172 -63139 36204
rect -63511 35928 -63447 36172
rect -63203 35928 -63139 36172
rect -63511 35896 -63139 35928
rect -62511 36172 -62139 36204
rect -62511 35928 -62447 36172
rect -62203 35928 -62139 36172
rect -62511 35896 -62139 35928
rect -61511 36172 -61139 36204
rect -61511 35928 -61447 36172
rect -61203 35928 -61139 36172
rect -61511 35896 -61139 35928
rect -60511 36172 -60139 36204
rect -60511 35928 -60447 36172
rect -60203 35928 -60139 36172
rect -60511 35896 -60139 35928
rect -59511 36172 -59139 36204
rect -59511 35928 -59447 36172
rect -59203 35928 -59139 36172
rect -59511 35896 -59139 35928
rect -58831 35896 -58825 36204
rect -74825 35890 -58825 35896
rect 9654 36204 34654 36210
rect 9654 35896 9660 36204
rect 9968 36172 10340 36204
rect 9968 35928 10032 36172
rect 10276 35928 10340 36172
rect 9968 35896 10340 35928
rect 10968 36172 11340 36204
rect 10968 35928 11032 36172
rect 11276 35928 11340 36172
rect 10968 35896 11340 35928
rect 11968 36172 12340 36204
rect 11968 35928 12032 36172
rect 12276 35928 12340 36172
rect 11968 35896 12340 35928
rect 12968 36172 13340 36204
rect 12968 35928 13032 36172
rect 13276 35928 13340 36172
rect 12968 35896 13340 35928
rect 13968 36172 14340 36204
rect 13968 35928 14032 36172
rect 14276 35928 14340 36172
rect 13968 35896 14340 35928
rect 14968 36172 15340 36204
rect 14968 35928 15032 36172
rect 15276 35928 15340 36172
rect 14968 35896 15340 35928
rect 15968 36172 16340 36204
rect 15968 35928 16032 36172
rect 16276 35928 16340 36172
rect 15968 35896 16340 35928
rect 16968 36172 17340 36204
rect 16968 35928 17032 36172
rect 17276 35928 17340 36172
rect 16968 35896 17340 35928
rect 17968 36172 18340 36204
rect 17968 35928 18032 36172
rect 18276 35928 18340 36172
rect 17968 35896 18340 35928
rect 18968 36172 19340 36204
rect 18968 35928 19032 36172
rect 19276 35928 19340 36172
rect 18968 35896 19340 35928
rect 19968 36172 20340 36204
rect 19968 35928 20032 36172
rect 20276 35928 20340 36172
rect 19968 35896 20340 35928
rect 20968 36172 21340 36204
rect 20968 35928 21032 36172
rect 21276 35928 21340 36172
rect 20968 35896 21340 35928
rect 21968 36172 22340 36204
rect 21968 35928 22032 36172
rect 22276 35928 22340 36172
rect 21968 35896 22340 35928
rect 22968 36172 23340 36204
rect 22968 35928 23032 36172
rect 23276 35928 23340 36172
rect 22968 35896 23340 35928
rect 23968 36172 24340 36204
rect 23968 35928 24032 36172
rect 24276 35928 24340 36172
rect 23968 35896 24340 35928
rect 24968 36172 25340 36204
rect 24968 35928 25032 36172
rect 25276 35928 25340 36172
rect 24968 35896 25340 35928
rect 25968 36172 26340 36204
rect 25968 35928 26032 36172
rect 26276 35928 26340 36172
rect 25968 35896 26340 35928
rect 26968 36172 27340 36204
rect 26968 35928 27032 36172
rect 27276 35928 27340 36172
rect 26968 35896 27340 35928
rect 27968 36172 28340 36204
rect 27968 35928 28032 36172
rect 28276 35928 28340 36172
rect 27968 35896 28340 35928
rect 28968 36172 29340 36204
rect 28968 35928 29032 36172
rect 29276 35928 29340 36172
rect 28968 35896 29340 35928
rect 29968 36172 30340 36204
rect 29968 35928 30032 36172
rect 30276 35928 30340 36172
rect 29968 35896 30340 35928
rect 30968 36172 31340 36204
rect 30968 35928 31032 36172
rect 31276 35928 31340 36172
rect 30968 35896 31340 35928
rect 31968 36172 32340 36204
rect 31968 35928 32032 36172
rect 32276 35928 32340 36172
rect 31968 35896 32340 35928
rect 32968 36172 33340 36204
rect 32968 35928 33032 36172
rect 33276 35928 33340 36172
rect 32968 35896 33340 35928
rect 33968 36172 34340 36204
rect 33968 35928 34032 36172
rect 34276 35928 34340 36172
rect 33968 35896 34340 35928
rect 34648 35896 34654 36204
rect 9654 35890 34654 35896
rect -74485 35864 -74165 35890
rect -74485 35236 -74479 35864
rect -74171 35236 -74165 35864
rect -74485 35210 -74165 35236
rect -73485 35864 -73165 35890
rect -73485 35236 -73479 35864
rect -73171 35236 -73165 35864
rect -73485 35210 -73165 35236
rect -72485 35864 -72165 35890
rect -72485 35236 -72479 35864
rect -72171 35236 -72165 35864
rect -72485 35210 -72165 35236
rect -71485 35864 -71165 35890
rect -71485 35236 -71479 35864
rect -71171 35236 -71165 35864
rect -71485 35210 -71165 35236
rect -70485 35864 -70165 35890
rect -70485 35236 -70479 35864
rect -70171 35236 -70165 35864
rect -70485 35210 -70165 35236
rect -69485 35864 -69165 35890
rect -69485 35236 -69479 35864
rect -69171 35236 -69165 35864
rect -69485 35210 -69165 35236
rect -68485 35864 -68165 35890
rect -68485 35236 -68479 35864
rect -68171 35236 -68165 35864
rect -68485 35210 -68165 35236
rect -67485 35864 -67165 35890
rect -67485 35236 -67479 35864
rect -67171 35236 -67165 35864
rect -67485 35210 -67165 35236
rect -66485 35864 -66165 35890
rect -66485 35236 -66479 35864
rect -66171 35236 -66165 35864
rect -66485 35210 -66165 35236
rect -65485 35864 -65165 35890
rect -65485 35236 -65479 35864
rect -65171 35236 -65165 35864
rect -65485 35210 -65165 35236
rect -64485 35864 -64165 35890
rect -64485 35236 -64479 35864
rect -64171 35236 -64165 35864
rect -64485 35210 -64165 35236
rect -63485 35864 -63165 35890
rect -63485 35236 -63479 35864
rect -63171 35236 -63165 35864
rect -63485 35210 -63165 35236
rect -62485 35864 -62165 35890
rect -62485 35236 -62479 35864
rect -62171 35236 -62165 35864
rect -62485 35210 -62165 35236
rect -61485 35864 -61165 35890
rect -61485 35236 -61479 35864
rect -61171 35236 -61165 35864
rect -61485 35210 -61165 35236
rect -60485 35864 -60165 35890
rect -60485 35236 -60479 35864
rect -60171 35236 -60165 35864
rect -60485 35210 -60165 35236
rect -59485 35864 -59165 35890
rect -59485 35236 -59479 35864
rect -59171 35236 -59165 35864
rect -59485 35210 -59165 35236
rect 9994 35864 10314 35890
rect 9994 35236 10000 35864
rect 10308 35236 10314 35864
rect 9994 35210 10314 35236
rect 10994 35864 11314 35890
rect 10994 35236 11000 35864
rect 11308 35236 11314 35864
rect 10994 35210 11314 35236
rect 11994 35864 12314 35890
rect 11994 35236 12000 35864
rect 12308 35236 12314 35864
rect 11994 35210 12314 35236
rect 12994 35864 13314 35890
rect 12994 35236 13000 35864
rect 13308 35236 13314 35864
rect 12994 35210 13314 35236
rect 13994 35864 14314 35890
rect 13994 35236 14000 35864
rect 14308 35236 14314 35864
rect 13994 35210 14314 35236
rect 14994 35864 15314 35890
rect 14994 35236 15000 35864
rect 15308 35236 15314 35864
rect 14994 35210 15314 35236
rect 15994 35864 16314 35890
rect 15994 35236 16000 35864
rect 16308 35236 16314 35864
rect 15994 35210 16314 35236
rect 16994 35864 17314 35890
rect 16994 35236 17000 35864
rect 17308 35236 17314 35864
rect 16994 35210 17314 35236
rect 17994 35864 18314 35890
rect 17994 35236 18000 35864
rect 18308 35236 18314 35864
rect 17994 35210 18314 35236
rect 18994 35864 19314 35890
rect 18994 35236 19000 35864
rect 19308 35236 19314 35864
rect 18994 35210 19314 35236
rect 19994 35864 20314 35890
rect 19994 35236 20000 35864
rect 20308 35236 20314 35864
rect 19994 35210 20314 35236
rect 20994 35864 21314 35890
rect 20994 35236 21000 35864
rect 21308 35236 21314 35864
rect 20994 35210 21314 35236
rect 21994 35864 22314 35890
rect 21994 35236 22000 35864
rect 22308 35236 22314 35864
rect 21994 35210 22314 35236
rect 22994 35864 23314 35890
rect 22994 35236 23000 35864
rect 23308 35236 23314 35864
rect 22994 35210 23314 35236
rect 23994 35864 24314 35890
rect 23994 35236 24000 35864
rect 24308 35236 24314 35864
rect 23994 35210 24314 35236
rect 24994 35864 25314 35890
rect 24994 35236 25000 35864
rect 25308 35236 25314 35864
rect 24994 35210 25314 35236
rect 25994 35864 26314 35890
rect 25994 35236 26000 35864
rect 26308 35236 26314 35864
rect 25994 35210 26314 35236
rect 26994 35864 27314 35890
rect 26994 35236 27000 35864
rect 27308 35236 27314 35864
rect 26994 35210 27314 35236
rect 27994 35864 28314 35890
rect 27994 35236 28000 35864
rect 28308 35236 28314 35864
rect 27994 35210 28314 35236
rect 28994 35864 29314 35890
rect 28994 35236 29000 35864
rect 29308 35236 29314 35864
rect 28994 35210 29314 35236
rect 29994 35864 30314 35890
rect 29994 35236 30000 35864
rect 30308 35236 30314 35864
rect 29994 35210 30314 35236
rect 30994 35864 31314 35890
rect 30994 35236 31000 35864
rect 31308 35236 31314 35864
rect 30994 35210 31314 35236
rect 31994 35864 32314 35890
rect 31994 35236 32000 35864
rect 32308 35236 32314 35864
rect 31994 35210 32314 35236
rect 32994 35864 33314 35890
rect 32994 35236 33000 35864
rect 33308 35236 33314 35864
rect 32994 35210 33314 35236
rect 33994 35864 34314 35890
rect 33994 35236 34000 35864
rect 34308 35236 34314 35864
rect 33994 35210 34314 35236
rect -74825 35204 -58825 35210
rect -74825 34896 -74819 35204
rect -74511 35172 -74139 35204
rect -74511 34928 -74447 35172
rect -74203 34928 -74139 35172
rect -74511 34896 -74139 34928
rect -73511 35172 -73139 35204
rect -73511 34928 -73447 35172
rect -73203 34928 -73139 35172
rect -73511 34896 -73139 34928
rect -72511 35172 -72139 35204
rect -72511 34928 -72447 35172
rect -72203 34928 -72139 35172
rect -72511 34896 -72139 34928
rect -71511 35172 -71139 35204
rect -71511 34928 -71447 35172
rect -71203 34928 -71139 35172
rect -71511 34896 -71139 34928
rect -70511 35172 -70139 35204
rect -70511 34928 -70447 35172
rect -70203 34928 -70139 35172
rect -70511 34896 -70139 34928
rect -69511 35172 -69139 35204
rect -69511 34928 -69447 35172
rect -69203 34928 -69139 35172
rect -69511 34896 -69139 34928
rect -68511 35172 -68139 35204
rect -68511 34928 -68447 35172
rect -68203 34928 -68139 35172
rect -68511 34896 -68139 34928
rect -67511 35172 -67139 35204
rect -67511 34928 -67447 35172
rect -67203 34928 -67139 35172
rect -67511 34896 -67139 34928
rect -66511 35172 -66139 35204
rect -66511 34928 -66447 35172
rect -66203 34928 -66139 35172
rect -66511 34896 -66139 34928
rect -65511 35172 -65139 35204
rect -65511 34928 -65447 35172
rect -65203 34928 -65139 35172
rect -65511 34896 -65139 34928
rect -64511 35172 -64139 35204
rect -64511 34928 -64447 35172
rect -64203 34928 -64139 35172
rect -64511 34896 -64139 34928
rect -63511 35172 -63139 35204
rect -63511 34928 -63447 35172
rect -63203 34928 -63139 35172
rect -63511 34896 -63139 34928
rect -62511 35172 -62139 35204
rect -62511 34928 -62447 35172
rect -62203 34928 -62139 35172
rect -62511 34896 -62139 34928
rect -61511 35172 -61139 35204
rect -61511 34928 -61447 35172
rect -61203 34928 -61139 35172
rect -61511 34896 -61139 34928
rect -60511 35172 -60139 35204
rect -60511 34928 -60447 35172
rect -60203 34928 -60139 35172
rect -60511 34896 -60139 34928
rect -59511 35172 -59139 35204
rect -59511 34928 -59447 35172
rect -59203 34928 -59139 35172
rect -59511 34896 -59139 34928
rect -58831 34896 -58825 35204
rect -74825 34890 -58825 34896
rect 9654 35204 34654 35210
rect 9654 34896 9660 35204
rect 9968 35172 10340 35204
rect 9968 34928 10032 35172
rect 10276 34928 10340 35172
rect 9968 34896 10340 34928
rect 10968 35172 11340 35204
rect 10968 34928 11032 35172
rect 11276 34928 11340 35172
rect 10968 34896 11340 34928
rect 11968 35172 12340 35204
rect 11968 34928 12032 35172
rect 12276 34928 12340 35172
rect 11968 34896 12340 34928
rect 12968 35172 13340 35204
rect 12968 34928 13032 35172
rect 13276 34928 13340 35172
rect 12968 34896 13340 34928
rect 13968 35172 14340 35204
rect 13968 34928 14032 35172
rect 14276 34928 14340 35172
rect 13968 34896 14340 34928
rect 14968 35172 15340 35204
rect 14968 34928 15032 35172
rect 15276 34928 15340 35172
rect 14968 34896 15340 34928
rect 15968 35172 16340 35204
rect 15968 34928 16032 35172
rect 16276 34928 16340 35172
rect 15968 34896 16340 34928
rect 16968 35172 17340 35204
rect 16968 34928 17032 35172
rect 17276 34928 17340 35172
rect 16968 34896 17340 34928
rect 17968 35172 18340 35204
rect 17968 34928 18032 35172
rect 18276 34928 18340 35172
rect 17968 34896 18340 34928
rect 18968 35172 19340 35204
rect 18968 34928 19032 35172
rect 19276 34928 19340 35172
rect 18968 34896 19340 34928
rect 19968 35172 20340 35204
rect 19968 34928 20032 35172
rect 20276 34928 20340 35172
rect 19968 34896 20340 34928
rect 20968 35172 21340 35204
rect 20968 34928 21032 35172
rect 21276 34928 21340 35172
rect 20968 34896 21340 34928
rect 21968 35172 22340 35204
rect 21968 34928 22032 35172
rect 22276 34928 22340 35172
rect 21968 34896 22340 34928
rect 22968 35172 23340 35204
rect 22968 34928 23032 35172
rect 23276 34928 23340 35172
rect 22968 34896 23340 34928
rect 23968 35172 24340 35204
rect 23968 34928 24032 35172
rect 24276 34928 24340 35172
rect 23968 34896 24340 34928
rect 24968 35172 25340 35204
rect 24968 34928 25032 35172
rect 25276 34928 25340 35172
rect 24968 34896 25340 34928
rect 25968 35172 26340 35204
rect 25968 34928 26032 35172
rect 26276 34928 26340 35172
rect 25968 34896 26340 34928
rect 26968 35172 27340 35204
rect 26968 34928 27032 35172
rect 27276 34928 27340 35172
rect 26968 34896 27340 34928
rect 27968 35172 28340 35204
rect 27968 34928 28032 35172
rect 28276 34928 28340 35172
rect 27968 34896 28340 34928
rect 28968 35172 29340 35204
rect 28968 34928 29032 35172
rect 29276 34928 29340 35172
rect 28968 34896 29340 34928
rect 29968 35172 30340 35204
rect 29968 34928 30032 35172
rect 30276 34928 30340 35172
rect 29968 34896 30340 34928
rect 30968 35172 31340 35204
rect 30968 34928 31032 35172
rect 31276 34928 31340 35172
rect 30968 34896 31340 34928
rect 31968 35172 32340 35204
rect 31968 34928 32032 35172
rect 32276 34928 32340 35172
rect 31968 34896 32340 34928
rect 32968 35172 33340 35204
rect 32968 34928 33032 35172
rect 33276 34928 33340 35172
rect 32968 34896 33340 34928
rect 33968 35172 34340 35204
rect 33968 34928 34032 35172
rect 34276 34928 34340 35172
rect 33968 34896 34340 34928
rect 34648 34896 34654 35204
rect 9654 34890 34654 34896
rect -74485 34864 -74165 34890
rect -74485 34236 -74479 34864
rect -74171 34236 -74165 34864
rect -74485 34210 -74165 34236
rect -73485 34864 -73165 34890
rect -73485 34236 -73479 34864
rect -73171 34236 -73165 34864
rect -73485 34210 -73165 34236
rect -72485 34864 -72165 34890
rect -72485 34236 -72479 34864
rect -72171 34236 -72165 34864
rect -72485 34210 -72165 34236
rect -71485 34864 -71165 34890
rect -71485 34236 -71479 34864
rect -71171 34236 -71165 34864
rect -71485 34210 -71165 34236
rect -70485 34864 -70165 34890
rect -70485 34236 -70479 34864
rect -70171 34236 -70165 34864
rect -70485 34210 -70165 34236
rect -69485 34864 -69165 34890
rect -69485 34236 -69479 34864
rect -69171 34236 -69165 34864
rect -69485 34210 -69165 34236
rect -68485 34864 -68165 34890
rect -68485 34236 -68479 34864
rect -68171 34236 -68165 34864
rect -68485 34210 -68165 34236
rect -67485 34864 -67165 34890
rect -67485 34236 -67479 34864
rect -67171 34236 -67165 34864
rect -67485 34210 -67165 34236
rect -66485 34864 -66165 34890
rect -66485 34236 -66479 34864
rect -66171 34236 -66165 34864
rect -66485 34210 -66165 34236
rect -65485 34864 -65165 34890
rect -65485 34236 -65479 34864
rect -65171 34236 -65165 34864
rect -65485 34210 -65165 34236
rect -64485 34864 -64165 34890
rect -64485 34236 -64479 34864
rect -64171 34236 -64165 34864
rect -64485 34210 -64165 34236
rect -63485 34864 -63165 34890
rect -63485 34236 -63479 34864
rect -63171 34236 -63165 34864
rect -63485 34210 -63165 34236
rect -62485 34864 -62165 34890
rect -62485 34236 -62479 34864
rect -62171 34236 -62165 34864
rect -62485 34210 -62165 34236
rect -61485 34864 -61165 34890
rect -61485 34236 -61479 34864
rect -61171 34236 -61165 34864
rect -61485 34210 -61165 34236
rect -60485 34864 -60165 34890
rect -60485 34236 -60479 34864
rect -60171 34236 -60165 34864
rect -60485 34210 -60165 34236
rect -59485 34864 -59165 34890
rect -59485 34236 -59479 34864
rect -59171 34236 -59165 34864
rect -59485 34210 -59165 34236
rect 9994 34864 10314 34890
rect 9994 34236 10000 34864
rect 10308 34236 10314 34864
rect 9994 34210 10314 34236
rect 10994 34864 11314 34890
rect 10994 34236 11000 34864
rect 11308 34236 11314 34864
rect 10994 34210 11314 34236
rect 11994 34864 12314 34890
rect 11994 34236 12000 34864
rect 12308 34236 12314 34864
rect 11994 34210 12314 34236
rect 12994 34864 13314 34890
rect 12994 34236 13000 34864
rect 13308 34236 13314 34864
rect 12994 34210 13314 34236
rect 13994 34864 14314 34890
rect 13994 34236 14000 34864
rect 14308 34236 14314 34864
rect 13994 34210 14314 34236
rect 14994 34864 15314 34890
rect 14994 34236 15000 34864
rect 15308 34236 15314 34864
rect 14994 34210 15314 34236
rect 15994 34864 16314 34890
rect 15994 34236 16000 34864
rect 16308 34236 16314 34864
rect 15994 34210 16314 34236
rect 16994 34864 17314 34890
rect 16994 34236 17000 34864
rect 17308 34236 17314 34864
rect 16994 34210 17314 34236
rect 17994 34864 18314 34890
rect 17994 34236 18000 34864
rect 18308 34236 18314 34864
rect 17994 34210 18314 34236
rect 18994 34864 19314 34890
rect 18994 34236 19000 34864
rect 19308 34236 19314 34864
rect 18994 34210 19314 34236
rect 19994 34864 20314 34890
rect 19994 34236 20000 34864
rect 20308 34236 20314 34864
rect 19994 34210 20314 34236
rect 20994 34864 21314 34890
rect 20994 34236 21000 34864
rect 21308 34236 21314 34864
rect 20994 34210 21314 34236
rect 21994 34864 22314 34890
rect 21994 34236 22000 34864
rect 22308 34236 22314 34864
rect 21994 34210 22314 34236
rect 22994 34864 23314 34890
rect 22994 34236 23000 34864
rect 23308 34236 23314 34864
rect 22994 34210 23314 34236
rect 23994 34864 24314 34890
rect 23994 34236 24000 34864
rect 24308 34236 24314 34864
rect 23994 34210 24314 34236
rect 24994 34864 25314 34890
rect 24994 34236 25000 34864
rect 25308 34236 25314 34864
rect 24994 34210 25314 34236
rect 25994 34864 26314 34890
rect 25994 34236 26000 34864
rect 26308 34236 26314 34864
rect 25994 34210 26314 34236
rect 26994 34864 27314 34890
rect 26994 34236 27000 34864
rect 27308 34236 27314 34864
rect 26994 34210 27314 34236
rect 27994 34864 28314 34890
rect 27994 34236 28000 34864
rect 28308 34236 28314 34864
rect 27994 34210 28314 34236
rect 28994 34864 29314 34890
rect 28994 34236 29000 34864
rect 29308 34236 29314 34864
rect 28994 34210 29314 34236
rect 29994 34864 30314 34890
rect 29994 34236 30000 34864
rect 30308 34236 30314 34864
rect 29994 34210 30314 34236
rect 30994 34864 31314 34890
rect 30994 34236 31000 34864
rect 31308 34236 31314 34864
rect 30994 34210 31314 34236
rect 31994 34864 32314 34890
rect 31994 34236 32000 34864
rect 32308 34236 32314 34864
rect 31994 34210 32314 34236
rect 32994 34864 33314 34890
rect 32994 34236 33000 34864
rect 33308 34236 33314 34864
rect 32994 34210 33314 34236
rect 33994 34864 34314 34890
rect 33994 34236 34000 34864
rect 34308 34236 34314 34864
rect 33994 34210 34314 34236
rect -74825 34204 -58825 34210
rect -74825 33896 -74819 34204
rect -74511 34172 -74139 34204
rect -74511 33928 -74447 34172
rect -74203 33928 -74139 34172
rect -74511 33896 -74139 33928
rect -73511 34172 -73139 34204
rect -73511 33928 -73447 34172
rect -73203 33928 -73139 34172
rect -73511 33896 -73139 33928
rect -72511 34172 -72139 34204
rect -72511 33928 -72447 34172
rect -72203 33928 -72139 34172
rect -72511 33896 -72139 33928
rect -71511 34172 -71139 34204
rect -71511 33928 -71447 34172
rect -71203 33928 -71139 34172
rect -71511 33896 -71139 33928
rect -70511 34172 -70139 34204
rect -70511 33928 -70447 34172
rect -70203 33928 -70139 34172
rect -70511 33896 -70139 33928
rect -69511 34172 -69139 34204
rect -69511 33928 -69447 34172
rect -69203 33928 -69139 34172
rect -69511 33896 -69139 33928
rect -68511 34172 -68139 34204
rect -68511 33928 -68447 34172
rect -68203 33928 -68139 34172
rect -68511 33896 -68139 33928
rect -67511 34172 -67139 34204
rect -67511 33928 -67447 34172
rect -67203 33928 -67139 34172
rect -67511 33896 -67139 33928
rect -66511 34172 -66139 34204
rect -66511 33928 -66447 34172
rect -66203 33928 -66139 34172
rect -66511 33896 -66139 33928
rect -65511 34172 -65139 34204
rect -65511 33928 -65447 34172
rect -65203 33928 -65139 34172
rect -65511 33896 -65139 33928
rect -64511 34172 -64139 34204
rect -64511 33928 -64447 34172
rect -64203 33928 -64139 34172
rect -64511 33896 -64139 33928
rect -63511 34172 -63139 34204
rect -63511 33928 -63447 34172
rect -63203 33928 -63139 34172
rect -63511 33896 -63139 33928
rect -62511 34172 -62139 34204
rect -62511 33928 -62447 34172
rect -62203 33928 -62139 34172
rect -62511 33896 -62139 33928
rect -61511 34172 -61139 34204
rect -61511 33928 -61447 34172
rect -61203 33928 -61139 34172
rect -61511 33896 -61139 33928
rect -60511 34172 -60139 34204
rect -60511 33928 -60447 34172
rect -60203 33928 -60139 34172
rect -60511 33896 -60139 33928
rect -59511 34172 -59139 34204
rect -59511 33928 -59447 34172
rect -59203 33928 -59139 34172
rect -59511 33896 -59139 33928
rect -58831 33896 -58825 34204
rect 9654 34204 34654 34210
rect -74825 33890 -58825 33896
rect -50472 34170 -48808 34176
rect -74485 33864 -74165 33890
rect -74485 33236 -74479 33864
rect -74171 33236 -74165 33864
rect -74485 33210 -74165 33236
rect -73485 33864 -73165 33890
rect -73485 33236 -73479 33864
rect -73171 33236 -73165 33864
rect -73485 33210 -73165 33236
rect -72485 33864 -72165 33890
rect -72485 33236 -72479 33864
rect -72171 33236 -72165 33864
rect -72485 33210 -72165 33236
rect -71485 33864 -71165 33890
rect -71485 33236 -71479 33864
rect -71171 33236 -71165 33864
rect -71485 33210 -71165 33236
rect -70485 33864 -70165 33890
rect -70485 33236 -70479 33864
rect -70171 33236 -70165 33864
rect -70485 33210 -70165 33236
rect -69485 33864 -69165 33890
rect -69485 33236 -69479 33864
rect -69171 33236 -69165 33864
rect -69485 33210 -69165 33236
rect -68485 33864 -68165 33890
rect -68485 33236 -68479 33864
rect -68171 33236 -68165 33864
rect -68485 33210 -68165 33236
rect -67485 33864 -67165 33890
rect -67485 33236 -67479 33864
rect -67171 33236 -67165 33864
rect -67485 33210 -67165 33236
rect -66485 33864 -66165 33890
rect -66485 33236 -66479 33864
rect -66171 33236 -66165 33864
rect -66485 33210 -66165 33236
rect -65485 33864 -65165 33890
rect -65485 33236 -65479 33864
rect -65171 33236 -65165 33864
rect -65485 33210 -65165 33236
rect -64485 33864 -64165 33890
rect -64485 33236 -64479 33864
rect -64171 33236 -64165 33864
rect -64485 33210 -64165 33236
rect -63485 33864 -63165 33890
rect -63485 33236 -63479 33864
rect -63171 33236 -63165 33864
rect -63485 33210 -63165 33236
rect -62485 33864 -62165 33890
rect -62485 33236 -62479 33864
rect -62171 33236 -62165 33864
rect -62485 33210 -62165 33236
rect -61485 33864 -61165 33890
rect -61485 33236 -61479 33864
rect -61171 33236 -61165 33864
rect -61485 33210 -61165 33236
rect -60485 33864 -60165 33890
rect -60485 33236 -60479 33864
rect -60171 33236 -60165 33864
rect -60485 33210 -60165 33236
rect -59485 33864 -59165 33890
rect -59485 33236 -59479 33864
rect -59171 33236 -59165 33864
rect -50472 33542 -50466 34170
rect -48814 33542 -48808 34170
rect -50472 33536 -48808 33542
rect 2875 34170 4539 34176
rect 2875 33542 2881 34170
rect 4533 33542 4539 34170
rect 9654 33896 9660 34204
rect 9968 34172 10340 34204
rect 9968 33928 10032 34172
rect 10276 33928 10340 34172
rect 9968 33896 10340 33928
rect 10968 34172 11340 34204
rect 10968 33928 11032 34172
rect 11276 33928 11340 34172
rect 10968 33896 11340 33928
rect 11968 34172 12340 34204
rect 11968 33928 12032 34172
rect 12276 33928 12340 34172
rect 11968 33896 12340 33928
rect 12968 34172 13340 34204
rect 12968 33928 13032 34172
rect 13276 33928 13340 34172
rect 12968 33896 13340 33928
rect 13968 34172 14340 34204
rect 13968 33928 14032 34172
rect 14276 33928 14340 34172
rect 13968 33896 14340 33928
rect 14968 34172 15340 34204
rect 14968 33928 15032 34172
rect 15276 33928 15340 34172
rect 14968 33896 15340 33928
rect 15968 34172 16340 34204
rect 15968 33928 16032 34172
rect 16276 33928 16340 34172
rect 15968 33896 16340 33928
rect 16968 34172 17340 34204
rect 16968 33928 17032 34172
rect 17276 33928 17340 34172
rect 16968 33896 17340 33928
rect 17968 34172 18340 34204
rect 17968 33928 18032 34172
rect 18276 33928 18340 34172
rect 17968 33896 18340 33928
rect 18968 34172 19340 34204
rect 18968 33928 19032 34172
rect 19276 33928 19340 34172
rect 18968 33896 19340 33928
rect 19968 34172 20340 34204
rect 19968 33928 20032 34172
rect 20276 33928 20340 34172
rect 19968 33896 20340 33928
rect 20968 34172 21340 34204
rect 20968 33928 21032 34172
rect 21276 33928 21340 34172
rect 20968 33896 21340 33928
rect 21968 34172 22340 34204
rect 21968 33928 22032 34172
rect 22276 33928 22340 34172
rect 21968 33896 22340 33928
rect 22968 34172 23340 34204
rect 22968 33928 23032 34172
rect 23276 33928 23340 34172
rect 22968 33896 23340 33928
rect 23968 34172 24340 34204
rect 23968 33928 24032 34172
rect 24276 33928 24340 34172
rect 23968 33896 24340 33928
rect 24968 34172 25340 34204
rect 24968 33928 25032 34172
rect 25276 33928 25340 34172
rect 24968 33896 25340 33928
rect 25968 34172 26340 34204
rect 25968 33928 26032 34172
rect 26276 33928 26340 34172
rect 25968 33896 26340 33928
rect 26968 34172 27340 34204
rect 26968 33928 27032 34172
rect 27276 33928 27340 34172
rect 26968 33896 27340 33928
rect 27968 34172 28340 34204
rect 27968 33928 28032 34172
rect 28276 33928 28340 34172
rect 27968 33896 28340 33928
rect 28968 34172 29340 34204
rect 28968 33928 29032 34172
rect 29276 33928 29340 34172
rect 28968 33896 29340 33928
rect 29968 34172 30340 34204
rect 29968 33928 30032 34172
rect 30276 33928 30340 34172
rect 29968 33896 30340 33928
rect 30968 34172 31340 34204
rect 30968 33928 31032 34172
rect 31276 33928 31340 34172
rect 30968 33896 31340 33928
rect 31968 34172 32340 34204
rect 31968 33928 32032 34172
rect 32276 33928 32340 34172
rect 31968 33896 32340 33928
rect 32968 34172 33340 34204
rect 32968 33928 33032 34172
rect 33276 33928 33340 34172
rect 32968 33896 33340 33928
rect 33968 34172 34340 34204
rect 33968 33928 34032 34172
rect 34276 33928 34340 34172
rect 33968 33896 34340 33928
rect 34648 33896 34654 34204
rect 9654 33890 34654 33896
rect 2875 33536 4539 33542
rect 9994 33864 10314 33890
rect -59485 33210 -59165 33236
rect -50461 33524 -48819 33536
rect -50461 33418 -50449 33524
rect -48831 33418 -48819 33524
rect -50461 33406 -48819 33418
rect -50461 33273 -50407 33406
rect -50295 33304 -50249 33312
rect -50461 33239 -50447 33273
rect -50413 33239 -50407 33273
rect -74825 33204 -58825 33210
rect -74825 32896 -74819 33204
rect -74511 33172 -74139 33204
rect -74511 32928 -74447 33172
rect -74203 32928 -74139 33172
rect -74511 32896 -74139 32928
rect -73511 33172 -73139 33204
rect -73511 32928 -73447 33172
rect -73203 32928 -73139 33172
rect -73511 32896 -73139 32928
rect -72511 33172 -72139 33204
rect -72511 32928 -72447 33172
rect -72203 32928 -72139 33172
rect -72511 32896 -72139 32928
rect -71511 33172 -71139 33204
rect -71511 32928 -71447 33172
rect -71203 32928 -71139 33172
rect -71511 32896 -71139 32928
rect -70511 33172 -70139 33204
rect -70511 32928 -70447 33172
rect -70203 32928 -70139 33172
rect -70511 32896 -70139 32928
rect -69511 33172 -69139 33204
rect -69511 32928 -69447 33172
rect -69203 32928 -69139 33172
rect -69511 32896 -69139 32928
rect -68511 33172 -68139 33204
rect -68511 32928 -68447 33172
rect -68203 32928 -68139 33172
rect -68511 32896 -68139 32928
rect -67511 33172 -67139 33204
rect -67511 32928 -67447 33172
rect -67203 32928 -67139 33172
rect -67511 32896 -67139 32928
rect -66511 33172 -66139 33204
rect -66511 32928 -66447 33172
rect -66203 32928 -66139 33172
rect -66511 32896 -66139 32928
rect -65511 33172 -65139 33204
rect -65511 32928 -65447 33172
rect -65203 32928 -65139 33172
rect -65511 32896 -65139 32928
rect -64511 33172 -64139 33204
rect -64511 32928 -64447 33172
rect -64203 32928 -64139 33172
rect -64511 32896 -64139 32928
rect -63511 33172 -63139 33204
rect -63511 32928 -63447 33172
rect -63203 32928 -63139 33172
rect -63511 32896 -63139 32928
rect -62511 33172 -62139 33204
rect -62511 32928 -62447 33172
rect -62203 32928 -62139 33172
rect -62511 32896 -62139 32928
rect -61511 33172 -61139 33204
rect -61511 32928 -61447 33172
rect -61203 32928 -61139 33172
rect -61511 32896 -61139 32928
rect -60511 33172 -60139 33204
rect -60511 32928 -60447 33172
rect -60203 32928 -60139 33172
rect -60511 32896 -60139 32928
rect -59511 33172 -59139 33204
rect -59511 32928 -59447 33172
rect -59203 32928 -59139 33172
rect -59511 32896 -59139 32928
rect -58831 32896 -58825 33204
rect -50461 33201 -50407 33239
rect -50461 33167 -50447 33201
rect -50413 33167 -50407 33201
rect -50461 33129 -50407 33167
rect -50461 33095 -50447 33129
rect -50413 33095 -50407 33129
rect -50461 33057 -50407 33095
rect -50461 33023 -50447 33057
rect -50413 33023 -50407 33057
rect -50461 32985 -50407 33023
rect -74825 32890 -58825 32896
rect -50957 32965 -50573 32971
rect -74485 32864 -74165 32890
rect -74485 32236 -74479 32864
rect -74171 32236 -74165 32864
rect -74485 32210 -74165 32236
rect -73485 32864 -73165 32890
rect -73485 32236 -73479 32864
rect -73171 32236 -73165 32864
rect -73485 32210 -73165 32236
rect -72485 32864 -72165 32890
rect -72485 32236 -72479 32864
rect -72171 32236 -72165 32864
rect -72485 32210 -72165 32236
rect -71485 32864 -71165 32890
rect -71485 32236 -71479 32864
rect -71171 32236 -71165 32864
rect -71485 32210 -71165 32236
rect -70485 32864 -70165 32890
rect -70485 32236 -70479 32864
rect -70171 32236 -70165 32864
rect -70485 32210 -70165 32236
rect -69485 32864 -69165 32890
rect -69485 32236 -69479 32864
rect -69171 32236 -69165 32864
rect -69485 32210 -69165 32236
rect -68485 32864 -68165 32890
rect -68485 32236 -68479 32864
rect -68171 32236 -68165 32864
rect -68485 32210 -68165 32236
rect -67485 32864 -67165 32890
rect -67485 32236 -67479 32864
rect -67171 32236 -67165 32864
rect -67485 32210 -67165 32236
rect -66485 32864 -66165 32890
rect -66485 32236 -66479 32864
rect -66171 32236 -66165 32864
rect -66485 32210 -66165 32236
rect -65485 32864 -65165 32890
rect -65485 32236 -65479 32864
rect -65171 32236 -65165 32864
rect -65485 32210 -65165 32236
rect -64485 32864 -64165 32890
rect -64485 32236 -64479 32864
rect -64171 32236 -64165 32864
rect -64485 32210 -64165 32236
rect -63485 32864 -63165 32890
rect -63485 32236 -63479 32864
rect -63171 32236 -63165 32864
rect -63485 32210 -63165 32236
rect -62485 32864 -62165 32890
rect -62485 32236 -62479 32864
rect -62171 32236 -62165 32864
rect -62485 32210 -62165 32236
rect -61485 32864 -61165 32890
rect -61485 32236 -61479 32864
rect -61171 32236 -61165 32864
rect -61485 32210 -61165 32236
rect -60485 32864 -60165 32890
rect -60485 32236 -60479 32864
rect -60171 32236 -60165 32864
rect -60485 32210 -60165 32236
rect -59485 32864 -59165 32890
rect -59485 32236 -59479 32864
rect -59171 32236 -59165 32864
rect -50957 32593 -50951 32965
rect -50579 32593 -50573 32965
rect -50461 32951 -50447 32985
rect -50413 32951 -50407 32985
rect -50461 32912 -50407 32951
rect -50304 33298 -50240 33304
rect -50304 33246 -50298 33298
rect -50246 33246 -50240 33298
rect -50304 33239 -50289 33246
rect -50255 33239 -50240 33246
rect -50304 33234 -50240 33239
rect -50304 33182 -50298 33234
rect -50246 33182 -50240 33234
rect -50304 33170 -50289 33182
rect -50255 33170 -50240 33182
rect -50304 33118 -50298 33170
rect -50246 33118 -50240 33170
rect -50304 33106 -50289 33118
rect -50255 33106 -50240 33118
rect -50304 33054 -50298 33106
rect -50246 33054 -50240 33106
rect -50304 33042 -50289 33054
rect -50255 33042 -50240 33054
rect -50304 32990 -50298 33042
rect -50246 32990 -50240 33042
rect -50304 32985 -50240 32990
rect -50304 32978 -50289 32985
rect -50255 32978 -50240 32985
rect -50304 32926 -50298 32978
rect -50246 32926 -50240 32978
rect -50304 32920 -50240 32926
rect -50137 33273 -50091 33406
rect -49979 33304 -49933 33312
rect -50137 33239 -50131 33273
rect -50097 33239 -50091 33273
rect -50137 33201 -50091 33239
rect -50137 33167 -50131 33201
rect -50097 33167 -50091 33201
rect -50137 33129 -50091 33167
rect -50137 33095 -50131 33129
rect -50097 33095 -50091 33129
rect -50137 33057 -50091 33095
rect -50137 33023 -50131 33057
rect -50097 33023 -50091 33057
rect -50137 32985 -50091 33023
rect -50137 32951 -50131 32985
rect -50097 32951 -50091 32985
rect -50295 32912 -50249 32920
rect -50137 32912 -50091 32951
rect -49988 33298 -49924 33304
rect -49988 33246 -49982 33298
rect -49930 33246 -49924 33298
rect -49988 33239 -49973 33246
rect -49939 33239 -49924 33246
rect -49988 33234 -49924 33239
rect -49988 33182 -49982 33234
rect -49930 33182 -49924 33234
rect -49988 33170 -49973 33182
rect -49939 33170 -49924 33182
rect -49988 33118 -49982 33170
rect -49930 33118 -49924 33170
rect -49988 33106 -49973 33118
rect -49939 33106 -49924 33118
rect -49988 33054 -49982 33106
rect -49930 33054 -49924 33106
rect -49988 33042 -49973 33054
rect -49939 33042 -49924 33054
rect -49988 32990 -49982 33042
rect -49930 32990 -49924 33042
rect -49988 32985 -49924 32990
rect -49988 32978 -49973 32985
rect -49939 32978 -49924 32985
rect -49988 32926 -49982 32978
rect -49930 32926 -49924 32978
rect -49988 32920 -49924 32926
rect -49821 33273 -49775 33406
rect -49663 33304 -49617 33312
rect -49821 33239 -49815 33273
rect -49781 33239 -49775 33273
rect -49821 33201 -49775 33239
rect -49821 33167 -49815 33201
rect -49781 33167 -49775 33201
rect -49821 33129 -49775 33167
rect -49821 33095 -49815 33129
rect -49781 33095 -49775 33129
rect -49821 33057 -49775 33095
rect -49821 33023 -49815 33057
rect -49781 33023 -49775 33057
rect -49821 32985 -49775 33023
rect -49821 32951 -49815 32985
rect -49781 32951 -49775 32985
rect -49979 32912 -49933 32920
rect -49821 32912 -49775 32951
rect -49672 33298 -49608 33304
rect -49672 33246 -49666 33298
rect -49614 33246 -49608 33298
rect -49672 33239 -49657 33246
rect -49623 33239 -49608 33246
rect -49672 33234 -49608 33239
rect -49672 33182 -49666 33234
rect -49614 33182 -49608 33234
rect -49672 33170 -49657 33182
rect -49623 33170 -49608 33182
rect -49672 33118 -49666 33170
rect -49614 33118 -49608 33170
rect -49672 33106 -49657 33118
rect -49623 33106 -49608 33118
rect -49672 33054 -49666 33106
rect -49614 33054 -49608 33106
rect -49672 33042 -49657 33054
rect -49623 33042 -49608 33054
rect -49672 32990 -49666 33042
rect -49614 32990 -49608 33042
rect -49672 32985 -49608 32990
rect -49672 32978 -49657 32985
rect -49623 32978 -49608 32985
rect -49672 32926 -49666 32978
rect -49614 32926 -49608 32978
rect -49672 32920 -49608 32926
rect -49505 33273 -49459 33406
rect -49347 33304 -49301 33312
rect -49505 33239 -49499 33273
rect -49465 33239 -49459 33273
rect -49505 33201 -49459 33239
rect -49505 33167 -49499 33201
rect -49465 33167 -49459 33201
rect -49505 33129 -49459 33167
rect -49505 33095 -49499 33129
rect -49465 33095 -49459 33129
rect -49505 33057 -49459 33095
rect -49505 33023 -49499 33057
rect -49465 33023 -49459 33057
rect -49505 32985 -49459 33023
rect -49505 32951 -49499 32985
rect -49465 32951 -49459 32985
rect -49663 32912 -49617 32920
rect -49505 32912 -49459 32951
rect -49356 33298 -49292 33304
rect -49356 33246 -49350 33298
rect -49298 33246 -49292 33298
rect -49356 33239 -49341 33246
rect -49307 33239 -49292 33246
rect -49356 33234 -49292 33239
rect -49356 33182 -49350 33234
rect -49298 33182 -49292 33234
rect -49356 33170 -49341 33182
rect -49307 33170 -49292 33182
rect -49356 33118 -49350 33170
rect -49298 33118 -49292 33170
rect -49356 33106 -49341 33118
rect -49307 33106 -49292 33118
rect -49356 33054 -49350 33106
rect -49298 33054 -49292 33106
rect -49356 33042 -49341 33054
rect -49307 33042 -49292 33054
rect -49356 32990 -49350 33042
rect -49298 32990 -49292 33042
rect -49356 32985 -49292 32990
rect -49356 32978 -49341 32985
rect -49307 32978 -49292 32985
rect -49356 32926 -49350 32978
rect -49298 32926 -49292 32978
rect -49356 32920 -49292 32926
rect -49189 33273 -49143 33406
rect -49031 33304 -48985 33312
rect -49189 33239 -49183 33273
rect -49149 33239 -49143 33273
rect -49189 33201 -49143 33239
rect -49189 33167 -49183 33201
rect -49149 33167 -49143 33201
rect -49189 33129 -49143 33167
rect -49189 33095 -49183 33129
rect -49149 33095 -49143 33129
rect -49189 33057 -49143 33095
rect -49189 33023 -49183 33057
rect -49149 33023 -49143 33057
rect -49189 32985 -49143 33023
rect -49189 32951 -49183 32985
rect -49149 32951 -49143 32985
rect -49347 32912 -49301 32920
rect -49189 32912 -49143 32951
rect -49040 33298 -48976 33304
rect -49040 33246 -49034 33298
rect -48982 33246 -48976 33298
rect -49040 33239 -49025 33246
rect -48991 33239 -48976 33246
rect -49040 33234 -48976 33239
rect -49040 33182 -49034 33234
rect -48982 33182 -48976 33234
rect -49040 33170 -49025 33182
rect -48991 33170 -48976 33182
rect -49040 33118 -49034 33170
rect -48982 33118 -48976 33170
rect -49040 33106 -49025 33118
rect -48991 33106 -48976 33118
rect -49040 33054 -49034 33106
rect -48982 33054 -48976 33106
rect -49040 33042 -49025 33054
rect -48991 33042 -48976 33054
rect -49040 32990 -49034 33042
rect -48982 32990 -48976 33042
rect -49040 32985 -48976 32990
rect -49040 32978 -49025 32985
rect -48991 32978 -48976 32985
rect -49040 32926 -49034 32978
rect -48982 32926 -48976 32978
rect -49040 32920 -48976 32926
rect -48873 33273 -48819 33406
rect -48873 33239 -48867 33273
rect -48833 33239 -48819 33273
rect -48873 33201 -48819 33239
rect -48873 33167 -48867 33201
rect -48833 33167 -48819 33201
rect -48873 33129 -48819 33167
rect -48873 33095 -48867 33129
rect -48833 33095 -48819 33129
rect -48873 33057 -48819 33095
rect -48873 33023 -48867 33057
rect -48833 33023 -48819 33057
rect -48873 32985 -48819 33023
rect -48873 32951 -48867 32985
rect -48833 32951 -48819 32985
rect 2886 33524 4528 33536
rect 2886 33418 2898 33524
rect 4516 33418 4528 33524
rect 2886 33406 4528 33418
rect 2886 33273 2940 33406
rect 3052 33304 3098 33312
rect 2886 33239 2900 33273
rect 2934 33239 2940 33273
rect 2886 33201 2940 33239
rect 2886 33167 2900 33201
rect 2934 33167 2940 33201
rect 2886 33129 2940 33167
rect 2886 33095 2900 33129
rect 2934 33095 2940 33129
rect 2886 33057 2940 33095
rect 2886 33023 2900 33057
rect 2934 33023 2940 33057
rect 2886 32985 2940 33023
rect -49031 32912 -48985 32920
rect -48873 32912 -48819 32951
rect 2390 32965 2774 32971
rect -50397 32865 -50305 32871
rect -50397 32831 -50368 32865
rect -50334 32831 -50305 32865
rect -50397 32825 -50305 32831
rect -50239 32865 -50147 32871
rect -50239 32831 -50210 32865
rect -50176 32831 -50147 32865
rect -50239 32825 -50147 32831
rect -50081 32865 -49989 32871
rect -50081 32831 -50052 32865
rect -50018 32831 -49989 32865
rect -50081 32825 -49989 32831
rect -49923 32865 -49831 32871
rect -49923 32831 -49894 32865
rect -49860 32831 -49831 32865
rect -49923 32825 -49831 32831
rect -49765 32865 -49673 32871
rect -49765 32831 -49736 32865
rect -49702 32831 -49673 32865
rect -49765 32825 -49673 32831
rect -49607 32865 -49515 32871
rect -49607 32831 -49578 32865
rect -49544 32831 -49515 32865
rect -49607 32825 -49515 32831
rect -49449 32865 -49357 32871
rect -49449 32831 -49420 32865
rect -49386 32831 -49357 32865
rect -49449 32825 -49357 32831
rect -49291 32865 -49199 32871
rect -49291 32831 -49262 32865
rect -49228 32831 -49199 32865
rect -49291 32825 -49199 32831
rect -49133 32865 -49041 32871
rect -49133 32831 -49104 32865
rect -49070 32831 -49041 32865
rect -49133 32825 -49041 32831
rect -48975 32865 -48883 32871
rect -48975 32831 -48946 32865
rect -48912 32831 -48883 32865
rect -48975 32825 -48883 32831
rect -50397 32727 -50305 32733
rect -50397 32693 -50368 32727
rect -50334 32693 -50305 32727
rect -50397 32687 -50305 32693
rect -50239 32727 -50147 32733
rect -50239 32693 -50210 32727
rect -50176 32693 -50147 32727
rect -50239 32687 -50147 32693
rect -50081 32727 -49989 32733
rect -50081 32693 -50052 32727
rect -50018 32693 -49989 32727
rect -50081 32687 -49989 32693
rect -49923 32727 -49831 32733
rect -49923 32693 -49894 32727
rect -49860 32693 -49831 32727
rect -49923 32687 -49831 32693
rect -49765 32727 -49673 32733
rect -49765 32693 -49736 32727
rect -49702 32693 -49673 32727
rect -49765 32687 -49673 32693
rect -49607 32727 -49515 32733
rect -49607 32693 -49578 32727
rect -49544 32693 -49515 32727
rect -49607 32687 -49515 32693
rect -49449 32727 -49357 32733
rect -49449 32693 -49420 32727
rect -49386 32693 -49357 32727
rect -49449 32687 -49357 32693
rect -49291 32727 -49199 32733
rect -49291 32693 -49262 32727
rect -49228 32693 -49199 32727
rect -49291 32687 -49199 32693
rect -49133 32727 -49041 32733
rect -49133 32693 -49104 32727
rect -49070 32693 -49041 32727
rect -49133 32687 -49041 32693
rect -48975 32727 -48883 32733
rect -48975 32693 -48946 32727
rect -48912 32693 -48883 32727
rect -48975 32687 -48883 32693
rect 2390 32657 2396 32965
rect -50957 32587 -50573 32593
rect -50461 32608 -50407 32655
rect -50295 32651 -50249 32655
rect -59485 32210 -59165 32236
rect -74825 32204 -58825 32210
rect -74825 31896 -74819 32204
rect -74511 32172 -74139 32204
rect -74511 31928 -74447 32172
rect -74203 31928 -74139 32172
rect -74511 31896 -74139 31928
rect -73511 32172 -73139 32204
rect -73511 31928 -73447 32172
rect -73203 31928 -73139 32172
rect -73511 31896 -73139 31928
rect -72511 32172 -72139 32204
rect -72511 31928 -72447 32172
rect -72203 31928 -72139 32172
rect -72511 31896 -72139 31928
rect -71511 32172 -71139 32204
rect -71511 31928 -71447 32172
rect -71203 31928 -71139 32172
rect -71511 31896 -71139 31928
rect -70511 32172 -70139 32204
rect -70511 31928 -70447 32172
rect -70203 31928 -70139 32172
rect -70511 31896 -70139 31928
rect -69511 32172 -69139 32204
rect -69511 31928 -69447 32172
rect -69203 31928 -69139 32172
rect -69511 31896 -69139 31928
rect -68511 32172 -68139 32204
rect -68511 31928 -68447 32172
rect -68203 31928 -68139 32172
rect -68511 31896 -68139 31928
rect -67511 32172 -67139 32204
rect -67511 31928 -67447 32172
rect -67203 31928 -67139 32172
rect -67511 31896 -67139 31928
rect -66511 32172 -66139 32204
rect -66511 31928 -66447 32172
rect -66203 31928 -66139 32172
rect -66511 31896 -66139 31928
rect -65511 32172 -65139 32204
rect -65511 31928 -65447 32172
rect -65203 31928 -65139 32172
rect -65511 31896 -65139 31928
rect -64511 32172 -64139 32204
rect -64511 31928 -64447 32172
rect -64203 31928 -64139 32172
rect -64511 31896 -64139 31928
rect -63511 32172 -63139 32204
rect -63511 31928 -63447 32172
rect -63203 31928 -63139 32172
rect -63511 31896 -63139 31928
rect -62511 32172 -62139 32204
rect -62511 31928 -62447 32172
rect -62203 31928 -62139 32172
rect -62511 31896 -62139 31928
rect -61511 32172 -61139 32204
rect -61511 31928 -61447 32172
rect -61203 31928 -61139 32172
rect -61511 31896 -61139 31928
rect -60511 32172 -60139 32204
rect -60511 31928 -60447 32172
rect -60203 31928 -60139 32172
rect -60511 31896 -60139 31928
rect -59511 32172 -59139 32204
rect -59511 31928 -59447 32172
rect -59203 31928 -59139 32172
rect -59511 31896 -59139 31928
rect -58831 31896 -58825 32204
rect -50797 32035 -50707 32587
rect -50461 32574 -50447 32608
rect -50413 32574 -50407 32608
rect -50461 32536 -50407 32574
rect -50461 32502 -50447 32536
rect -50413 32502 -50407 32536
rect -50461 32361 -50407 32502
rect -50304 32645 -50240 32651
rect -50304 32593 -50298 32645
rect -50246 32593 -50240 32645
rect -50304 32581 -50289 32593
rect -50255 32581 -50240 32593
rect -50304 32529 -50298 32581
rect -50246 32529 -50240 32581
rect -50304 32517 -50289 32529
rect -50255 32517 -50240 32529
rect -50304 32465 -50298 32517
rect -50246 32465 -50240 32517
rect -50304 32459 -50240 32465
rect -50137 32608 -50091 32655
rect -49979 32651 -49933 32655
rect -50137 32574 -50131 32608
rect -50097 32574 -50091 32608
rect -50137 32536 -50091 32574
rect -50137 32502 -50131 32536
rect -50097 32502 -50091 32536
rect -50295 32455 -50249 32459
rect -50137 32361 -50091 32502
rect -49988 32645 -49924 32651
rect -49988 32593 -49982 32645
rect -49930 32593 -49924 32645
rect -49988 32581 -49973 32593
rect -49939 32581 -49924 32593
rect -49988 32529 -49982 32581
rect -49930 32529 -49924 32581
rect -49988 32517 -49973 32529
rect -49939 32517 -49924 32529
rect -49988 32465 -49982 32517
rect -49930 32465 -49924 32517
rect -49988 32459 -49924 32465
rect -49821 32608 -49775 32655
rect -49663 32651 -49617 32655
rect -49821 32574 -49815 32608
rect -49781 32574 -49775 32608
rect -49821 32536 -49775 32574
rect -49821 32502 -49815 32536
rect -49781 32502 -49775 32536
rect -49979 32455 -49933 32459
rect -49821 32361 -49775 32502
rect -49672 32645 -49608 32651
rect -49672 32593 -49666 32645
rect -49614 32593 -49608 32645
rect -49672 32581 -49657 32593
rect -49623 32581 -49608 32593
rect -49672 32529 -49666 32581
rect -49614 32529 -49608 32581
rect -49672 32517 -49657 32529
rect -49623 32517 -49608 32529
rect -49672 32465 -49666 32517
rect -49614 32465 -49608 32517
rect -49672 32459 -49608 32465
rect -49505 32608 -49459 32655
rect -49347 32651 -49301 32655
rect -49505 32574 -49499 32608
rect -49465 32574 -49459 32608
rect -49505 32536 -49459 32574
rect -49505 32502 -49499 32536
rect -49465 32502 -49459 32536
rect -49663 32455 -49617 32459
rect -49505 32361 -49459 32502
rect -49356 32645 -49292 32651
rect -49356 32593 -49350 32645
rect -49298 32593 -49292 32645
rect -49356 32581 -49341 32593
rect -49307 32581 -49292 32593
rect -49356 32529 -49350 32581
rect -49298 32529 -49292 32581
rect -49356 32517 -49341 32529
rect -49307 32517 -49292 32529
rect -49356 32465 -49350 32517
rect -49298 32465 -49292 32517
rect -49356 32459 -49292 32465
rect -49189 32608 -49143 32655
rect -49031 32651 -48985 32655
rect -49189 32574 -49183 32608
rect -49149 32574 -49143 32608
rect -49189 32536 -49143 32574
rect -49189 32502 -49183 32536
rect -49149 32502 -49143 32536
rect -49347 32455 -49301 32459
rect -49189 32361 -49143 32502
rect -49040 32645 -48976 32651
rect -49040 32593 -49034 32645
rect -48982 32593 -48976 32645
rect -49040 32581 -49025 32593
rect -48991 32581 -48976 32593
rect -49040 32529 -49034 32581
rect -48982 32529 -48976 32581
rect -49040 32517 -49025 32529
rect -48991 32517 -48976 32529
rect -49040 32465 -49034 32517
rect -48982 32465 -48976 32517
rect -49040 32459 -48976 32465
rect -48873 32608 -48819 32655
rect -48873 32574 -48867 32608
rect -48833 32574 -48819 32608
rect -48873 32536 -48819 32574
rect -48873 32502 -48867 32536
rect -48833 32502 -48819 32536
rect -49031 32455 -48985 32459
rect -48873 32361 -48819 32502
rect 2131 32593 2396 32657
rect 2768 32593 2774 32965
rect 2886 32951 2900 32985
rect 2934 32951 2940 32985
rect 2886 32912 2940 32951
rect 3043 33298 3107 33304
rect 3043 33246 3049 33298
rect 3101 33246 3107 33298
rect 3043 33239 3058 33246
rect 3092 33239 3107 33246
rect 3043 33234 3107 33239
rect 3043 33182 3049 33234
rect 3101 33182 3107 33234
rect 3043 33170 3058 33182
rect 3092 33170 3107 33182
rect 3043 33118 3049 33170
rect 3101 33118 3107 33170
rect 3043 33106 3058 33118
rect 3092 33106 3107 33118
rect 3043 33054 3049 33106
rect 3101 33054 3107 33106
rect 3043 33042 3058 33054
rect 3092 33042 3107 33054
rect 3043 32990 3049 33042
rect 3101 32990 3107 33042
rect 3043 32985 3107 32990
rect 3043 32978 3058 32985
rect 3092 32978 3107 32985
rect 3043 32926 3049 32978
rect 3101 32926 3107 32978
rect 3043 32920 3107 32926
rect 3210 33273 3256 33406
rect 3368 33304 3414 33312
rect 3210 33239 3216 33273
rect 3250 33239 3256 33273
rect 3210 33201 3256 33239
rect 3210 33167 3216 33201
rect 3250 33167 3256 33201
rect 3210 33129 3256 33167
rect 3210 33095 3216 33129
rect 3250 33095 3256 33129
rect 3210 33057 3256 33095
rect 3210 33023 3216 33057
rect 3250 33023 3256 33057
rect 3210 32985 3256 33023
rect 3210 32951 3216 32985
rect 3250 32951 3256 32985
rect 3052 32912 3098 32920
rect 3210 32912 3256 32951
rect 3359 33298 3423 33304
rect 3359 33246 3365 33298
rect 3417 33246 3423 33298
rect 3359 33239 3374 33246
rect 3408 33239 3423 33246
rect 3359 33234 3423 33239
rect 3359 33182 3365 33234
rect 3417 33182 3423 33234
rect 3359 33170 3374 33182
rect 3408 33170 3423 33182
rect 3359 33118 3365 33170
rect 3417 33118 3423 33170
rect 3359 33106 3374 33118
rect 3408 33106 3423 33118
rect 3359 33054 3365 33106
rect 3417 33054 3423 33106
rect 3359 33042 3374 33054
rect 3408 33042 3423 33054
rect 3359 32990 3365 33042
rect 3417 32990 3423 33042
rect 3359 32985 3423 32990
rect 3359 32978 3374 32985
rect 3408 32978 3423 32985
rect 3359 32926 3365 32978
rect 3417 32926 3423 32978
rect 3359 32920 3423 32926
rect 3526 33273 3572 33406
rect 3684 33304 3730 33312
rect 3526 33239 3532 33273
rect 3566 33239 3572 33273
rect 3526 33201 3572 33239
rect 3526 33167 3532 33201
rect 3566 33167 3572 33201
rect 3526 33129 3572 33167
rect 3526 33095 3532 33129
rect 3566 33095 3572 33129
rect 3526 33057 3572 33095
rect 3526 33023 3532 33057
rect 3566 33023 3572 33057
rect 3526 32985 3572 33023
rect 3526 32951 3532 32985
rect 3566 32951 3572 32985
rect 3368 32912 3414 32920
rect 3526 32912 3572 32951
rect 3675 33298 3739 33304
rect 3675 33246 3681 33298
rect 3733 33246 3739 33298
rect 3675 33239 3690 33246
rect 3724 33239 3739 33246
rect 3675 33234 3739 33239
rect 3675 33182 3681 33234
rect 3733 33182 3739 33234
rect 3675 33170 3690 33182
rect 3724 33170 3739 33182
rect 3675 33118 3681 33170
rect 3733 33118 3739 33170
rect 3675 33106 3690 33118
rect 3724 33106 3739 33118
rect 3675 33054 3681 33106
rect 3733 33054 3739 33106
rect 3675 33042 3690 33054
rect 3724 33042 3739 33054
rect 3675 32990 3681 33042
rect 3733 32990 3739 33042
rect 3675 32985 3739 32990
rect 3675 32978 3690 32985
rect 3724 32978 3739 32985
rect 3675 32926 3681 32978
rect 3733 32926 3739 32978
rect 3675 32920 3739 32926
rect 3842 33273 3888 33406
rect 4000 33304 4046 33312
rect 3842 33239 3848 33273
rect 3882 33239 3888 33273
rect 3842 33201 3888 33239
rect 3842 33167 3848 33201
rect 3882 33167 3888 33201
rect 3842 33129 3888 33167
rect 3842 33095 3848 33129
rect 3882 33095 3888 33129
rect 3842 33057 3888 33095
rect 3842 33023 3848 33057
rect 3882 33023 3888 33057
rect 3842 32985 3888 33023
rect 3842 32951 3848 32985
rect 3882 32951 3888 32985
rect 3684 32912 3730 32920
rect 3842 32912 3888 32951
rect 3991 33298 4055 33304
rect 3991 33246 3997 33298
rect 4049 33246 4055 33298
rect 3991 33239 4006 33246
rect 4040 33239 4055 33246
rect 3991 33234 4055 33239
rect 3991 33182 3997 33234
rect 4049 33182 4055 33234
rect 3991 33170 4006 33182
rect 4040 33170 4055 33182
rect 3991 33118 3997 33170
rect 4049 33118 4055 33170
rect 3991 33106 4006 33118
rect 4040 33106 4055 33118
rect 3991 33054 3997 33106
rect 4049 33054 4055 33106
rect 3991 33042 4006 33054
rect 4040 33042 4055 33054
rect 3991 32990 3997 33042
rect 4049 32990 4055 33042
rect 3991 32985 4055 32990
rect 3991 32978 4006 32985
rect 4040 32978 4055 32985
rect 3991 32926 3997 32978
rect 4049 32926 4055 32978
rect 3991 32920 4055 32926
rect 4158 33273 4204 33406
rect 4316 33304 4362 33312
rect 4158 33239 4164 33273
rect 4198 33239 4204 33273
rect 4158 33201 4204 33239
rect 4158 33167 4164 33201
rect 4198 33167 4204 33201
rect 4158 33129 4204 33167
rect 4158 33095 4164 33129
rect 4198 33095 4204 33129
rect 4158 33057 4204 33095
rect 4158 33023 4164 33057
rect 4198 33023 4204 33057
rect 4158 32985 4204 33023
rect 4158 32951 4164 32985
rect 4198 32951 4204 32985
rect 4000 32912 4046 32920
rect 4158 32912 4204 32951
rect 4307 33298 4371 33304
rect 4307 33246 4313 33298
rect 4365 33246 4371 33298
rect 4307 33239 4322 33246
rect 4356 33239 4371 33246
rect 4307 33234 4371 33239
rect 4307 33182 4313 33234
rect 4365 33182 4371 33234
rect 4307 33170 4322 33182
rect 4356 33170 4371 33182
rect 4307 33118 4313 33170
rect 4365 33118 4371 33170
rect 4307 33106 4322 33118
rect 4356 33106 4371 33118
rect 4307 33054 4313 33106
rect 4365 33054 4371 33106
rect 4307 33042 4322 33054
rect 4356 33042 4371 33054
rect 4307 32990 4313 33042
rect 4365 32990 4371 33042
rect 4307 32985 4371 32990
rect 4307 32978 4322 32985
rect 4356 32978 4371 32985
rect 4307 32926 4313 32978
rect 4365 32926 4371 32978
rect 4307 32920 4371 32926
rect 4474 33273 4528 33406
rect 4474 33239 4480 33273
rect 4514 33239 4528 33273
rect 4474 33201 4528 33239
rect 9994 33236 10000 33864
rect 10308 33236 10314 33864
rect 9994 33210 10314 33236
rect 10994 33864 11314 33890
rect 10994 33236 11000 33864
rect 11308 33236 11314 33864
rect 10994 33210 11314 33236
rect 11994 33864 12314 33890
rect 11994 33236 12000 33864
rect 12308 33236 12314 33864
rect 11994 33210 12314 33236
rect 12994 33864 13314 33890
rect 12994 33236 13000 33864
rect 13308 33236 13314 33864
rect 12994 33210 13314 33236
rect 13994 33864 14314 33890
rect 13994 33236 14000 33864
rect 14308 33236 14314 33864
rect 13994 33210 14314 33236
rect 14994 33864 15314 33890
rect 14994 33236 15000 33864
rect 15308 33236 15314 33864
rect 14994 33210 15314 33236
rect 15994 33864 16314 33890
rect 15994 33236 16000 33864
rect 16308 33236 16314 33864
rect 15994 33210 16314 33236
rect 16994 33864 17314 33890
rect 16994 33236 17000 33864
rect 17308 33236 17314 33864
rect 16994 33210 17314 33236
rect 17994 33864 18314 33890
rect 17994 33236 18000 33864
rect 18308 33236 18314 33864
rect 17994 33210 18314 33236
rect 18994 33864 19314 33890
rect 18994 33236 19000 33864
rect 19308 33236 19314 33864
rect 18994 33210 19314 33236
rect 19994 33864 20314 33890
rect 19994 33236 20000 33864
rect 20308 33236 20314 33864
rect 19994 33210 20314 33236
rect 20994 33864 21314 33890
rect 20994 33236 21000 33864
rect 21308 33236 21314 33864
rect 20994 33210 21314 33236
rect 21994 33864 22314 33890
rect 21994 33236 22000 33864
rect 22308 33236 22314 33864
rect 21994 33210 22314 33236
rect 22994 33864 23314 33890
rect 22994 33236 23000 33864
rect 23308 33236 23314 33864
rect 22994 33210 23314 33236
rect 23994 33864 24314 33890
rect 23994 33236 24000 33864
rect 24308 33236 24314 33864
rect 23994 33210 24314 33236
rect 24994 33864 25314 33890
rect 24994 33236 25000 33864
rect 25308 33236 25314 33864
rect 24994 33210 25314 33236
rect 25994 33864 26314 33890
rect 25994 33236 26000 33864
rect 26308 33236 26314 33864
rect 25994 33210 26314 33236
rect 26994 33864 27314 33890
rect 26994 33236 27000 33864
rect 27308 33236 27314 33864
rect 26994 33210 27314 33236
rect 27994 33864 28314 33890
rect 27994 33236 28000 33864
rect 28308 33236 28314 33864
rect 27994 33210 28314 33236
rect 28994 33864 29314 33890
rect 28994 33236 29000 33864
rect 29308 33236 29314 33864
rect 28994 33210 29314 33236
rect 29994 33864 30314 33890
rect 29994 33236 30000 33864
rect 30308 33236 30314 33864
rect 29994 33210 30314 33236
rect 30994 33864 31314 33890
rect 30994 33236 31000 33864
rect 31308 33236 31314 33864
rect 30994 33210 31314 33236
rect 31994 33864 32314 33890
rect 31994 33236 32000 33864
rect 32308 33236 32314 33864
rect 31994 33210 32314 33236
rect 32994 33864 33314 33890
rect 32994 33236 33000 33864
rect 33308 33236 33314 33864
rect 32994 33210 33314 33236
rect 33994 33864 34314 33890
rect 33994 33236 34000 33864
rect 34308 33236 34314 33864
rect 33994 33210 34314 33236
rect 4474 33167 4480 33201
rect 4514 33167 4528 33201
rect 4474 33129 4528 33167
rect 4474 33095 4480 33129
rect 4514 33095 4528 33129
rect 4474 33057 4528 33095
rect 4474 33023 4480 33057
rect 4514 33023 4528 33057
rect 4474 32985 4528 33023
rect 4474 32951 4480 32985
rect 4514 32951 4528 32985
rect 4316 32912 4362 32920
rect 4474 32912 4528 32951
rect 9654 33204 34654 33210
rect 9654 32896 9660 33204
rect 9968 33172 10340 33204
rect 9968 32928 10032 33172
rect 10276 32928 10340 33172
rect 9968 32896 10340 32928
rect 10968 33172 11340 33204
rect 10968 32928 11032 33172
rect 11276 32928 11340 33172
rect 10968 32896 11340 32928
rect 11968 33172 12340 33204
rect 11968 32928 12032 33172
rect 12276 32928 12340 33172
rect 11968 32896 12340 32928
rect 12968 33172 13340 33204
rect 12968 32928 13032 33172
rect 13276 32928 13340 33172
rect 12968 32896 13340 32928
rect 13968 33172 14340 33204
rect 13968 32928 14032 33172
rect 14276 32928 14340 33172
rect 13968 32896 14340 32928
rect 14968 33172 15340 33204
rect 14968 32928 15032 33172
rect 15276 32928 15340 33172
rect 14968 32896 15340 32928
rect 15968 33172 16340 33204
rect 15968 32928 16032 33172
rect 16276 32928 16340 33172
rect 15968 32896 16340 32928
rect 16968 33172 17340 33204
rect 16968 32928 17032 33172
rect 17276 32928 17340 33172
rect 16968 32896 17340 32928
rect 17968 33172 18340 33204
rect 17968 32928 18032 33172
rect 18276 32928 18340 33172
rect 17968 32896 18340 32928
rect 18968 33172 19340 33204
rect 18968 32928 19032 33172
rect 19276 32928 19340 33172
rect 18968 32896 19340 32928
rect 19968 33172 20340 33204
rect 19968 32928 20032 33172
rect 20276 32928 20340 33172
rect 19968 32896 20340 32928
rect 20968 33172 21340 33204
rect 20968 32928 21032 33172
rect 21276 32928 21340 33172
rect 20968 32896 21340 32928
rect 21968 33172 22340 33204
rect 21968 32928 22032 33172
rect 22276 32928 22340 33172
rect 21968 32896 22340 32928
rect 22968 33172 23340 33204
rect 22968 32928 23032 33172
rect 23276 32928 23340 33172
rect 22968 32896 23340 32928
rect 23968 33172 24340 33204
rect 23968 32928 24032 33172
rect 24276 32928 24340 33172
rect 23968 32896 24340 32928
rect 24968 33172 25340 33204
rect 24968 32928 25032 33172
rect 25276 32928 25340 33172
rect 24968 32896 25340 32928
rect 25968 33172 26340 33204
rect 25968 32928 26032 33172
rect 26276 32928 26340 33172
rect 25968 32896 26340 32928
rect 26968 33172 27340 33204
rect 26968 32928 27032 33172
rect 27276 32928 27340 33172
rect 26968 32896 27340 32928
rect 27968 33172 28340 33204
rect 27968 32928 28032 33172
rect 28276 32928 28340 33172
rect 27968 32896 28340 32928
rect 28968 33172 29340 33204
rect 28968 32928 29032 33172
rect 29276 32928 29340 33172
rect 28968 32896 29340 32928
rect 29968 33172 30340 33204
rect 29968 32928 30032 33172
rect 30276 32928 30340 33172
rect 29968 32896 30340 32928
rect 30968 33172 31340 33204
rect 30968 32928 31032 33172
rect 31276 32928 31340 33172
rect 30968 32896 31340 32928
rect 31968 33172 32340 33204
rect 31968 32928 32032 33172
rect 32276 32928 32340 33172
rect 31968 32896 32340 32928
rect 32968 33172 33340 33204
rect 32968 32928 33032 33172
rect 33276 32928 33340 33172
rect 32968 32896 33340 32928
rect 33968 33172 34340 33204
rect 33968 32928 34032 33172
rect 34276 32928 34340 33172
rect 33968 32896 34340 32928
rect 34648 32896 34654 33204
rect 9654 32890 34654 32896
rect 2950 32865 3042 32871
rect 2950 32831 2979 32865
rect 3013 32831 3042 32865
rect 2950 32825 3042 32831
rect 3108 32865 3200 32871
rect 3108 32831 3137 32865
rect 3171 32831 3200 32865
rect 3108 32825 3200 32831
rect 3266 32865 3358 32871
rect 3266 32831 3295 32865
rect 3329 32831 3358 32865
rect 3266 32825 3358 32831
rect 3424 32865 3516 32871
rect 3424 32831 3453 32865
rect 3487 32831 3516 32865
rect 3424 32825 3516 32831
rect 3582 32865 3674 32871
rect 3582 32831 3611 32865
rect 3645 32831 3674 32865
rect 3582 32825 3674 32831
rect 3740 32865 3832 32871
rect 3740 32831 3769 32865
rect 3803 32831 3832 32865
rect 3740 32825 3832 32831
rect 3898 32865 3990 32871
rect 3898 32831 3927 32865
rect 3961 32831 3990 32865
rect 3898 32825 3990 32831
rect 4056 32865 4148 32871
rect 4056 32831 4085 32865
rect 4119 32831 4148 32865
rect 4056 32825 4148 32831
rect 4214 32865 4306 32871
rect 4214 32831 4243 32865
rect 4277 32831 4306 32865
rect 4214 32825 4306 32831
rect 4372 32865 4464 32871
rect 4372 32831 4401 32865
rect 4435 32831 4464 32865
rect 4372 32825 4464 32831
rect 9994 32864 10314 32890
rect 2950 32727 3042 32733
rect 2950 32693 2979 32727
rect 3013 32693 3042 32727
rect 2950 32687 3042 32693
rect 3108 32727 3200 32733
rect 3108 32693 3137 32727
rect 3171 32693 3200 32727
rect 3108 32687 3200 32693
rect 3266 32727 3358 32733
rect 3266 32693 3295 32727
rect 3329 32693 3358 32727
rect 3266 32687 3358 32693
rect 3424 32727 3516 32733
rect 3424 32693 3453 32727
rect 3487 32693 3516 32727
rect 3424 32687 3516 32693
rect 3582 32727 3674 32733
rect 3582 32693 3611 32727
rect 3645 32693 3674 32727
rect 3582 32687 3674 32693
rect 3740 32727 3832 32733
rect 3740 32693 3769 32727
rect 3803 32693 3832 32727
rect 3740 32687 3832 32693
rect 3898 32727 3990 32733
rect 3898 32693 3927 32727
rect 3961 32693 3990 32727
rect 3898 32687 3990 32693
rect 4056 32727 4148 32733
rect 4056 32693 4085 32727
rect 4119 32693 4148 32727
rect 4056 32687 4148 32693
rect 4214 32727 4306 32733
rect 4214 32693 4243 32727
rect 4277 32693 4306 32727
rect 4214 32687 4306 32693
rect 4372 32727 4464 32733
rect 4372 32693 4401 32727
rect 4435 32693 4464 32727
rect 4372 32687 4464 32693
rect 2131 32567 2774 32593
rect 2886 32608 2940 32655
rect 3052 32651 3098 32655
rect 2886 32574 2900 32608
rect 2934 32574 2940 32608
rect 2131 32539 2209 32567
rect 2131 32505 2153 32539
rect 2187 32505 2209 32539
rect 2131 32477 2209 32505
rect 2886 32536 2940 32574
rect 2886 32502 2900 32536
rect 2934 32502 2940 32536
rect -50461 32349 -48819 32361
rect -50461 32243 -50449 32349
rect -48831 32243 -48819 32349
rect -50461 32231 -48819 32243
rect 1967 32359 2313 32371
rect 1967 32253 1979 32359
rect 2301 32253 2313 32359
rect 1967 32231 2313 32253
rect 2886 32361 2940 32502
rect 3043 32645 3107 32651
rect 3043 32593 3049 32645
rect 3101 32593 3107 32645
rect 3043 32581 3058 32593
rect 3092 32581 3107 32593
rect 3043 32529 3049 32581
rect 3101 32529 3107 32581
rect 3043 32517 3058 32529
rect 3092 32517 3107 32529
rect 3043 32465 3049 32517
rect 3101 32465 3107 32517
rect 3043 32459 3107 32465
rect 3210 32608 3256 32655
rect 3368 32651 3414 32655
rect 3210 32574 3216 32608
rect 3250 32574 3256 32608
rect 3210 32536 3256 32574
rect 3210 32502 3216 32536
rect 3250 32502 3256 32536
rect 3052 32455 3098 32459
rect 3210 32361 3256 32502
rect 3359 32645 3423 32651
rect 3359 32593 3365 32645
rect 3417 32593 3423 32645
rect 3359 32581 3374 32593
rect 3408 32581 3423 32593
rect 3359 32529 3365 32581
rect 3417 32529 3423 32581
rect 3359 32517 3374 32529
rect 3408 32517 3423 32529
rect 3359 32465 3365 32517
rect 3417 32465 3423 32517
rect 3359 32459 3423 32465
rect 3526 32608 3572 32655
rect 3684 32651 3730 32655
rect 3526 32574 3532 32608
rect 3566 32574 3572 32608
rect 3526 32536 3572 32574
rect 3526 32502 3532 32536
rect 3566 32502 3572 32536
rect 3368 32455 3414 32459
rect 3526 32361 3572 32502
rect 3675 32645 3739 32651
rect 3675 32593 3681 32645
rect 3733 32593 3739 32645
rect 3675 32581 3690 32593
rect 3724 32581 3739 32593
rect 3675 32529 3681 32581
rect 3733 32529 3739 32581
rect 3675 32517 3690 32529
rect 3724 32517 3739 32529
rect 3675 32465 3681 32517
rect 3733 32465 3739 32517
rect 3675 32459 3739 32465
rect 3842 32608 3888 32655
rect 4000 32651 4046 32655
rect 3842 32574 3848 32608
rect 3882 32574 3888 32608
rect 3842 32536 3888 32574
rect 3842 32502 3848 32536
rect 3882 32502 3888 32536
rect 3684 32455 3730 32459
rect 3842 32361 3888 32502
rect 3991 32645 4055 32651
rect 3991 32593 3997 32645
rect 4049 32593 4055 32645
rect 3991 32581 4006 32593
rect 4040 32581 4055 32593
rect 3991 32529 3997 32581
rect 4049 32529 4055 32581
rect 3991 32517 4006 32529
rect 4040 32517 4055 32529
rect 3991 32465 3997 32517
rect 4049 32465 4055 32517
rect 3991 32459 4055 32465
rect 4158 32608 4204 32655
rect 4316 32651 4362 32655
rect 4158 32574 4164 32608
rect 4198 32574 4204 32608
rect 4158 32536 4204 32574
rect 4158 32502 4164 32536
rect 4198 32502 4204 32536
rect 4000 32455 4046 32459
rect 4158 32361 4204 32502
rect 4307 32645 4371 32651
rect 4307 32593 4313 32645
rect 4365 32593 4371 32645
rect 4307 32581 4322 32593
rect 4356 32581 4371 32593
rect 4307 32529 4313 32581
rect 4365 32529 4371 32581
rect 4307 32517 4322 32529
rect 4356 32517 4371 32529
rect 4307 32465 4313 32517
rect 4365 32465 4371 32517
rect 4307 32459 4371 32465
rect 4474 32608 4528 32655
rect 4474 32574 4480 32608
rect 4514 32574 4528 32608
rect 4474 32536 4528 32574
rect 4474 32502 4480 32536
rect 4514 32502 4528 32536
rect 4316 32455 4362 32459
rect 4474 32361 4528 32502
rect 2886 32349 4528 32361
rect 2886 32243 2898 32349
rect 4516 32243 4528 32349
rect 2886 32231 4528 32243
rect 9994 32236 10000 32864
rect 10308 32236 10314 32864
rect -50461 32210 9654 32231
rect 9994 32210 10314 32236
rect 10994 32864 11314 32890
rect 10994 32236 11000 32864
rect 11308 32236 11314 32864
rect 10994 32210 11314 32236
rect 11994 32864 12314 32890
rect 11994 32236 12000 32864
rect 12308 32236 12314 32864
rect 11994 32210 12314 32236
rect 12994 32864 13314 32890
rect 12994 32236 13000 32864
rect 13308 32236 13314 32864
rect 12994 32210 13314 32236
rect 13994 32864 14314 32890
rect 13994 32236 14000 32864
rect 14308 32236 14314 32864
rect 13994 32210 14314 32236
rect 14994 32864 15314 32890
rect 14994 32236 15000 32864
rect 15308 32236 15314 32864
rect 14994 32210 15314 32236
rect 15994 32864 16314 32890
rect 15994 32236 16000 32864
rect 16308 32236 16314 32864
rect 15994 32210 16314 32236
rect 16994 32864 17314 32890
rect 16994 32236 17000 32864
rect 17308 32236 17314 32864
rect 16994 32210 17314 32236
rect 17994 32864 18314 32890
rect 17994 32236 18000 32864
rect 18308 32236 18314 32864
rect 17994 32210 18314 32236
rect 18994 32864 19314 32890
rect 18994 32236 19000 32864
rect 19308 32236 19314 32864
rect 18994 32210 19314 32236
rect 19994 32864 20314 32890
rect 19994 32236 20000 32864
rect 20308 32236 20314 32864
rect 19994 32210 20314 32236
rect 20994 32864 21314 32890
rect 20994 32236 21000 32864
rect 21308 32236 21314 32864
rect 20994 32210 21314 32236
rect 21994 32864 22314 32890
rect 21994 32236 22000 32864
rect 22308 32236 22314 32864
rect 21994 32210 22314 32236
rect 22994 32864 23314 32890
rect 22994 32236 23000 32864
rect 23308 32236 23314 32864
rect 22994 32210 23314 32236
rect 23994 32864 24314 32890
rect 23994 32236 24000 32864
rect 24308 32236 24314 32864
rect 23994 32210 24314 32236
rect 24994 32864 25314 32890
rect 24994 32236 25000 32864
rect 25308 32236 25314 32864
rect 24994 32210 25314 32236
rect 25994 32864 26314 32890
rect 25994 32236 26000 32864
rect 26308 32236 26314 32864
rect 25994 32210 26314 32236
rect 26994 32864 27314 32890
rect 26994 32236 27000 32864
rect 27308 32236 27314 32864
rect 26994 32210 27314 32236
rect 27994 32864 28314 32890
rect 27994 32236 28000 32864
rect 28308 32236 28314 32864
rect 27994 32210 28314 32236
rect 28994 32864 29314 32890
rect 28994 32236 29000 32864
rect 29308 32236 29314 32864
rect 28994 32210 29314 32236
rect 29994 32864 30314 32890
rect 29994 32236 30000 32864
rect 30308 32236 30314 32864
rect 29994 32210 30314 32236
rect 30994 32864 31314 32890
rect 30994 32236 31000 32864
rect 31308 32236 31314 32864
rect 30994 32210 31314 32236
rect 31994 32864 32314 32890
rect 31994 32236 32000 32864
rect 32308 32236 32314 32864
rect 31994 32210 32314 32236
rect 32994 32864 33314 32890
rect 32994 32236 33000 32864
rect 33308 32236 33314 32864
rect 32994 32210 33314 32236
rect 33994 32864 34314 32890
rect 33994 32236 34000 32864
rect 34308 32236 34314 32864
rect 33994 32210 34314 32236
rect -50461 32204 34654 32210
rect -50461 32161 9660 32204
rect -50797 32001 -50769 32035
rect -50735 32001 -50707 32035
rect -50797 31979 -50707 32001
rect -50601 32149 9660 32161
rect -74825 31890 -58825 31896
rect -74485 31864 -74165 31890
rect -74485 31236 -74479 31864
rect -74171 31236 -74165 31864
rect -74485 31210 -74165 31236
rect -73485 31864 -73165 31890
rect -73485 31236 -73479 31864
rect -73171 31236 -73165 31864
rect -73485 31210 -73165 31236
rect -72485 31864 -72165 31890
rect -72485 31236 -72479 31864
rect -72171 31236 -72165 31864
rect -72485 31210 -72165 31236
rect -71485 31864 -71165 31890
rect -71485 31236 -71479 31864
rect -71171 31236 -71165 31864
rect -71485 31210 -71165 31236
rect -70485 31864 -70165 31890
rect -70485 31236 -70479 31864
rect -70171 31236 -70165 31864
rect -70485 31210 -70165 31236
rect -69485 31864 -69165 31890
rect -69485 31236 -69479 31864
rect -69171 31236 -69165 31864
rect -69485 31210 -69165 31236
rect -68485 31864 -68165 31890
rect -68485 31236 -68479 31864
rect -68171 31236 -68165 31864
rect -68485 31210 -68165 31236
rect -67485 31864 -67165 31890
rect -67485 31236 -67479 31864
rect -67171 31236 -67165 31864
rect -67485 31210 -67165 31236
rect -66485 31864 -66165 31890
rect -66485 31236 -66479 31864
rect -66171 31236 -66165 31864
rect -66485 31210 -66165 31236
rect -65485 31864 -65165 31890
rect -65485 31236 -65479 31864
rect -65171 31236 -65165 31864
rect -65485 31210 -65165 31236
rect -64485 31864 -64165 31890
rect -64485 31236 -64479 31864
rect -64171 31236 -64165 31864
rect -64485 31210 -64165 31236
rect -63485 31864 -63165 31890
rect -63485 31236 -63479 31864
rect -63171 31236 -63165 31864
rect -63485 31210 -63165 31236
rect -62485 31864 -62165 31890
rect -62485 31236 -62479 31864
rect -62171 31236 -62165 31864
rect -62485 31210 -62165 31236
rect -61485 31864 -61165 31890
rect -61485 31236 -61479 31864
rect -61171 31236 -61165 31864
rect -61485 31210 -61165 31236
rect -60485 31864 -60165 31890
rect -60485 31236 -60479 31864
rect -60171 31236 -60165 31864
rect -60485 31210 -60165 31236
rect -59485 31864 -59165 31890
rect -59485 31236 -59479 31864
rect -59171 31236 -59165 31864
rect -50601 31827 -50589 32149
rect -50483 31896 9660 32149
rect 9968 32172 10340 32204
rect 9968 31928 10032 32172
rect 10276 31928 10340 32172
rect 9968 31896 10340 31928
rect 10968 32172 11340 32204
rect 10968 31928 11032 32172
rect 11276 31928 11340 32172
rect 10968 31896 11340 31928
rect 11968 32172 12340 32204
rect 11968 31928 12032 32172
rect 12276 31928 12340 32172
rect 11968 31896 12340 31928
rect 12968 32172 13340 32204
rect 12968 31928 13032 32172
rect 13276 31928 13340 32172
rect 12968 31896 13340 31928
rect 13968 32172 14340 32204
rect 13968 31928 14032 32172
rect 14276 31928 14340 32172
rect 13968 31896 14340 31928
rect 14968 32172 15340 32204
rect 14968 31928 15032 32172
rect 15276 31928 15340 32172
rect 14968 31896 15340 31928
rect 15968 32172 16340 32204
rect 15968 31928 16032 32172
rect 16276 31928 16340 32172
rect 15968 31896 16340 31928
rect 16968 32172 17340 32204
rect 16968 31928 17032 32172
rect 17276 31928 17340 32172
rect 16968 31896 17340 31928
rect 17968 32172 18340 32204
rect 17968 31928 18032 32172
rect 18276 31928 18340 32172
rect 17968 31896 18340 31928
rect 18968 32172 19340 32204
rect 18968 31928 19032 32172
rect 19276 31928 19340 32172
rect 18968 31896 19340 31928
rect 19968 32172 20340 32204
rect 19968 31928 20032 32172
rect 20276 31928 20340 32172
rect 19968 31896 20340 31928
rect 20968 32172 21340 32204
rect 20968 31928 21032 32172
rect 21276 31928 21340 32172
rect 20968 31896 21340 31928
rect 21968 32172 22340 32204
rect 21968 31928 22032 32172
rect 22276 31928 22340 32172
rect 21968 31896 22340 31928
rect 22968 32172 23340 32204
rect 22968 31928 23032 32172
rect 23276 31928 23340 32172
rect 22968 31896 23340 31928
rect 23968 32172 24340 32204
rect 23968 31928 24032 32172
rect 24276 31928 24340 32172
rect 23968 31896 24340 31928
rect 24968 32172 25340 32204
rect 24968 31928 25032 32172
rect 25276 31928 25340 32172
rect 24968 31896 25340 31928
rect 25968 32172 26340 32204
rect 25968 31928 26032 32172
rect 26276 31928 26340 32172
rect 25968 31896 26340 31928
rect 26968 32172 27340 32204
rect 26968 31928 27032 32172
rect 27276 31928 27340 32172
rect 26968 31896 27340 31928
rect 27968 32172 28340 32204
rect 27968 31928 28032 32172
rect 28276 31928 28340 32172
rect 27968 31896 28340 31928
rect 28968 32172 29340 32204
rect 28968 31928 29032 32172
rect 29276 31928 29340 32172
rect 28968 31896 29340 31928
rect 29968 32172 30340 32204
rect 29968 31928 30032 32172
rect 30276 31928 30340 32172
rect 29968 31896 30340 31928
rect 30968 32172 31340 32204
rect 30968 31928 31032 32172
rect 31276 31928 31340 32172
rect 30968 31896 31340 31928
rect 31968 32172 32340 32204
rect 31968 31928 32032 32172
rect 32276 31928 32340 32172
rect 31968 31896 32340 31928
rect 32968 32172 33340 32204
rect 32968 31928 33032 32172
rect 33276 31928 33340 32172
rect 32968 31896 33340 31928
rect 33968 32172 34340 32204
rect 33968 31928 34032 32172
rect 34276 31928 34340 32172
rect 33968 31896 34340 31928
rect 34648 31896 34654 32204
rect -50483 31890 34654 31896
rect -50483 31827 9654 31890
rect -50601 31815 9654 31827
rect -59485 31210 -59165 31236
rect -50461 31210 9654 31815
rect 9994 31864 10314 31890
rect 9994 31236 10000 31864
rect 10308 31236 10314 31864
rect 9994 31210 10314 31236
rect 10994 31864 11314 31890
rect 10994 31236 11000 31864
rect 11308 31236 11314 31864
rect 10994 31210 11314 31236
rect 11994 31864 12314 31890
rect 11994 31236 12000 31864
rect 12308 31236 12314 31864
rect 11994 31210 12314 31236
rect 12994 31864 13314 31890
rect 12994 31236 13000 31864
rect 13308 31236 13314 31864
rect 12994 31210 13314 31236
rect 13994 31864 14314 31890
rect 13994 31236 14000 31864
rect 14308 31236 14314 31864
rect 13994 31210 14314 31236
rect 14994 31864 15314 31890
rect 14994 31236 15000 31864
rect 15308 31236 15314 31864
rect 14994 31210 15314 31236
rect 15994 31864 16314 31890
rect 15994 31236 16000 31864
rect 16308 31236 16314 31864
rect 15994 31210 16314 31236
rect 16994 31864 17314 31890
rect 16994 31236 17000 31864
rect 17308 31236 17314 31864
rect 16994 31210 17314 31236
rect 17994 31864 18314 31890
rect 17994 31236 18000 31864
rect 18308 31236 18314 31864
rect 17994 31210 18314 31236
rect 18994 31864 19314 31890
rect 18994 31236 19000 31864
rect 19308 31236 19314 31864
rect 18994 31210 19314 31236
rect 19994 31864 20314 31890
rect 19994 31236 20000 31864
rect 20308 31236 20314 31864
rect 19994 31210 20314 31236
rect 20994 31864 21314 31890
rect 20994 31236 21000 31864
rect 21308 31236 21314 31864
rect 20994 31210 21314 31236
rect 21994 31864 22314 31890
rect 21994 31236 22000 31864
rect 22308 31236 22314 31864
rect 21994 31210 22314 31236
rect 22994 31864 23314 31890
rect 22994 31236 23000 31864
rect 23308 31236 23314 31864
rect 22994 31210 23314 31236
rect 23994 31864 24314 31890
rect 23994 31236 24000 31864
rect 24308 31236 24314 31864
rect 23994 31210 24314 31236
rect 24994 31864 25314 31890
rect 24994 31236 25000 31864
rect 25308 31236 25314 31864
rect 24994 31210 25314 31236
rect 25994 31864 26314 31890
rect 25994 31236 26000 31864
rect 26308 31236 26314 31864
rect 25994 31210 26314 31236
rect 26994 31864 27314 31890
rect 26994 31236 27000 31864
rect 27308 31236 27314 31864
rect 26994 31210 27314 31236
rect 27994 31864 28314 31890
rect 27994 31236 28000 31864
rect 28308 31236 28314 31864
rect 27994 31210 28314 31236
rect 28994 31864 29314 31890
rect 28994 31236 29000 31864
rect 29308 31236 29314 31864
rect 28994 31210 29314 31236
rect 29994 31864 30314 31890
rect 29994 31236 30000 31864
rect 30308 31236 30314 31864
rect 29994 31210 30314 31236
rect 30994 31864 31314 31890
rect 30994 31236 31000 31864
rect 31308 31236 31314 31864
rect 30994 31210 31314 31236
rect 31994 31864 32314 31890
rect 31994 31236 32000 31864
rect 32308 31236 32314 31864
rect 31994 31210 32314 31236
rect 32994 31864 33314 31890
rect 32994 31236 33000 31864
rect 33308 31236 33314 31864
rect 32994 31210 33314 31236
rect 33994 31864 34314 31890
rect 33994 31236 34000 31864
rect 34308 31236 34314 31864
rect 33994 31210 34314 31236
rect -74825 31204 -58825 31210
rect -74825 30896 -74819 31204
rect -74511 31172 -74139 31204
rect -74511 30928 -74447 31172
rect -74203 30928 -74139 31172
rect -74511 30896 -74139 30928
rect -73511 31172 -73139 31204
rect -73511 30928 -73447 31172
rect -73203 30928 -73139 31172
rect -73511 30896 -73139 30928
rect -72511 31172 -72139 31204
rect -72511 30928 -72447 31172
rect -72203 30928 -72139 31172
rect -72511 30896 -72139 30928
rect -71511 31172 -71139 31204
rect -71511 30928 -71447 31172
rect -71203 30928 -71139 31172
rect -71511 30896 -71139 30928
rect -70511 31172 -70139 31204
rect -70511 30928 -70447 31172
rect -70203 30928 -70139 31172
rect -70511 30896 -70139 30928
rect -69511 31172 -69139 31204
rect -69511 30928 -69447 31172
rect -69203 30928 -69139 31172
rect -69511 30896 -69139 30928
rect -68511 31172 -68139 31204
rect -68511 30928 -68447 31172
rect -68203 30928 -68139 31172
rect -68511 30896 -68139 30928
rect -67511 31172 -67139 31204
rect -67511 30928 -67447 31172
rect -67203 30928 -67139 31172
rect -67511 30896 -67139 30928
rect -66511 31172 -66139 31204
rect -66511 30928 -66447 31172
rect -66203 30928 -66139 31172
rect -66511 30896 -66139 30928
rect -65511 31172 -65139 31204
rect -65511 30928 -65447 31172
rect -65203 30928 -65139 31172
rect -65511 30896 -65139 30928
rect -64511 31172 -64139 31204
rect -64511 30928 -64447 31172
rect -64203 30928 -64139 31172
rect -64511 30896 -64139 30928
rect -63511 31172 -63139 31204
rect -63511 30928 -63447 31172
rect -63203 30928 -63139 31172
rect -63511 30896 -63139 30928
rect -62511 31172 -62139 31204
rect -62511 30928 -62447 31172
rect -62203 30928 -62139 31172
rect -62511 30896 -62139 30928
rect -61511 31172 -61139 31204
rect -61511 30928 -61447 31172
rect -61203 30928 -61139 31172
rect -61511 30896 -61139 30928
rect -60511 31172 -60139 31204
rect -60511 30928 -60447 31172
rect -60203 30928 -60139 31172
rect -60511 30896 -60139 30928
rect -59511 31172 -59139 31204
rect -59511 30928 -59447 31172
rect -59203 30928 -59139 31172
rect -59511 30896 -59139 30928
rect -58831 30896 -58825 31204
rect -74825 30890 -58825 30896
rect -50461 31204 34654 31210
rect -50461 30896 9660 31204
rect 9968 31172 10340 31204
rect 9968 30928 10032 31172
rect 10276 30928 10340 31172
rect 9968 30896 10340 30928
rect 10968 31172 11340 31204
rect 10968 30928 11032 31172
rect 11276 30928 11340 31172
rect 10968 30896 11340 30928
rect 11968 31172 12340 31204
rect 11968 30928 12032 31172
rect 12276 30928 12340 31172
rect 11968 30896 12340 30928
rect 12968 31172 13340 31204
rect 12968 30928 13032 31172
rect 13276 30928 13340 31172
rect 12968 30896 13340 30928
rect 13968 31172 14340 31204
rect 13968 30928 14032 31172
rect 14276 30928 14340 31172
rect 13968 30896 14340 30928
rect 14968 31172 15340 31204
rect 14968 30928 15032 31172
rect 15276 30928 15340 31172
rect 14968 30896 15340 30928
rect 15968 31172 16340 31204
rect 15968 30928 16032 31172
rect 16276 30928 16340 31172
rect 15968 30896 16340 30928
rect 16968 31172 17340 31204
rect 16968 30928 17032 31172
rect 17276 30928 17340 31172
rect 16968 30896 17340 30928
rect 17968 31172 18340 31204
rect 17968 30928 18032 31172
rect 18276 30928 18340 31172
rect 17968 30896 18340 30928
rect 18968 31172 19340 31204
rect 18968 30928 19032 31172
rect 19276 30928 19340 31172
rect 18968 30896 19340 30928
rect 19968 31172 20340 31204
rect 19968 30928 20032 31172
rect 20276 30928 20340 31172
rect 19968 30896 20340 30928
rect 20968 31172 21340 31204
rect 20968 30928 21032 31172
rect 21276 30928 21340 31172
rect 20968 30896 21340 30928
rect 21968 31172 22340 31204
rect 21968 30928 22032 31172
rect 22276 30928 22340 31172
rect 21968 30896 22340 30928
rect 22968 31172 23340 31204
rect 22968 30928 23032 31172
rect 23276 30928 23340 31172
rect 22968 30896 23340 30928
rect 23968 31172 24340 31204
rect 23968 30928 24032 31172
rect 24276 30928 24340 31172
rect 23968 30896 24340 30928
rect 24968 31172 25340 31204
rect 24968 30928 25032 31172
rect 25276 30928 25340 31172
rect 24968 30896 25340 30928
rect 25968 31172 26340 31204
rect 25968 30928 26032 31172
rect 26276 30928 26340 31172
rect 25968 30896 26340 30928
rect 26968 31172 27340 31204
rect 26968 30928 27032 31172
rect 27276 30928 27340 31172
rect 26968 30896 27340 30928
rect 27968 31172 28340 31204
rect 27968 30928 28032 31172
rect 28276 30928 28340 31172
rect 27968 30896 28340 30928
rect 28968 31172 29340 31204
rect 28968 30928 29032 31172
rect 29276 30928 29340 31172
rect 28968 30896 29340 30928
rect 29968 31172 30340 31204
rect 29968 30928 30032 31172
rect 30276 30928 30340 31172
rect 29968 30896 30340 30928
rect 30968 31172 31340 31204
rect 30968 30928 31032 31172
rect 31276 30928 31340 31172
rect 30968 30896 31340 30928
rect 31968 31172 32340 31204
rect 31968 30928 32032 31172
rect 32276 30928 32340 31172
rect 31968 30896 32340 30928
rect 32968 31172 33340 31204
rect 32968 30928 33032 31172
rect 33276 30928 33340 31172
rect 32968 30896 33340 30928
rect 33968 31172 34340 31204
rect 33968 30928 34032 31172
rect 34276 30928 34340 31172
rect 33968 30896 34340 30928
rect 34648 30896 34654 31204
rect -50461 30890 34654 30896
rect -74485 30864 -74165 30890
rect -74485 30236 -74479 30864
rect -74171 30236 -74165 30864
rect -74485 30210 -74165 30236
rect -73485 30864 -73165 30890
rect -73485 30236 -73479 30864
rect -73171 30236 -73165 30864
rect -73485 30210 -73165 30236
rect -72485 30864 -72165 30890
rect -72485 30236 -72479 30864
rect -72171 30236 -72165 30864
rect -72485 30210 -72165 30236
rect -71485 30864 -71165 30890
rect -71485 30236 -71479 30864
rect -71171 30236 -71165 30864
rect -71485 30210 -71165 30236
rect -70485 30864 -70165 30890
rect -70485 30236 -70479 30864
rect -70171 30236 -70165 30864
rect -70485 30210 -70165 30236
rect -69485 30864 -69165 30890
rect -69485 30236 -69479 30864
rect -69171 30236 -69165 30864
rect -69485 30210 -69165 30236
rect -68485 30864 -68165 30890
rect -68485 30236 -68479 30864
rect -68171 30236 -68165 30864
rect -68485 30210 -68165 30236
rect -67485 30864 -67165 30890
rect -67485 30236 -67479 30864
rect -67171 30236 -67165 30864
rect -67485 30210 -67165 30236
rect -66485 30864 -66165 30890
rect -66485 30236 -66479 30864
rect -66171 30236 -66165 30864
rect -66485 30210 -66165 30236
rect -65485 30864 -65165 30890
rect -65485 30236 -65479 30864
rect -65171 30236 -65165 30864
rect -65485 30210 -65165 30236
rect -64485 30864 -64165 30890
rect -64485 30236 -64479 30864
rect -64171 30236 -64165 30864
rect -64485 30210 -64165 30236
rect -63485 30864 -63165 30890
rect -63485 30236 -63479 30864
rect -63171 30236 -63165 30864
rect -63485 30210 -63165 30236
rect -62485 30864 -62165 30890
rect -62485 30236 -62479 30864
rect -62171 30236 -62165 30864
rect -62485 30210 -62165 30236
rect -61485 30864 -61165 30890
rect -61485 30236 -61479 30864
rect -61171 30236 -61165 30864
rect -61485 30210 -61165 30236
rect -60485 30864 -60165 30890
rect -60485 30236 -60479 30864
rect -60171 30236 -60165 30864
rect -60485 30210 -60165 30236
rect -59485 30864 -59165 30890
rect -59485 30236 -59479 30864
rect -59171 30236 -59165 30864
rect -59485 30210 -59165 30236
rect -50461 30210 9654 30890
rect 9994 30864 10314 30890
rect 9994 30236 10000 30864
rect 10308 30236 10314 30864
rect 9994 30210 10314 30236
rect 10994 30864 11314 30890
rect 10994 30236 11000 30864
rect 11308 30236 11314 30864
rect 10994 30210 11314 30236
rect 11994 30864 12314 30890
rect 11994 30236 12000 30864
rect 12308 30236 12314 30864
rect 11994 30210 12314 30236
rect 12994 30864 13314 30890
rect 12994 30236 13000 30864
rect 13308 30236 13314 30864
rect 12994 30210 13314 30236
rect 13994 30864 14314 30890
rect 13994 30236 14000 30864
rect 14308 30236 14314 30864
rect 13994 30210 14314 30236
rect 14994 30864 15314 30890
rect 14994 30236 15000 30864
rect 15308 30236 15314 30864
rect 14994 30210 15314 30236
rect 15994 30864 16314 30890
rect 15994 30236 16000 30864
rect 16308 30236 16314 30864
rect 15994 30210 16314 30236
rect 16994 30864 17314 30890
rect 16994 30236 17000 30864
rect 17308 30236 17314 30864
rect 16994 30210 17314 30236
rect 17994 30864 18314 30890
rect 17994 30236 18000 30864
rect 18308 30236 18314 30864
rect 17994 30210 18314 30236
rect 18994 30864 19314 30890
rect 18994 30236 19000 30864
rect 19308 30236 19314 30864
rect 18994 30210 19314 30236
rect 19994 30864 20314 30890
rect 19994 30236 20000 30864
rect 20308 30236 20314 30864
rect 19994 30210 20314 30236
rect 20994 30864 21314 30890
rect 20994 30236 21000 30864
rect 21308 30236 21314 30864
rect 20994 30210 21314 30236
rect 21994 30864 22314 30890
rect 21994 30236 22000 30864
rect 22308 30236 22314 30864
rect 21994 30210 22314 30236
rect 22994 30864 23314 30890
rect 22994 30236 23000 30864
rect 23308 30236 23314 30864
rect 22994 30210 23314 30236
rect 23994 30864 24314 30890
rect 23994 30236 24000 30864
rect 24308 30236 24314 30864
rect 23994 30210 24314 30236
rect 24994 30864 25314 30890
rect 24994 30236 25000 30864
rect 25308 30236 25314 30864
rect 24994 30210 25314 30236
rect 25994 30864 26314 30890
rect 25994 30236 26000 30864
rect 26308 30236 26314 30864
rect 25994 30210 26314 30236
rect 26994 30864 27314 30890
rect 26994 30236 27000 30864
rect 27308 30236 27314 30864
rect 26994 30210 27314 30236
rect 27994 30864 28314 30890
rect 27994 30236 28000 30864
rect 28308 30236 28314 30864
rect 27994 30210 28314 30236
rect 28994 30864 29314 30890
rect 28994 30236 29000 30864
rect 29308 30236 29314 30864
rect 28994 30210 29314 30236
rect 29994 30864 30314 30890
rect 29994 30236 30000 30864
rect 30308 30236 30314 30864
rect 29994 30210 30314 30236
rect 30994 30864 31314 30890
rect 30994 30236 31000 30864
rect 31308 30236 31314 30864
rect 30994 30210 31314 30236
rect 31994 30864 32314 30890
rect 31994 30236 32000 30864
rect 32308 30236 32314 30864
rect 31994 30210 32314 30236
rect 32994 30864 33314 30890
rect 32994 30236 33000 30864
rect 33308 30236 33314 30864
rect 32994 30210 33314 30236
rect 33994 30864 34314 30890
rect 33994 30236 34000 30864
rect 34308 30236 34314 30864
rect 33994 30210 34314 30236
rect -74825 30204 -58825 30210
rect -74825 29896 -74819 30204
rect -74511 30172 -74139 30204
rect -74511 29928 -74447 30172
rect -74203 29928 -74139 30172
rect -74511 29896 -74139 29928
rect -73511 30172 -73139 30204
rect -73511 29928 -73447 30172
rect -73203 29928 -73139 30172
rect -73511 29896 -73139 29928
rect -72511 30172 -72139 30204
rect -72511 29928 -72447 30172
rect -72203 29928 -72139 30172
rect -72511 29896 -72139 29928
rect -71511 30172 -71139 30204
rect -71511 29928 -71447 30172
rect -71203 29928 -71139 30172
rect -71511 29896 -71139 29928
rect -70511 30172 -70139 30204
rect -70511 29928 -70447 30172
rect -70203 29928 -70139 30172
rect -70511 29896 -70139 29928
rect -69511 30172 -69139 30204
rect -69511 29928 -69447 30172
rect -69203 29928 -69139 30172
rect -69511 29896 -69139 29928
rect -68511 30172 -68139 30204
rect -68511 29928 -68447 30172
rect -68203 29928 -68139 30172
rect -68511 29896 -68139 29928
rect -67511 30172 -67139 30204
rect -67511 29928 -67447 30172
rect -67203 29928 -67139 30172
rect -67511 29896 -67139 29928
rect -66511 30172 -66139 30204
rect -66511 29928 -66447 30172
rect -66203 29928 -66139 30172
rect -66511 29896 -66139 29928
rect -65511 30172 -65139 30204
rect -65511 29928 -65447 30172
rect -65203 29928 -65139 30172
rect -65511 29896 -65139 29928
rect -64511 30172 -64139 30204
rect -64511 29928 -64447 30172
rect -64203 29928 -64139 30172
rect -64511 29896 -64139 29928
rect -63511 30172 -63139 30204
rect -63511 29928 -63447 30172
rect -63203 29928 -63139 30172
rect -63511 29896 -63139 29928
rect -62511 30172 -62139 30204
rect -62511 29928 -62447 30172
rect -62203 29928 -62139 30172
rect -62511 29896 -62139 29928
rect -61511 30172 -61139 30204
rect -61511 29928 -61447 30172
rect -61203 29928 -61139 30172
rect -61511 29896 -61139 29928
rect -60511 30172 -60139 30204
rect -60511 29928 -60447 30172
rect -60203 29928 -60139 30172
rect -60511 29896 -60139 29928
rect -59511 30172 -59139 30204
rect -59511 29928 -59447 30172
rect -59203 29928 -59139 30172
rect -59511 29896 -59139 29928
rect -58831 29896 -58825 30204
rect -74825 29890 -58825 29896
rect -50461 30204 34654 30210
rect -50461 29896 9660 30204
rect 9968 30172 10340 30204
rect 9968 29928 10032 30172
rect 10276 29928 10340 30172
rect 9968 29896 10340 29928
rect 10968 30172 11340 30204
rect 10968 29928 11032 30172
rect 11276 29928 11340 30172
rect 10968 29896 11340 29928
rect 11968 30172 12340 30204
rect 11968 29928 12032 30172
rect 12276 29928 12340 30172
rect 11968 29896 12340 29928
rect 12968 30172 13340 30204
rect 12968 29928 13032 30172
rect 13276 29928 13340 30172
rect 12968 29896 13340 29928
rect 13968 30172 14340 30204
rect 13968 29928 14032 30172
rect 14276 29928 14340 30172
rect 13968 29896 14340 29928
rect 14968 30172 15340 30204
rect 14968 29928 15032 30172
rect 15276 29928 15340 30172
rect 14968 29896 15340 29928
rect 15968 30172 16340 30204
rect 15968 29928 16032 30172
rect 16276 29928 16340 30172
rect 15968 29896 16340 29928
rect 16968 30172 17340 30204
rect 16968 29928 17032 30172
rect 17276 29928 17340 30172
rect 16968 29896 17340 29928
rect 17968 30172 18340 30204
rect 17968 29928 18032 30172
rect 18276 29928 18340 30172
rect 17968 29896 18340 29928
rect 18968 30172 19340 30204
rect 18968 29928 19032 30172
rect 19276 29928 19340 30172
rect 18968 29896 19340 29928
rect 19968 30172 20340 30204
rect 19968 29928 20032 30172
rect 20276 29928 20340 30172
rect 19968 29896 20340 29928
rect 20968 30172 21340 30204
rect 20968 29928 21032 30172
rect 21276 29928 21340 30172
rect 20968 29896 21340 29928
rect 21968 30172 22340 30204
rect 21968 29928 22032 30172
rect 22276 29928 22340 30172
rect 21968 29896 22340 29928
rect 22968 30172 23340 30204
rect 22968 29928 23032 30172
rect 23276 29928 23340 30172
rect 22968 29896 23340 29928
rect 23968 30172 24340 30204
rect 23968 29928 24032 30172
rect 24276 29928 24340 30172
rect 23968 29896 24340 29928
rect 24968 30172 25340 30204
rect 24968 29928 25032 30172
rect 25276 29928 25340 30172
rect 24968 29896 25340 29928
rect 25968 30172 26340 30204
rect 25968 29928 26032 30172
rect 26276 29928 26340 30172
rect 25968 29896 26340 29928
rect 26968 30172 27340 30204
rect 26968 29928 27032 30172
rect 27276 29928 27340 30172
rect 26968 29896 27340 29928
rect 27968 30172 28340 30204
rect 27968 29928 28032 30172
rect 28276 29928 28340 30172
rect 27968 29896 28340 29928
rect 28968 30172 29340 30204
rect 28968 29928 29032 30172
rect 29276 29928 29340 30172
rect 28968 29896 29340 29928
rect 29968 30172 30340 30204
rect 29968 29928 30032 30172
rect 30276 29928 30340 30172
rect 29968 29896 30340 29928
rect 30968 30172 31340 30204
rect 30968 29928 31032 30172
rect 31276 29928 31340 30172
rect 30968 29896 31340 29928
rect 31968 30172 32340 30204
rect 31968 29928 32032 30172
rect 32276 29928 32340 30172
rect 31968 29896 32340 29928
rect 32968 30172 33340 30204
rect 32968 29928 33032 30172
rect 33276 29928 33340 30172
rect 32968 29896 33340 29928
rect 33968 30172 34340 30204
rect 33968 29928 34032 30172
rect 34276 29928 34340 30172
rect 33968 29896 34340 29928
rect 34648 29896 34654 30204
rect -50461 29890 34654 29896
rect -74485 29864 -74165 29890
rect -74485 29236 -74479 29864
rect -74171 29236 -74165 29864
rect -74485 29210 -74165 29236
rect -73485 29864 -73165 29890
rect -73485 29236 -73479 29864
rect -73171 29236 -73165 29864
rect -73485 29210 -73165 29236
rect -72485 29864 -72165 29890
rect -72485 29236 -72479 29864
rect -72171 29236 -72165 29864
rect -72485 29210 -72165 29236
rect -71485 29864 -71165 29890
rect -71485 29236 -71479 29864
rect -71171 29236 -71165 29864
rect -71485 29210 -71165 29236
rect -70485 29864 -70165 29890
rect -70485 29236 -70479 29864
rect -70171 29236 -70165 29864
rect -70485 29210 -70165 29236
rect -69485 29864 -69165 29890
rect -69485 29236 -69479 29864
rect -69171 29236 -69165 29864
rect -69485 29210 -69165 29236
rect -68485 29864 -68165 29890
rect -68485 29236 -68479 29864
rect -68171 29236 -68165 29864
rect -68485 29210 -68165 29236
rect -67485 29864 -67165 29890
rect -67485 29236 -67479 29864
rect -67171 29236 -67165 29864
rect -67485 29210 -67165 29236
rect -66485 29864 -66165 29890
rect -66485 29236 -66479 29864
rect -66171 29236 -66165 29864
rect -66485 29210 -66165 29236
rect -65485 29864 -65165 29890
rect -65485 29236 -65479 29864
rect -65171 29236 -65165 29864
rect -65485 29210 -65165 29236
rect -64485 29864 -64165 29890
rect -64485 29236 -64479 29864
rect -64171 29236 -64165 29864
rect -64485 29210 -64165 29236
rect -63485 29864 -63165 29890
rect -63485 29236 -63479 29864
rect -63171 29236 -63165 29864
rect -63485 29210 -63165 29236
rect -62485 29864 -62165 29890
rect -62485 29236 -62479 29864
rect -62171 29236 -62165 29864
rect -62485 29210 -62165 29236
rect -61485 29864 -61165 29890
rect -61485 29236 -61479 29864
rect -61171 29236 -61165 29864
rect -61485 29210 -61165 29236
rect -60485 29864 -60165 29890
rect -60485 29236 -60479 29864
rect -60171 29236 -60165 29864
rect -60485 29210 -60165 29236
rect -59485 29864 -59165 29890
rect -59485 29236 -59479 29864
rect -59171 29236 -59165 29864
rect -59485 29210 -59165 29236
rect -50461 29210 9654 29890
rect 9994 29864 10314 29890
rect 9994 29236 10000 29864
rect 10308 29236 10314 29864
rect 9994 29210 10314 29236
rect 10994 29864 11314 29890
rect 10994 29236 11000 29864
rect 11308 29236 11314 29864
rect 10994 29210 11314 29236
rect 11994 29864 12314 29890
rect 11994 29236 12000 29864
rect 12308 29236 12314 29864
rect 11994 29210 12314 29236
rect 12994 29864 13314 29890
rect 12994 29236 13000 29864
rect 13308 29236 13314 29864
rect 12994 29210 13314 29236
rect 13994 29864 14314 29890
rect 13994 29236 14000 29864
rect 14308 29236 14314 29864
rect 13994 29210 14314 29236
rect 14994 29864 15314 29890
rect 14994 29236 15000 29864
rect 15308 29236 15314 29864
rect 14994 29210 15314 29236
rect 15994 29864 16314 29890
rect 15994 29236 16000 29864
rect 16308 29236 16314 29864
rect 15994 29210 16314 29236
rect 16994 29864 17314 29890
rect 16994 29236 17000 29864
rect 17308 29236 17314 29864
rect 16994 29210 17314 29236
rect 17994 29864 18314 29890
rect 17994 29236 18000 29864
rect 18308 29236 18314 29864
rect 17994 29210 18314 29236
rect 18994 29864 19314 29890
rect 18994 29236 19000 29864
rect 19308 29236 19314 29864
rect 18994 29210 19314 29236
rect 19994 29864 20314 29890
rect 19994 29236 20000 29864
rect 20308 29236 20314 29864
rect 19994 29210 20314 29236
rect 20994 29864 21314 29890
rect 20994 29236 21000 29864
rect 21308 29236 21314 29864
rect 20994 29210 21314 29236
rect 21994 29864 22314 29890
rect 21994 29236 22000 29864
rect 22308 29236 22314 29864
rect 21994 29210 22314 29236
rect 22994 29864 23314 29890
rect 22994 29236 23000 29864
rect 23308 29236 23314 29864
rect 22994 29210 23314 29236
rect 23994 29864 24314 29890
rect 23994 29236 24000 29864
rect 24308 29236 24314 29864
rect 23994 29210 24314 29236
rect 24994 29864 25314 29890
rect 24994 29236 25000 29864
rect 25308 29236 25314 29864
rect 24994 29210 25314 29236
rect 25994 29864 26314 29890
rect 25994 29236 26000 29864
rect 26308 29236 26314 29864
rect 25994 29210 26314 29236
rect 26994 29864 27314 29890
rect 26994 29236 27000 29864
rect 27308 29236 27314 29864
rect 26994 29210 27314 29236
rect 27994 29864 28314 29890
rect 27994 29236 28000 29864
rect 28308 29236 28314 29864
rect 27994 29210 28314 29236
rect 28994 29864 29314 29890
rect 28994 29236 29000 29864
rect 29308 29236 29314 29864
rect 28994 29210 29314 29236
rect 29994 29864 30314 29890
rect 29994 29236 30000 29864
rect 30308 29236 30314 29864
rect 29994 29210 30314 29236
rect 30994 29864 31314 29890
rect 30994 29236 31000 29864
rect 31308 29236 31314 29864
rect 30994 29210 31314 29236
rect 31994 29864 32314 29890
rect 31994 29236 32000 29864
rect 32308 29236 32314 29864
rect 31994 29210 32314 29236
rect 32994 29864 33314 29890
rect 32994 29236 33000 29864
rect 33308 29236 33314 29864
rect 32994 29210 33314 29236
rect 33994 29864 34314 29890
rect 33994 29236 34000 29864
rect 34308 29236 34314 29864
rect 33994 29210 34314 29236
rect -74825 29204 -58825 29210
rect -74825 28896 -74819 29204
rect -74511 29172 -74139 29204
rect -74511 28928 -74447 29172
rect -74203 28928 -74139 29172
rect -74511 28896 -74139 28928
rect -73511 29172 -73139 29204
rect -73511 28928 -73447 29172
rect -73203 28928 -73139 29172
rect -73511 28896 -73139 28928
rect -72511 29172 -72139 29204
rect -72511 28928 -72447 29172
rect -72203 28928 -72139 29172
rect -72511 28896 -72139 28928
rect -71511 29172 -71139 29204
rect -71511 28928 -71447 29172
rect -71203 28928 -71139 29172
rect -71511 28896 -71139 28928
rect -70511 29172 -70139 29204
rect -70511 28928 -70447 29172
rect -70203 28928 -70139 29172
rect -70511 28896 -70139 28928
rect -69511 29172 -69139 29204
rect -69511 28928 -69447 29172
rect -69203 28928 -69139 29172
rect -69511 28896 -69139 28928
rect -68511 29172 -68139 29204
rect -68511 28928 -68447 29172
rect -68203 28928 -68139 29172
rect -68511 28896 -68139 28928
rect -67511 29172 -67139 29204
rect -67511 28928 -67447 29172
rect -67203 28928 -67139 29172
rect -67511 28896 -67139 28928
rect -66511 29172 -66139 29204
rect -66511 28928 -66447 29172
rect -66203 28928 -66139 29172
rect -66511 28896 -66139 28928
rect -65511 29172 -65139 29204
rect -65511 28928 -65447 29172
rect -65203 28928 -65139 29172
rect -65511 28896 -65139 28928
rect -64511 29172 -64139 29204
rect -64511 28928 -64447 29172
rect -64203 28928 -64139 29172
rect -64511 28896 -64139 28928
rect -63511 29172 -63139 29204
rect -63511 28928 -63447 29172
rect -63203 28928 -63139 29172
rect -63511 28896 -63139 28928
rect -62511 29172 -62139 29204
rect -62511 28928 -62447 29172
rect -62203 28928 -62139 29172
rect -62511 28896 -62139 28928
rect -61511 29172 -61139 29204
rect -61511 28928 -61447 29172
rect -61203 28928 -61139 29172
rect -61511 28896 -61139 28928
rect -60511 29172 -60139 29204
rect -60511 28928 -60447 29172
rect -60203 28928 -60139 29172
rect -60511 28896 -60139 28928
rect -59511 29172 -59139 29204
rect -59511 28928 -59447 29172
rect -59203 28928 -59139 29172
rect -59511 28896 -59139 28928
rect -58831 28896 -58825 29204
rect -74825 28890 -58825 28896
rect -50461 29204 34654 29210
rect -50461 28896 9660 29204
rect 9968 29172 10340 29204
rect 9968 28928 10032 29172
rect 10276 28928 10340 29172
rect 9968 28896 10340 28928
rect 10968 29172 11340 29204
rect 10968 28928 11032 29172
rect 11276 28928 11340 29172
rect 10968 28896 11340 28928
rect 11968 29172 12340 29204
rect 11968 28928 12032 29172
rect 12276 28928 12340 29172
rect 11968 28896 12340 28928
rect 12968 29172 13340 29204
rect 12968 28928 13032 29172
rect 13276 28928 13340 29172
rect 12968 28896 13340 28928
rect 13968 29172 14340 29204
rect 13968 28928 14032 29172
rect 14276 28928 14340 29172
rect 13968 28896 14340 28928
rect 14968 29172 15340 29204
rect 14968 28928 15032 29172
rect 15276 28928 15340 29172
rect 14968 28896 15340 28928
rect 15968 29172 16340 29204
rect 15968 28928 16032 29172
rect 16276 28928 16340 29172
rect 15968 28896 16340 28928
rect 16968 29172 17340 29204
rect 16968 28928 17032 29172
rect 17276 28928 17340 29172
rect 16968 28896 17340 28928
rect 17968 29172 18340 29204
rect 17968 28928 18032 29172
rect 18276 28928 18340 29172
rect 17968 28896 18340 28928
rect 18968 29172 19340 29204
rect 18968 28928 19032 29172
rect 19276 28928 19340 29172
rect 18968 28896 19340 28928
rect 19968 29172 20340 29204
rect 19968 28928 20032 29172
rect 20276 28928 20340 29172
rect 19968 28896 20340 28928
rect 20968 29172 21340 29204
rect 20968 28928 21032 29172
rect 21276 28928 21340 29172
rect 20968 28896 21340 28928
rect 21968 29172 22340 29204
rect 21968 28928 22032 29172
rect 22276 28928 22340 29172
rect 21968 28896 22340 28928
rect 22968 29172 23340 29204
rect 22968 28928 23032 29172
rect 23276 28928 23340 29172
rect 22968 28896 23340 28928
rect 23968 29172 24340 29204
rect 23968 28928 24032 29172
rect 24276 28928 24340 29172
rect 23968 28896 24340 28928
rect 24968 29172 25340 29204
rect 24968 28928 25032 29172
rect 25276 28928 25340 29172
rect 24968 28896 25340 28928
rect 25968 29172 26340 29204
rect 25968 28928 26032 29172
rect 26276 28928 26340 29172
rect 25968 28896 26340 28928
rect 26968 29172 27340 29204
rect 26968 28928 27032 29172
rect 27276 28928 27340 29172
rect 26968 28896 27340 28928
rect 27968 29172 28340 29204
rect 27968 28928 28032 29172
rect 28276 28928 28340 29172
rect 27968 28896 28340 28928
rect 28968 29172 29340 29204
rect 28968 28928 29032 29172
rect 29276 28928 29340 29172
rect 28968 28896 29340 28928
rect 29968 29172 30340 29204
rect 29968 28928 30032 29172
rect 30276 28928 30340 29172
rect 29968 28896 30340 28928
rect 30968 29172 31340 29204
rect 30968 28928 31032 29172
rect 31276 28928 31340 29172
rect 30968 28896 31340 28928
rect 31968 29172 32340 29204
rect 31968 28928 32032 29172
rect 32276 28928 32340 29172
rect 31968 28896 32340 28928
rect 32968 29172 33340 29204
rect 32968 28928 33032 29172
rect 33276 28928 33340 29172
rect 32968 28896 33340 28928
rect 33968 29172 34340 29204
rect 33968 28928 34032 29172
rect 34276 28928 34340 29172
rect 33968 28896 34340 28928
rect 34648 28896 34654 29204
rect -50461 28890 34654 28896
rect -74485 28864 -74165 28890
rect -74485 28556 -74479 28864
rect -74171 28556 -74165 28864
rect -74485 28550 -74165 28556
rect -73485 28864 -73165 28890
rect -73485 28556 -73479 28864
rect -73171 28556 -73165 28864
rect -73485 28550 -73165 28556
rect -72485 28864 -72165 28890
rect -72485 28556 -72479 28864
rect -72171 28556 -72165 28864
rect -72485 28550 -72165 28556
rect -71485 28864 -71165 28890
rect -71485 28556 -71479 28864
rect -71171 28556 -71165 28864
rect -71485 28550 -71165 28556
rect -70485 28864 -70165 28890
rect -70485 28556 -70479 28864
rect -70171 28556 -70165 28864
rect -70485 28550 -70165 28556
rect -69485 28864 -69165 28890
rect -69485 28556 -69479 28864
rect -69171 28556 -69165 28864
rect -69485 28550 -69165 28556
rect -68485 28864 -68165 28890
rect -68485 28556 -68479 28864
rect -68171 28556 -68165 28864
rect -68485 28550 -68165 28556
rect -67485 28864 -67165 28890
rect -67485 28556 -67479 28864
rect -67171 28556 -67165 28864
rect -67485 28550 -67165 28556
rect -66485 28864 -66165 28890
rect -66485 28556 -66479 28864
rect -66171 28556 -66165 28864
rect -66485 28550 -66165 28556
rect -65485 28864 -65165 28890
rect -65485 28556 -65479 28864
rect -65171 28556 -65165 28864
rect -65485 28550 -65165 28556
rect -64485 28864 -64165 28890
rect -64485 28556 -64479 28864
rect -64171 28556 -64165 28864
rect -64485 28550 -64165 28556
rect -63485 28864 -63165 28890
rect -63485 28556 -63479 28864
rect -63171 28556 -63165 28864
rect -63485 28550 -63165 28556
rect -62485 28864 -62165 28890
rect -62485 28556 -62479 28864
rect -62171 28556 -62165 28864
rect -62485 28550 -62165 28556
rect -61485 28864 -61165 28890
rect -61485 28556 -61479 28864
rect -61171 28556 -61165 28864
rect -61485 28550 -61165 28556
rect -60485 28864 -60165 28890
rect -60485 28556 -60479 28864
rect -60171 28556 -60165 28864
rect -60485 28550 -60165 28556
rect -59485 28864 -59165 28890
rect -59485 28556 -59479 28864
rect -59171 28556 -59165 28864
rect -59485 28550 -59165 28556
rect -50461 28000 9654 28890
rect 9994 28864 10314 28890
rect 9994 28556 10000 28864
rect 10308 28556 10314 28864
rect 9994 28550 10314 28556
rect 10994 28864 11314 28890
rect 10994 28556 11000 28864
rect 11308 28556 11314 28864
rect 10994 28550 11314 28556
rect 11994 28864 12314 28890
rect 11994 28556 12000 28864
rect 12308 28556 12314 28864
rect 11994 28550 12314 28556
rect 12994 28864 13314 28890
rect 12994 28556 13000 28864
rect 13308 28556 13314 28864
rect 12994 28550 13314 28556
rect 13994 28864 14314 28890
rect 13994 28556 14000 28864
rect 14308 28556 14314 28864
rect 13994 28550 14314 28556
rect 14994 28864 15314 28890
rect 14994 28556 15000 28864
rect 15308 28556 15314 28864
rect 14994 28550 15314 28556
rect 15994 28864 16314 28890
rect 15994 28556 16000 28864
rect 16308 28556 16314 28864
rect 15994 28550 16314 28556
rect 16994 28864 17314 28890
rect 16994 28556 17000 28864
rect 17308 28556 17314 28864
rect 16994 28550 17314 28556
rect 17994 28864 18314 28890
rect 17994 28556 18000 28864
rect 18308 28556 18314 28864
rect 17994 28550 18314 28556
rect 18994 28864 19314 28890
rect 18994 28556 19000 28864
rect 19308 28556 19314 28864
rect 18994 28550 19314 28556
rect 19994 28864 20314 28890
rect 19994 28556 20000 28864
rect 20308 28556 20314 28864
rect 19994 28550 20314 28556
rect 20994 28864 21314 28890
rect 20994 28556 21000 28864
rect 21308 28556 21314 28864
rect 20994 28550 21314 28556
rect 21994 28864 22314 28890
rect 21994 28556 22000 28864
rect 22308 28556 22314 28864
rect 21994 28550 22314 28556
rect 22994 28864 23314 28890
rect 22994 28556 23000 28864
rect 23308 28556 23314 28864
rect 22994 28550 23314 28556
rect 23994 28864 24314 28890
rect 23994 28556 24000 28864
rect 24308 28556 24314 28864
rect 23994 28550 24314 28556
rect 24994 28864 25314 28890
rect 24994 28556 25000 28864
rect 25308 28556 25314 28864
rect 24994 28550 25314 28556
rect 25994 28864 26314 28890
rect 25994 28556 26000 28864
rect 26308 28556 26314 28864
rect 25994 28550 26314 28556
rect 26994 28864 27314 28890
rect 26994 28556 27000 28864
rect 27308 28556 27314 28864
rect 26994 28550 27314 28556
rect 27994 28864 28314 28890
rect 27994 28556 28000 28864
rect 28308 28556 28314 28864
rect 27994 28550 28314 28556
rect 28994 28864 29314 28890
rect 28994 28556 29000 28864
rect 29308 28556 29314 28864
rect 28994 28550 29314 28556
rect 29994 28864 30314 28890
rect 29994 28556 30000 28864
rect 30308 28556 30314 28864
rect 29994 28550 30314 28556
rect 30994 28864 31314 28890
rect 30994 28556 31000 28864
rect 31308 28556 31314 28864
rect 30994 28550 31314 28556
rect 31994 28864 32314 28890
rect 31994 28556 32000 28864
rect 32308 28556 32314 28864
rect 31994 28550 32314 28556
rect 32994 28864 33314 28890
rect 32994 28556 33000 28864
rect 33308 28556 33314 28864
rect 32994 28550 33314 28556
rect 33994 28864 34314 28890
rect 33994 28556 34000 28864
rect 34308 28556 34314 28864
rect 33994 28550 34314 28556
rect -47613 26087 -47037 26093
rect -72825 25949 -60825 26000
rect -72825 16041 -72776 25949
rect -60884 16041 -60825 25949
rect -47613 25523 -47607 26087
rect -47043 25523 -47037 26087
rect -47613 25517 -47037 25523
rect -47396 24973 -47254 25517
rect -47396 24939 -47340 24973
rect -47306 24939 -47254 24973
rect -47396 24901 -47254 24939
rect -47396 24867 -47340 24901
rect -47306 24867 -47254 24901
rect -47396 24829 -47254 24867
rect -47396 24795 -47340 24829
rect -47306 24795 -47254 24829
rect -47396 24757 -47254 24795
rect -47396 24723 -47340 24757
rect -47306 24723 -47254 24757
rect -47396 24692 -47254 24723
rect -72825 7600 -60825 16041
rect -21272 15124 -19272 28000
rect 6632 26131 7208 26137
rect 6632 25567 6638 26131
rect 7202 25567 7208 26131
rect 6632 25561 7208 25567
rect 20275 25954 32275 26000
rect 6824 24953 6966 25561
rect 6824 24919 6874 24953
rect 6908 24919 6966 24953
rect 6824 24881 6966 24919
rect 6824 24847 6874 24881
rect 6908 24847 6966 24881
rect 6824 24809 6966 24847
rect 6824 24775 6874 24809
rect 6908 24775 6966 24809
rect 6824 24737 6966 24775
rect 6824 24703 6874 24737
rect 6908 24703 6966 24737
rect 6824 24692 6966 24703
rect -21272 13856 -21212 15124
rect -19304 13856 -19272 15124
rect -21272 13850 -19272 13856
rect 20275 16046 20324 25954
rect 32216 16046 32275 25954
rect -72825 -7600 -71325 7600
rect -70525 -7600 -69025 7600
rect -68225 -7600 -66725 7600
rect -65925 -7600 -64425 7600
rect -63625 -7600 -62125 7600
rect -72825 -16046 -60825 -7600
rect -57085 -13850 -57015 13850
rect -56425 -13850 -56355 13850
rect -55765 -13850 -55695 13850
rect -55105 -13850 -55035 13850
rect -54445 -13850 -54375 13850
rect -53785 -13850 -53715 13850
rect -53125 -13850 -53055 13850
rect -52465 -13850 -52395 13850
rect -51805 -13850 -51735 13850
rect -51145 -13850 -51075 13850
rect -50485 -13850 -50415 13850
rect -49825 -13850 -49755 13850
rect -49165 -13850 -49095 13850
rect -48505 -13850 -48435 13850
rect -47845 -13850 -47775 13850
rect -47185 -13850 -47115 13850
rect -46525 -13850 -46455 13850
rect -45865 -13850 -45795 13850
rect -45205 -13850 -45135 13850
rect -44545 -13850 -44475 13850
rect -43885 -13850 -43815 13850
rect -43225 -13850 -43155 13850
rect -42440 13820 -40660 13850
rect -42440 7880 -42408 13820
rect -40692 7880 -40660 13820
rect -42440 5808 -40660 7880
rect -42530 5734 -40660 5808
rect 110 13820 1890 13850
rect 110 7880 142 13820
rect 1858 7880 1890 13820
rect 110 5938 1890 7880
rect 110 5734 1970 5938
rect -42530 5631 -40756 5734
rect -42530 5414 -42484 5631
rect -42530 5380 -42524 5414
rect -42490 5380 -42484 5414
rect -42530 5342 -42484 5380
rect -42530 5308 -42524 5342
rect -42490 5308 -42484 5342
rect -42530 5270 -42484 5308
rect -42530 5236 -42524 5270
rect -42490 5236 -42484 5270
rect -42530 5198 -42484 5236
rect -42530 5164 -42524 5198
rect -42490 5164 -42484 5198
rect -42530 5126 -42484 5164
rect -42530 5092 -42524 5126
rect -42490 5092 -42484 5126
rect -42530 5054 -42484 5092
rect -42530 5020 -42524 5054
rect -42490 5020 -42484 5054
rect -42530 4982 -42484 5020
rect -42530 4948 -42524 4982
rect -42490 4948 -42484 4982
rect -42530 4910 -42484 4948
rect -42530 4876 -42524 4910
rect -42490 4876 -42484 4910
rect -42530 4838 -42484 4876
rect -42530 4804 -42524 4838
rect -42490 4804 -42484 4838
rect -42530 4766 -42484 4804
rect -42530 4732 -42524 4766
rect -42490 4732 -42484 4766
rect -42530 4694 -42484 4732
rect -42530 4660 -42524 4694
rect -42490 4660 -42484 4694
rect -42530 4637 -42484 4660
rect -42434 5414 -42388 5437
rect -42434 5380 -42428 5414
rect -42394 5380 -42388 5414
rect -42434 5342 -42388 5380
rect -42434 5308 -42428 5342
rect -42394 5308 -42388 5342
rect -42434 5270 -42388 5308
rect -42434 5236 -42428 5270
rect -42394 5236 -42388 5270
rect -42434 5198 -42388 5236
rect -42434 5164 -42428 5198
rect -42394 5164 -42388 5198
rect -42434 5126 -42388 5164
rect -42434 5092 -42428 5126
rect -42394 5092 -42388 5126
rect -42434 5054 -42388 5092
rect -42434 5020 -42428 5054
rect -42394 5020 -42388 5054
rect -42434 4982 -42388 5020
rect -42434 4948 -42428 4982
rect -42394 4948 -42388 4982
rect -42434 4910 -42388 4948
rect -42434 4876 -42428 4910
rect -42394 4876 -42388 4910
rect -42434 4838 -42388 4876
rect -42434 4804 -42428 4838
rect -42394 4804 -42388 4838
rect -42434 4766 -42388 4804
rect -42434 4732 -42428 4766
rect -42394 4732 -42388 4766
rect -42434 4694 -42388 4732
rect -42434 4660 -42428 4694
rect -42394 4660 -42388 4694
rect -42434 4374 -42388 4660
rect -42338 5414 -42292 5631
rect -42338 5380 -42332 5414
rect -42298 5380 -42292 5414
rect -42338 5342 -42292 5380
rect -42338 5308 -42332 5342
rect -42298 5308 -42292 5342
rect -42338 5270 -42292 5308
rect -42338 5236 -42332 5270
rect -42298 5236 -42292 5270
rect -42338 5198 -42292 5236
rect -42338 5164 -42332 5198
rect -42298 5164 -42292 5198
rect -42338 5126 -42292 5164
rect -42338 5092 -42332 5126
rect -42298 5092 -42292 5126
rect -42338 5054 -42292 5092
rect -42338 5020 -42332 5054
rect -42298 5020 -42292 5054
rect -42338 4982 -42292 5020
rect -42338 4948 -42332 4982
rect -42298 4948 -42292 4982
rect -42338 4910 -42292 4948
rect -42338 4876 -42332 4910
rect -42298 4876 -42292 4910
rect -42338 4838 -42292 4876
rect -42338 4804 -42332 4838
rect -42298 4804 -42292 4838
rect -42338 4766 -42292 4804
rect -42338 4732 -42332 4766
rect -42298 4732 -42292 4766
rect -42338 4694 -42292 4732
rect -42338 4660 -42332 4694
rect -42298 4660 -42292 4694
rect -42338 4637 -42292 4660
rect -42242 5414 -42196 5437
rect -42242 5380 -42236 5414
rect -42202 5380 -42196 5414
rect -42242 5342 -42196 5380
rect -42242 5308 -42236 5342
rect -42202 5308 -42196 5342
rect -42242 5270 -42196 5308
rect -42242 5236 -42236 5270
rect -42202 5236 -42196 5270
rect -42242 5198 -42196 5236
rect -42242 5164 -42236 5198
rect -42202 5164 -42196 5198
rect -42242 5126 -42196 5164
rect -42242 5092 -42236 5126
rect -42202 5092 -42196 5126
rect -42242 5054 -42196 5092
rect -42242 5020 -42236 5054
rect -42202 5020 -42196 5054
rect -42242 4982 -42196 5020
rect -42242 4948 -42236 4982
rect -42202 4948 -42196 4982
rect -42242 4910 -42196 4948
rect -42242 4876 -42236 4910
rect -42202 4876 -42196 4910
rect -42242 4838 -42196 4876
rect -42242 4804 -42236 4838
rect -42202 4804 -42196 4838
rect -42242 4766 -42196 4804
rect -42242 4732 -42236 4766
rect -42202 4732 -42196 4766
rect -42242 4694 -42196 4732
rect -42242 4660 -42236 4694
rect -42202 4660 -42196 4694
rect -42242 4374 -42196 4660
rect -42146 5414 -42100 5631
rect -42146 5380 -42140 5414
rect -42106 5380 -42100 5414
rect -42146 5342 -42100 5380
rect -42146 5308 -42140 5342
rect -42106 5308 -42100 5342
rect -42146 5270 -42100 5308
rect -42146 5236 -42140 5270
rect -42106 5236 -42100 5270
rect -42146 5198 -42100 5236
rect -42146 5164 -42140 5198
rect -42106 5164 -42100 5198
rect -42146 5126 -42100 5164
rect -42146 5092 -42140 5126
rect -42106 5092 -42100 5126
rect -42146 5054 -42100 5092
rect -42146 5020 -42140 5054
rect -42106 5020 -42100 5054
rect -42146 4982 -42100 5020
rect -42146 4948 -42140 4982
rect -42106 4948 -42100 4982
rect -42146 4910 -42100 4948
rect -42146 4876 -42140 4910
rect -42106 4876 -42100 4910
rect -42146 4838 -42100 4876
rect -42146 4804 -42140 4838
rect -42106 4804 -42100 4838
rect -42146 4766 -42100 4804
rect -42146 4732 -42140 4766
rect -42106 4732 -42100 4766
rect -42146 4694 -42100 4732
rect -42146 4660 -42140 4694
rect -42106 4660 -42100 4694
rect -42146 4637 -42100 4660
rect -42050 5414 -42004 5437
rect -42050 5380 -42044 5414
rect -42010 5380 -42004 5414
rect -42050 5342 -42004 5380
rect -42050 5308 -42044 5342
rect -42010 5308 -42004 5342
rect -42050 5270 -42004 5308
rect -42050 5236 -42044 5270
rect -42010 5236 -42004 5270
rect -42050 5198 -42004 5236
rect -42050 5164 -42044 5198
rect -42010 5164 -42004 5198
rect -42050 5126 -42004 5164
rect -42050 5092 -42044 5126
rect -42010 5092 -42004 5126
rect -42050 5054 -42004 5092
rect -42050 5020 -42044 5054
rect -42010 5020 -42004 5054
rect -42050 4982 -42004 5020
rect -42050 4948 -42044 4982
rect -42010 4948 -42004 4982
rect -42050 4910 -42004 4948
rect -42050 4876 -42044 4910
rect -42010 4876 -42004 4910
rect -42050 4838 -42004 4876
rect -42050 4804 -42044 4838
rect -42010 4804 -42004 4838
rect -42050 4766 -42004 4804
rect -42050 4732 -42044 4766
rect -42010 4732 -42004 4766
rect -42050 4694 -42004 4732
rect -42050 4660 -42044 4694
rect -42010 4660 -42004 4694
rect -42050 4374 -42004 4660
rect -41954 5414 -41908 5631
rect -41954 5380 -41948 5414
rect -41914 5380 -41908 5414
rect -41954 5342 -41908 5380
rect -41954 5308 -41948 5342
rect -41914 5308 -41908 5342
rect -41954 5270 -41908 5308
rect -41954 5236 -41948 5270
rect -41914 5236 -41908 5270
rect -41954 5198 -41908 5236
rect -41954 5164 -41948 5198
rect -41914 5164 -41908 5198
rect -41954 5126 -41908 5164
rect -41954 5092 -41948 5126
rect -41914 5092 -41908 5126
rect -41954 5054 -41908 5092
rect -41954 5020 -41948 5054
rect -41914 5020 -41908 5054
rect -41954 4982 -41908 5020
rect -41954 4948 -41948 4982
rect -41914 4948 -41908 4982
rect -41954 4910 -41908 4948
rect -41954 4876 -41948 4910
rect -41914 4876 -41908 4910
rect -41954 4838 -41908 4876
rect -41954 4804 -41948 4838
rect -41914 4804 -41908 4838
rect -41954 4766 -41908 4804
rect -41954 4732 -41948 4766
rect -41914 4732 -41908 4766
rect -41954 4694 -41908 4732
rect -41954 4660 -41948 4694
rect -41914 4660 -41908 4694
rect -41954 4637 -41908 4660
rect -41858 5414 -41812 5437
rect -41858 5380 -41852 5414
rect -41818 5380 -41812 5414
rect -41858 5342 -41812 5380
rect -41858 5308 -41852 5342
rect -41818 5308 -41812 5342
rect -41858 5270 -41812 5308
rect -41858 5236 -41852 5270
rect -41818 5236 -41812 5270
rect -41858 5198 -41812 5236
rect -41858 5164 -41852 5198
rect -41818 5164 -41812 5198
rect -41858 5126 -41812 5164
rect -41858 5092 -41852 5126
rect -41818 5092 -41812 5126
rect -41858 5054 -41812 5092
rect -41858 5020 -41852 5054
rect -41818 5020 -41812 5054
rect -41858 4982 -41812 5020
rect -41858 4948 -41852 4982
rect -41818 4948 -41812 4982
rect -41858 4910 -41812 4948
rect -41858 4876 -41852 4910
rect -41818 4876 -41812 4910
rect -41858 4838 -41812 4876
rect -41858 4804 -41852 4838
rect -41818 4804 -41812 4838
rect -41858 4766 -41812 4804
rect -41858 4732 -41852 4766
rect -41818 4732 -41812 4766
rect -41858 4694 -41812 4732
rect -41858 4660 -41852 4694
rect -41818 4660 -41812 4694
rect -41858 4374 -41812 4660
rect -41762 5414 -41716 5631
rect -41762 5380 -41756 5414
rect -41722 5380 -41716 5414
rect -41762 5342 -41716 5380
rect -41762 5308 -41756 5342
rect -41722 5308 -41716 5342
rect -41762 5270 -41716 5308
rect -41762 5236 -41756 5270
rect -41722 5236 -41716 5270
rect -41762 5198 -41716 5236
rect -41762 5164 -41756 5198
rect -41722 5164 -41716 5198
rect -41762 5126 -41716 5164
rect -41762 5092 -41756 5126
rect -41722 5092 -41716 5126
rect -41762 5054 -41716 5092
rect -41762 5020 -41756 5054
rect -41722 5020 -41716 5054
rect -41762 4982 -41716 5020
rect -41762 4948 -41756 4982
rect -41722 4948 -41716 4982
rect -41762 4910 -41716 4948
rect -41762 4876 -41756 4910
rect -41722 4876 -41716 4910
rect -41762 4838 -41716 4876
rect -41762 4804 -41756 4838
rect -41722 4804 -41716 4838
rect -41762 4766 -41716 4804
rect -41762 4732 -41756 4766
rect -41722 4732 -41716 4766
rect -41762 4694 -41716 4732
rect -41762 4660 -41756 4694
rect -41722 4660 -41716 4694
rect -41762 4637 -41716 4660
rect -41666 5414 -41620 5437
rect -41666 5380 -41660 5414
rect -41626 5380 -41620 5414
rect -41666 5342 -41620 5380
rect -41666 5308 -41660 5342
rect -41626 5308 -41620 5342
rect -41666 5270 -41620 5308
rect -41666 5236 -41660 5270
rect -41626 5236 -41620 5270
rect -41666 5198 -41620 5236
rect -41666 5164 -41660 5198
rect -41626 5164 -41620 5198
rect -41666 5126 -41620 5164
rect -41666 5092 -41660 5126
rect -41626 5092 -41620 5126
rect -41666 5054 -41620 5092
rect -41666 5020 -41660 5054
rect -41626 5020 -41620 5054
rect -41666 4982 -41620 5020
rect -41666 4948 -41660 4982
rect -41626 4948 -41620 4982
rect -41666 4910 -41620 4948
rect -41666 4876 -41660 4910
rect -41626 4876 -41620 4910
rect -41666 4838 -41620 4876
rect -41666 4804 -41660 4838
rect -41626 4804 -41620 4838
rect -41666 4766 -41620 4804
rect -41666 4732 -41660 4766
rect -41626 4732 -41620 4766
rect -41666 4694 -41620 4732
rect -41666 4660 -41660 4694
rect -41626 4660 -41620 4694
rect -41666 4374 -41620 4660
rect -41570 5414 -41524 5631
rect -41570 5380 -41564 5414
rect -41530 5380 -41524 5414
rect -41570 5342 -41524 5380
rect -41570 5308 -41564 5342
rect -41530 5308 -41524 5342
rect -41570 5270 -41524 5308
rect -41570 5236 -41564 5270
rect -41530 5236 -41524 5270
rect -41570 5198 -41524 5236
rect -41570 5164 -41564 5198
rect -41530 5164 -41524 5198
rect -41570 5126 -41524 5164
rect -41570 5092 -41564 5126
rect -41530 5092 -41524 5126
rect -41570 5054 -41524 5092
rect -41570 5020 -41564 5054
rect -41530 5020 -41524 5054
rect -41570 4982 -41524 5020
rect -41570 4948 -41564 4982
rect -41530 4948 -41524 4982
rect -41570 4910 -41524 4948
rect -41570 4876 -41564 4910
rect -41530 4876 -41524 4910
rect -41570 4838 -41524 4876
rect -41570 4804 -41564 4838
rect -41530 4804 -41524 4838
rect -41570 4766 -41524 4804
rect -41570 4732 -41564 4766
rect -41530 4732 -41524 4766
rect -41570 4694 -41524 4732
rect -41570 4660 -41564 4694
rect -41530 4660 -41524 4694
rect -41570 4637 -41524 4660
rect -41474 5414 -41428 5437
rect -41474 5380 -41468 5414
rect -41434 5380 -41428 5414
rect -41474 5342 -41428 5380
rect -41474 5308 -41468 5342
rect -41434 5308 -41428 5342
rect -41474 5270 -41428 5308
rect -41474 5236 -41468 5270
rect -41434 5236 -41428 5270
rect -41474 5198 -41428 5236
rect -41474 5164 -41468 5198
rect -41434 5164 -41428 5198
rect -41474 5126 -41428 5164
rect -41474 5092 -41468 5126
rect -41434 5092 -41428 5126
rect -41474 5054 -41428 5092
rect -41474 5020 -41468 5054
rect -41434 5020 -41428 5054
rect -41474 4982 -41428 5020
rect -41474 4948 -41468 4982
rect -41434 4948 -41428 4982
rect -41474 4910 -41428 4948
rect -41474 4876 -41468 4910
rect -41434 4876 -41428 4910
rect -41474 4838 -41428 4876
rect -41474 4804 -41468 4838
rect -41434 4804 -41428 4838
rect -41474 4766 -41428 4804
rect -41474 4732 -41468 4766
rect -41434 4732 -41428 4766
rect -41474 4694 -41428 4732
rect -41474 4660 -41468 4694
rect -41434 4660 -41428 4694
rect -41474 4374 -41428 4660
rect -41378 5414 -41332 5631
rect -41378 5380 -41372 5414
rect -41338 5380 -41332 5414
rect -41378 5342 -41332 5380
rect -41378 5308 -41372 5342
rect -41338 5308 -41332 5342
rect -41378 5270 -41332 5308
rect -41378 5236 -41372 5270
rect -41338 5236 -41332 5270
rect -41378 5198 -41332 5236
rect -41378 5164 -41372 5198
rect -41338 5164 -41332 5198
rect -41378 5126 -41332 5164
rect -41378 5092 -41372 5126
rect -41338 5092 -41332 5126
rect -41378 5054 -41332 5092
rect -41378 5020 -41372 5054
rect -41338 5020 -41332 5054
rect -41378 4982 -41332 5020
rect -41378 4948 -41372 4982
rect -41338 4948 -41332 4982
rect -41378 4910 -41332 4948
rect -41378 4876 -41372 4910
rect -41338 4876 -41332 4910
rect -41378 4838 -41332 4876
rect -41378 4804 -41372 4838
rect -41338 4804 -41332 4838
rect -41378 4766 -41332 4804
rect -41378 4732 -41372 4766
rect -41338 4732 -41332 4766
rect -41378 4694 -41332 4732
rect -41378 4660 -41372 4694
rect -41338 4660 -41332 4694
rect -41378 4637 -41332 4660
rect -41282 5414 -41236 5437
rect -41282 5380 -41276 5414
rect -41242 5380 -41236 5414
rect -41282 5342 -41236 5380
rect -41282 5308 -41276 5342
rect -41242 5308 -41236 5342
rect -41282 5270 -41236 5308
rect -41282 5236 -41276 5270
rect -41242 5236 -41236 5270
rect -41282 5198 -41236 5236
rect -41282 5164 -41276 5198
rect -41242 5164 -41236 5198
rect -41282 5126 -41236 5164
rect -41282 5092 -41276 5126
rect -41242 5092 -41236 5126
rect -41282 5054 -41236 5092
rect -41282 5020 -41276 5054
rect -41242 5020 -41236 5054
rect -41282 4982 -41236 5020
rect -41282 4948 -41276 4982
rect -41242 4948 -41236 4982
rect -41282 4910 -41236 4948
rect -41282 4876 -41276 4910
rect -41242 4876 -41236 4910
rect -41282 4838 -41236 4876
rect -41282 4804 -41276 4838
rect -41242 4804 -41236 4838
rect -41282 4766 -41236 4804
rect -41282 4732 -41276 4766
rect -41242 4732 -41236 4766
rect -41282 4694 -41236 4732
rect -41282 4660 -41276 4694
rect -41242 4660 -41236 4694
rect -41282 4374 -41236 4660
rect -41186 5414 -41140 5631
rect -41186 5380 -41180 5414
rect -41146 5380 -41140 5414
rect -41186 5342 -41140 5380
rect -41186 5308 -41180 5342
rect -41146 5308 -41140 5342
rect -41186 5270 -41140 5308
rect -41186 5236 -41180 5270
rect -41146 5236 -41140 5270
rect -41186 5198 -41140 5236
rect -41186 5164 -41180 5198
rect -41146 5164 -41140 5198
rect -41186 5126 -41140 5164
rect -41186 5092 -41180 5126
rect -41146 5092 -41140 5126
rect -41186 5054 -41140 5092
rect -41186 5020 -41180 5054
rect -41146 5020 -41140 5054
rect -41186 4982 -41140 5020
rect -41186 4948 -41180 4982
rect -41146 4948 -41140 4982
rect -41186 4910 -41140 4948
rect -41186 4876 -41180 4910
rect -41146 4876 -41140 4910
rect -41186 4838 -41140 4876
rect -41186 4804 -41180 4838
rect -41146 4804 -41140 4838
rect -41186 4766 -41140 4804
rect -41186 4732 -41180 4766
rect -41146 4732 -41140 4766
rect -41186 4694 -41140 4732
rect -41186 4660 -41180 4694
rect -41146 4660 -41140 4694
rect -41186 4637 -41140 4660
rect -41090 5414 -41044 5437
rect -41090 5380 -41084 5414
rect -41050 5380 -41044 5414
rect -41090 5342 -41044 5380
rect -41090 5308 -41084 5342
rect -41050 5308 -41044 5342
rect -41090 5270 -41044 5308
rect -41090 5236 -41084 5270
rect -41050 5236 -41044 5270
rect -41090 5198 -41044 5236
rect -41090 5164 -41084 5198
rect -41050 5164 -41044 5198
rect -41090 5126 -41044 5164
rect -41090 5092 -41084 5126
rect -41050 5092 -41044 5126
rect -41090 5054 -41044 5092
rect -41090 5020 -41084 5054
rect -41050 5020 -41044 5054
rect -41090 4982 -41044 5020
rect -41090 4948 -41084 4982
rect -41050 4948 -41044 4982
rect -41090 4910 -41044 4948
rect -41090 4876 -41084 4910
rect -41050 4876 -41044 4910
rect -41090 4838 -41044 4876
rect -41090 4804 -41084 4838
rect -41050 4804 -41044 4838
rect -41090 4766 -41044 4804
rect -41090 4732 -41084 4766
rect -41050 4732 -41044 4766
rect -41090 4694 -41044 4732
rect -41090 4660 -41084 4694
rect -41050 4660 -41044 4694
rect -41090 4374 -41044 4660
rect -40994 5414 -40948 5631
rect -40994 5380 -40988 5414
rect -40954 5380 -40948 5414
rect -40994 5342 -40948 5380
rect -40994 5308 -40988 5342
rect -40954 5308 -40948 5342
rect -40994 5270 -40948 5308
rect -40994 5236 -40988 5270
rect -40954 5236 -40948 5270
rect -40994 5198 -40948 5236
rect -40994 5164 -40988 5198
rect -40954 5164 -40948 5198
rect -40994 5126 -40948 5164
rect -40994 5092 -40988 5126
rect -40954 5092 -40948 5126
rect -40994 5054 -40948 5092
rect -40994 5020 -40988 5054
rect -40954 5020 -40948 5054
rect -40994 4982 -40948 5020
rect -40994 4948 -40988 4982
rect -40954 4948 -40948 4982
rect -40994 4910 -40948 4948
rect -40994 4876 -40988 4910
rect -40954 4876 -40948 4910
rect -40994 4838 -40948 4876
rect -40994 4804 -40988 4838
rect -40954 4804 -40948 4838
rect -40994 4766 -40948 4804
rect -40994 4732 -40988 4766
rect -40954 4732 -40948 4766
rect -40994 4694 -40948 4732
rect -40994 4660 -40988 4694
rect -40954 4660 -40948 4694
rect -40994 4637 -40948 4660
rect -40898 5414 -40852 5437
rect -40898 5380 -40892 5414
rect -40858 5380 -40852 5414
rect -40898 5342 -40852 5380
rect -40898 5308 -40892 5342
rect -40858 5308 -40852 5342
rect -40898 5270 -40852 5308
rect -40898 5236 -40892 5270
rect -40858 5236 -40852 5270
rect -40898 5198 -40852 5236
rect -40898 5164 -40892 5198
rect -40858 5164 -40852 5198
rect -40898 5126 -40852 5164
rect -40898 5092 -40892 5126
rect -40858 5092 -40852 5126
rect -40898 5054 -40852 5092
rect -40898 5020 -40892 5054
rect -40858 5020 -40852 5054
rect -40898 4982 -40852 5020
rect -40898 4948 -40892 4982
rect -40858 4948 -40852 4982
rect -40898 4910 -40852 4948
rect -40898 4876 -40892 4910
rect -40858 4876 -40852 4910
rect -40898 4838 -40852 4876
rect -40898 4804 -40892 4838
rect -40858 4804 -40852 4838
rect -40898 4766 -40852 4804
rect -40898 4732 -40892 4766
rect -40858 4732 -40852 4766
rect -40898 4694 -40852 4732
rect -40898 4660 -40892 4694
rect -40858 4660 -40852 4694
rect -40898 4374 -40852 4660
rect -40802 5414 -40756 5631
rect 194 5619 1968 5734
rect -40802 5380 -40796 5414
rect -40762 5380 -40756 5414
rect -40802 5342 -40756 5380
rect -40802 5308 -40796 5342
rect -40762 5308 -40756 5342
rect -40802 5270 -40756 5308
rect -40802 5236 -40796 5270
rect -40762 5236 -40756 5270
rect -40802 5198 -40756 5236
rect -40802 5164 -40796 5198
rect -40762 5164 -40756 5198
rect -40802 5126 -40756 5164
rect -40802 5092 -40796 5126
rect -40762 5092 -40756 5126
rect -40802 5054 -40756 5092
rect -40802 5020 -40796 5054
rect -40762 5020 -40756 5054
rect -40802 4982 -40756 5020
rect -40802 4948 -40796 4982
rect -40762 4948 -40756 4982
rect -40802 4910 -40756 4948
rect -40802 4876 -40796 4910
rect -40762 4876 -40756 4910
rect -40802 4838 -40756 4876
rect -40802 4804 -40796 4838
rect -40762 4804 -40756 4838
rect -40802 4766 -40756 4804
rect -40802 4732 -40796 4766
rect -40762 4732 -40756 4766
rect -40802 4694 -40756 4732
rect -40802 4660 -40796 4694
rect -40762 4660 -40756 4694
rect -40802 4637 -40756 4660
rect -40706 5414 -40660 5437
rect -40706 5380 -40700 5414
rect -40666 5380 -40660 5414
rect -40706 5342 -40660 5380
rect -40706 5308 -40700 5342
rect -40666 5308 -40660 5342
rect -40706 5270 -40660 5308
rect -40706 5236 -40700 5270
rect -40666 5236 -40660 5270
rect -40706 5198 -40660 5236
rect -40706 5164 -40700 5198
rect -40666 5164 -40660 5198
rect -40706 5126 -40660 5164
rect -40706 5092 -40700 5126
rect -40666 5092 -40660 5126
rect -40706 5054 -40660 5092
rect -40706 5020 -40700 5054
rect -40666 5020 -40660 5054
rect -40706 4982 -40660 5020
rect -40706 4948 -40700 4982
rect -40666 4948 -40660 4982
rect -40706 4910 -40660 4948
rect -40706 4876 -40700 4910
rect -40666 4876 -40660 4910
rect -40706 4838 -40660 4876
rect -40706 4804 -40700 4838
rect -40666 4804 -40660 4838
rect -40706 4766 -40660 4804
rect -40706 4732 -40700 4766
rect -40666 4732 -40660 4766
rect -40706 4694 -40660 4732
rect -40706 4660 -40700 4694
rect -40666 4660 -40660 4694
rect -40706 4374 -40660 4660
rect -42434 4240 -40660 4374
rect -42440 2298 -40660 4240
rect 98 5402 144 5430
rect 98 5368 104 5402
rect 138 5368 144 5402
rect 98 5330 144 5368
rect 98 5296 104 5330
rect 138 5296 144 5330
rect 98 5258 144 5296
rect 98 5224 104 5258
rect 138 5224 144 5258
rect 98 5186 144 5224
rect 98 5152 104 5186
rect 138 5152 144 5186
rect 98 5114 144 5152
rect 98 5080 104 5114
rect 138 5080 144 5114
rect 98 5042 144 5080
rect 98 5008 104 5042
rect 138 5008 144 5042
rect 98 4970 144 5008
rect 98 4936 104 4970
rect 138 4936 144 4970
rect 98 4898 144 4936
rect 98 4864 104 4898
rect 138 4864 144 4898
rect 98 4826 144 4864
rect 98 4792 104 4826
rect 138 4792 144 4826
rect 98 4754 144 4792
rect 98 4720 104 4754
rect 138 4720 144 4754
rect 98 4682 144 4720
rect 98 4648 104 4682
rect 138 4648 144 4682
rect 98 4367 144 4648
rect 194 5402 240 5619
rect 194 5368 200 5402
rect 234 5368 240 5402
rect 194 5330 240 5368
rect 194 5296 200 5330
rect 234 5296 240 5330
rect 194 5258 240 5296
rect 194 5224 200 5258
rect 234 5224 240 5258
rect 194 5186 240 5224
rect 194 5152 200 5186
rect 234 5152 240 5186
rect 194 5114 240 5152
rect 194 5080 200 5114
rect 234 5080 240 5114
rect 194 5042 240 5080
rect 194 5008 200 5042
rect 234 5008 240 5042
rect 194 4970 240 5008
rect 194 4936 200 4970
rect 234 4936 240 4970
rect 194 4898 240 4936
rect 194 4864 200 4898
rect 234 4864 240 4898
rect 194 4826 240 4864
rect 194 4792 200 4826
rect 234 4792 240 4826
rect 194 4754 240 4792
rect 194 4720 200 4754
rect 234 4720 240 4754
rect 194 4682 240 4720
rect 194 4648 200 4682
rect 234 4648 240 4682
rect 194 4625 240 4648
rect 290 5402 336 5430
rect 290 5368 296 5402
rect 330 5368 336 5402
rect 290 5330 336 5368
rect 290 5296 296 5330
rect 330 5296 336 5330
rect 290 5258 336 5296
rect 290 5224 296 5258
rect 330 5224 336 5258
rect 290 5186 336 5224
rect 290 5152 296 5186
rect 330 5152 336 5186
rect 290 5114 336 5152
rect 290 5080 296 5114
rect 330 5080 336 5114
rect 290 5042 336 5080
rect 290 5008 296 5042
rect 330 5008 336 5042
rect 290 4970 336 5008
rect 290 4936 296 4970
rect 330 4936 336 4970
rect 290 4898 336 4936
rect 290 4864 296 4898
rect 330 4864 336 4898
rect 290 4826 336 4864
rect 290 4792 296 4826
rect 330 4792 336 4826
rect 290 4754 336 4792
rect 290 4720 296 4754
rect 330 4720 336 4754
rect 290 4682 336 4720
rect 290 4648 296 4682
rect 330 4648 336 4682
rect 290 4367 336 4648
rect 386 5402 432 5619
rect 386 5368 392 5402
rect 426 5368 432 5402
rect 386 5330 432 5368
rect 386 5296 392 5330
rect 426 5296 432 5330
rect 386 5258 432 5296
rect 386 5224 392 5258
rect 426 5224 432 5258
rect 386 5186 432 5224
rect 386 5152 392 5186
rect 426 5152 432 5186
rect 386 5114 432 5152
rect 386 5080 392 5114
rect 426 5080 432 5114
rect 386 5042 432 5080
rect 386 5008 392 5042
rect 426 5008 432 5042
rect 386 4970 432 5008
rect 386 4936 392 4970
rect 426 4936 432 4970
rect 386 4898 432 4936
rect 386 4864 392 4898
rect 426 4864 432 4898
rect 386 4826 432 4864
rect 386 4792 392 4826
rect 426 4792 432 4826
rect 386 4754 432 4792
rect 386 4720 392 4754
rect 426 4720 432 4754
rect 386 4682 432 4720
rect 386 4648 392 4682
rect 426 4648 432 4682
rect 386 4625 432 4648
rect 482 5402 528 5430
rect 482 5368 488 5402
rect 522 5368 528 5402
rect 482 5330 528 5368
rect 482 5296 488 5330
rect 522 5296 528 5330
rect 482 5258 528 5296
rect 482 5224 488 5258
rect 522 5224 528 5258
rect 482 5186 528 5224
rect 482 5152 488 5186
rect 522 5152 528 5186
rect 482 5114 528 5152
rect 482 5080 488 5114
rect 522 5080 528 5114
rect 482 5042 528 5080
rect 482 5008 488 5042
rect 522 5008 528 5042
rect 482 4970 528 5008
rect 482 4936 488 4970
rect 522 4936 528 4970
rect 482 4898 528 4936
rect 482 4864 488 4898
rect 522 4864 528 4898
rect 482 4826 528 4864
rect 482 4792 488 4826
rect 522 4792 528 4826
rect 482 4754 528 4792
rect 482 4720 488 4754
rect 522 4720 528 4754
rect 482 4682 528 4720
rect 482 4648 488 4682
rect 522 4648 528 4682
rect 482 4367 528 4648
rect 578 5402 624 5619
rect 578 5368 584 5402
rect 618 5368 624 5402
rect 578 5330 624 5368
rect 578 5296 584 5330
rect 618 5296 624 5330
rect 578 5258 624 5296
rect 578 5224 584 5258
rect 618 5224 624 5258
rect 578 5186 624 5224
rect 578 5152 584 5186
rect 618 5152 624 5186
rect 578 5114 624 5152
rect 578 5080 584 5114
rect 618 5080 624 5114
rect 578 5042 624 5080
rect 578 5008 584 5042
rect 618 5008 624 5042
rect 578 4970 624 5008
rect 578 4936 584 4970
rect 618 4936 624 4970
rect 578 4898 624 4936
rect 578 4864 584 4898
rect 618 4864 624 4898
rect 578 4826 624 4864
rect 578 4792 584 4826
rect 618 4792 624 4826
rect 578 4754 624 4792
rect 578 4720 584 4754
rect 618 4720 624 4754
rect 578 4682 624 4720
rect 578 4648 584 4682
rect 618 4648 624 4682
rect 578 4625 624 4648
rect 674 5402 720 5430
rect 674 5368 680 5402
rect 714 5368 720 5402
rect 674 5330 720 5368
rect 674 5296 680 5330
rect 714 5296 720 5330
rect 674 5258 720 5296
rect 674 5224 680 5258
rect 714 5224 720 5258
rect 674 5186 720 5224
rect 674 5152 680 5186
rect 714 5152 720 5186
rect 674 5114 720 5152
rect 674 5080 680 5114
rect 714 5080 720 5114
rect 674 5042 720 5080
rect 674 5008 680 5042
rect 714 5008 720 5042
rect 674 4970 720 5008
rect 674 4936 680 4970
rect 714 4936 720 4970
rect 674 4898 720 4936
rect 674 4864 680 4898
rect 714 4864 720 4898
rect 674 4826 720 4864
rect 674 4792 680 4826
rect 714 4792 720 4826
rect 674 4754 720 4792
rect 674 4720 680 4754
rect 714 4720 720 4754
rect 674 4682 720 4720
rect 674 4648 680 4682
rect 714 4648 720 4682
rect 674 4367 720 4648
rect 770 5402 816 5619
rect 770 5368 776 5402
rect 810 5368 816 5402
rect 770 5330 816 5368
rect 770 5296 776 5330
rect 810 5296 816 5330
rect 770 5258 816 5296
rect 770 5224 776 5258
rect 810 5224 816 5258
rect 770 5186 816 5224
rect 770 5152 776 5186
rect 810 5152 816 5186
rect 770 5114 816 5152
rect 770 5080 776 5114
rect 810 5080 816 5114
rect 770 5042 816 5080
rect 770 5008 776 5042
rect 810 5008 816 5042
rect 770 4970 816 5008
rect 770 4936 776 4970
rect 810 4936 816 4970
rect 770 4898 816 4936
rect 770 4864 776 4898
rect 810 4864 816 4898
rect 770 4826 816 4864
rect 770 4792 776 4826
rect 810 4792 816 4826
rect 770 4754 816 4792
rect 770 4720 776 4754
rect 810 4720 816 4754
rect 770 4682 816 4720
rect 770 4648 776 4682
rect 810 4648 816 4682
rect 770 4625 816 4648
rect 866 5402 912 5430
rect 866 5368 872 5402
rect 906 5368 912 5402
rect 866 5330 912 5368
rect 866 5296 872 5330
rect 906 5296 912 5330
rect 866 5258 912 5296
rect 866 5224 872 5258
rect 906 5224 912 5258
rect 866 5186 912 5224
rect 866 5152 872 5186
rect 906 5152 912 5186
rect 866 5114 912 5152
rect 866 5080 872 5114
rect 906 5080 912 5114
rect 866 5042 912 5080
rect 866 5008 872 5042
rect 906 5008 912 5042
rect 866 4970 912 5008
rect 866 4936 872 4970
rect 906 4936 912 4970
rect 866 4898 912 4936
rect 866 4864 872 4898
rect 906 4864 912 4898
rect 866 4826 912 4864
rect 866 4792 872 4826
rect 906 4792 912 4826
rect 866 4754 912 4792
rect 866 4720 872 4754
rect 906 4720 912 4754
rect 866 4682 912 4720
rect 866 4648 872 4682
rect 906 4648 912 4682
rect 866 4367 912 4648
rect 962 5402 1008 5619
rect 962 5368 968 5402
rect 1002 5368 1008 5402
rect 962 5330 1008 5368
rect 962 5296 968 5330
rect 1002 5296 1008 5330
rect 962 5258 1008 5296
rect 962 5224 968 5258
rect 1002 5224 1008 5258
rect 962 5186 1008 5224
rect 962 5152 968 5186
rect 1002 5152 1008 5186
rect 962 5114 1008 5152
rect 962 5080 968 5114
rect 1002 5080 1008 5114
rect 962 5042 1008 5080
rect 962 5008 968 5042
rect 1002 5008 1008 5042
rect 962 4970 1008 5008
rect 962 4936 968 4970
rect 1002 4936 1008 4970
rect 962 4898 1008 4936
rect 962 4864 968 4898
rect 1002 4864 1008 4898
rect 962 4826 1008 4864
rect 962 4792 968 4826
rect 1002 4792 1008 4826
rect 962 4754 1008 4792
rect 962 4720 968 4754
rect 1002 4720 1008 4754
rect 962 4682 1008 4720
rect 962 4648 968 4682
rect 1002 4648 1008 4682
rect 962 4625 1008 4648
rect 1058 5402 1104 5430
rect 1058 5368 1064 5402
rect 1098 5368 1104 5402
rect 1058 5330 1104 5368
rect 1058 5296 1064 5330
rect 1098 5296 1104 5330
rect 1058 5258 1104 5296
rect 1058 5224 1064 5258
rect 1098 5224 1104 5258
rect 1058 5186 1104 5224
rect 1058 5152 1064 5186
rect 1098 5152 1104 5186
rect 1058 5114 1104 5152
rect 1058 5080 1064 5114
rect 1098 5080 1104 5114
rect 1058 5042 1104 5080
rect 1058 5008 1064 5042
rect 1098 5008 1104 5042
rect 1058 4970 1104 5008
rect 1058 4936 1064 4970
rect 1098 4936 1104 4970
rect 1058 4898 1104 4936
rect 1058 4864 1064 4898
rect 1098 4864 1104 4898
rect 1058 4826 1104 4864
rect 1058 4792 1064 4826
rect 1098 4792 1104 4826
rect 1058 4754 1104 4792
rect 1058 4720 1064 4754
rect 1098 4720 1104 4754
rect 1058 4682 1104 4720
rect 1058 4648 1064 4682
rect 1098 4648 1104 4682
rect 1058 4367 1104 4648
rect 1154 5402 1200 5619
rect 1154 5368 1160 5402
rect 1194 5368 1200 5402
rect 1154 5330 1200 5368
rect 1154 5296 1160 5330
rect 1194 5296 1200 5330
rect 1154 5258 1200 5296
rect 1154 5224 1160 5258
rect 1194 5224 1200 5258
rect 1154 5186 1200 5224
rect 1154 5152 1160 5186
rect 1194 5152 1200 5186
rect 1154 5114 1200 5152
rect 1154 5080 1160 5114
rect 1194 5080 1200 5114
rect 1154 5042 1200 5080
rect 1154 5008 1160 5042
rect 1194 5008 1200 5042
rect 1154 4970 1200 5008
rect 1154 4936 1160 4970
rect 1194 4936 1200 4970
rect 1154 4898 1200 4936
rect 1154 4864 1160 4898
rect 1194 4864 1200 4898
rect 1154 4826 1200 4864
rect 1154 4792 1160 4826
rect 1194 4792 1200 4826
rect 1154 4754 1200 4792
rect 1154 4720 1160 4754
rect 1194 4720 1200 4754
rect 1154 4682 1200 4720
rect 1154 4648 1160 4682
rect 1194 4648 1200 4682
rect 1154 4625 1200 4648
rect 1250 5402 1296 5430
rect 1250 5368 1256 5402
rect 1290 5368 1296 5402
rect 1250 5330 1296 5368
rect 1250 5296 1256 5330
rect 1290 5296 1296 5330
rect 1250 5258 1296 5296
rect 1250 5224 1256 5258
rect 1290 5224 1296 5258
rect 1250 5186 1296 5224
rect 1250 5152 1256 5186
rect 1290 5152 1296 5186
rect 1250 5114 1296 5152
rect 1250 5080 1256 5114
rect 1290 5080 1296 5114
rect 1250 5042 1296 5080
rect 1250 5008 1256 5042
rect 1290 5008 1296 5042
rect 1250 4970 1296 5008
rect 1250 4936 1256 4970
rect 1290 4936 1296 4970
rect 1250 4898 1296 4936
rect 1250 4864 1256 4898
rect 1290 4864 1296 4898
rect 1250 4826 1296 4864
rect 1250 4792 1256 4826
rect 1290 4792 1296 4826
rect 1250 4754 1296 4792
rect 1250 4720 1256 4754
rect 1290 4720 1296 4754
rect 1250 4682 1296 4720
rect 1250 4648 1256 4682
rect 1290 4648 1296 4682
rect 1250 4367 1296 4648
rect 1346 5402 1392 5619
rect 1346 5368 1352 5402
rect 1386 5368 1392 5402
rect 1346 5330 1392 5368
rect 1346 5296 1352 5330
rect 1386 5296 1392 5330
rect 1346 5258 1392 5296
rect 1346 5224 1352 5258
rect 1386 5224 1392 5258
rect 1346 5186 1392 5224
rect 1346 5152 1352 5186
rect 1386 5152 1392 5186
rect 1346 5114 1392 5152
rect 1346 5080 1352 5114
rect 1386 5080 1392 5114
rect 1346 5042 1392 5080
rect 1346 5008 1352 5042
rect 1386 5008 1392 5042
rect 1346 4970 1392 5008
rect 1346 4936 1352 4970
rect 1386 4936 1392 4970
rect 1346 4898 1392 4936
rect 1346 4864 1352 4898
rect 1386 4864 1392 4898
rect 1346 4826 1392 4864
rect 1346 4792 1352 4826
rect 1386 4792 1392 4826
rect 1346 4754 1392 4792
rect 1346 4720 1352 4754
rect 1386 4720 1392 4754
rect 1346 4682 1392 4720
rect 1346 4648 1352 4682
rect 1386 4648 1392 4682
rect 1346 4625 1392 4648
rect 1442 5402 1488 5430
rect 1442 5368 1448 5402
rect 1482 5368 1488 5402
rect 1442 5330 1488 5368
rect 1442 5296 1448 5330
rect 1482 5296 1488 5330
rect 1442 5258 1488 5296
rect 1442 5224 1448 5258
rect 1482 5224 1488 5258
rect 1442 5186 1488 5224
rect 1442 5152 1448 5186
rect 1482 5152 1488 5186
rect 1442 5114 1488 5152
rect 1442 5080 1448 5114
rect 1482 5080 1488 5114
rect 1442 5042 1488 5080
rect 1442 5008 1448 5042
rect 1482 5008 1488 5042
rect 1442 4970 1488 5008
rect 1442 4936 1448 4970
rect 1482 4936 1488 4970
rect 1442 4898 1488 4936
rect 1442 4864 1448 4898
rect 1482 4864 1488 4898
rect 1442 4826 1488 4864
rect 1442 4792 1448 4826
rect 1482 4792 1488 4826
rect 1442 4754 1488 4792
rect 1442 4720 1448 4754
rect 1482 4720 1488 4754
rect 1442 4682 1488 4720
rect 1442 4648 1448 4682
rect 1482 4648 1488 4682
rect 1442 4367 1488 4648
rect 1538 5402 1584 5619
rect 1538 5368 1544 5402
rect 1578 5368 1584 5402
rect 1538 5330 1584 5368
rect 1538 5296 1544 5330
rect 1578 5296 1584 5330
rect 1538 5258 1584 5296
rect 1538 5224 1544 5258
rect 1578 5224 1584 5258
rect 1538 5186 1584 5224
rect 1538 5152 1544 5186
rect 1578 5152 1584 5186
rect 1538 5114 1584 5152
rect 1538 5080 1544 5114
rect 1578 5080 1584 5114
rect 1538 5042 1584 5080
rect 1538 5008 1544 5042
rect 1578 5008 1584 5042
rect 1538 4970 1584 5008
rect 1538 4936 1544 4970
rect 1578 4936 1584 4970
rect 1538 4898 1584 4936
rect 1538 4864 1544 4898
rect 1578 4864 1584 4898
rect 1538 4826 1584 4864
rect 1538 4792 1544 4826
rect 1578 4792 1584 4826
rect 1538 4754 1584 4792
rect 1538 4720 1544 4754
rect 1578 4720 1584 4754
rect 1538 4682 1584 4720
rect 1538 4648 1544 4682
rect 1578 4648 1584 4682
rect 1538 4625 1584 4648
rect 1634 5402 1680 5430
rect 1634 5368 1640 5402
rect 1674 5368 1680 5402
rect 1634 5330 1680 5368
rect 1634 5296 1640 5330
rect 1674 5296 1680 5330
rect 1634 5258 1680 5296
rect 1634 5224 1640 5258
rect 1674 5224 1680 5258
rect 1634 5186 1680 5224
rect 1634 5152 1640 5186
rect 1674 5152 1680 5186
rect 1634 5114 1680 5152
rect 1634 5080 1640 5114
rect 1674 5080 1680 5114
rect 1634 5042 1680 5080
rect 1634 5008 1640 5042
rect 1674 5008 1680 5042
rect 1634 4970 1680 5008
rect 1634 4936 1640 4970
rect 1674 4936 1680 4970
rect 1634 4898 1680 4936
rect 1634 4864 1640 4898
rect 1674 4864 1680 4898
rect 1634 4826 1680 4864
rect 1634 4792 1640 4826
rect 1674 4792 1680 4826
rect 1634 4754 1680 4792
rect 1634 4720 1640 4754
rect 1674 4720 1680 4754
rect 1634 4682 1680 4720
rect 1634 4648 1640 4682
rect 1674 4648 1680 4682
rect 1634 4367 1680 4648
rect 1730 5402 1776 5619
rect 1730 5368 1736 5402
rect 1770 5368 1776 5402
rect 1730 5330 1776 5368
rect 1730 5296 1736 5330
rect 1770 5296 1776 5330
rect 1730 5258 1776 5296
rect 1730 5224 1736 5258
rect 1770 5224 1776 5258
rect 1730 5186 1776 5224
rect 1730 5152 1736 5186
rect 1770 5152 1776 5186
rect 1730 5114 1776 5152
rect 1730 5080 1736 5114
rect 1770 5080 1776 5114
rect 1730 5042 1776 5080
rect 1730 5008 1736 5042
rect 1770 5008 1776 5042
rect 1730 4970 1776 5008
rect 1730 4936 1736 4970
rect 1770 4936 1776 4970
rect 1730 4898 1776 4936
rect 1730 4864 1736 4898
rect 1770 4864 1776 4898
rect 1730 4826 1776 4864
rect 1730 4792 1736 4826
rect 1770 4792 1776 4826
rect 1730 4754 1776 4792
rect 1730 4720 1736 4754
rect 1770 4720 1776 4754
rect 1730 4682 1776 4720
rect 1730 4648 1736 4682
rect 1770 4648 1776 4682
rect 1730 4625 1776 4648
rect 1826 5402 1872 5430
rect 1826 5368 1832 5402
rect 1866 5368 1872 5402
rect 1826 5330 1872 5368
rect 1826 5296 1832 5330
rect 1866 5296 1872 5330
rect 1826 5258 1872 5296
rect 1826 5224 1832 5258
rect 1866 5224 1872 5258
rect 1826 5186 1872 5224
rect 1826 5152 1832 5186
rect 1866 5152 1872 5186
rect 1826 5114 1872 5152
rect 1826 5080 1832 5114
rect 1866 5080 1872 5114
rect 1826 5042 1872 5080
rect 1826 5008 1832 5042
rect 1866 5008 1872 5042
rect 1826 4970 1872 5008
rect 1826 4936 1832 4970
rect 1866 4936 1872 4970
rect 1826 4898 1872 4936
rect 1826 4864 1832 4898
rect 1866 4864 1872 4898
rect 1826 4826 1872 4864
rect 1826 4792 1832 4826
rect 1866 4792 1872 4826
rect 1826 4754 1872 4792
rect 1826 4720 1832 4754
rect 1866 4720 1872 4754
rect 1826 4682 1872 4720
rect 1826 4648 1832 4682
rect 1866 4648 1872 4682
rect 1826 4367 1872 4648
rect 1922 5402 1968 5619
rect 1922 5368 1928 5402
rect 1962 5368 1968 5402
rect 1922 5330 1968 5368
rect 1922 5296 1928 5330
rect 1962 5296 1968 5330
rect 1922 5258 1968 5296
rect 1922 5224 1928 5258
rect 1962 5224 1968 5258
rect 1922 5186 1968 5224
rect 1922 5152 1928 5186
rect 1962 5152 1968 5186
rect 1922 5114 1968 5152
rect 1922 5080 1928 5114
rect 1962 5080 1968 5114
rect 1922 5042 1968 5080
rect 1922 5008 1928 5042
rect 1962 5008 1968 5042
rect 1922 4970 1968 5008
rect 1922 4936 1928 4970
rect 1962 4936 1968 4970
rect 1922 4898 1968 4936
rect 1922 4864 1928 4898
rect 1962 4864 1968 4898
rect 1922 4826 1968 4864
rect 1922 4792 1928 4826
rect 1962 4792 1968 4826
rect 1922 4754 1968 4792
rect 1922 4720 1928 4754
rect 1962 4720 1968 4754
rect 1922 4682 1968 4720
rect 1922 4648 1928 4682
rect 1962 4648 1968 4682
rect 1922 4625 1968 4648
rect 98 4358 1872 4367
rect 98 4233 1890 4358
rect -42440 -2298 -42408 2298
rect -40692 -2298 -40660 2298
rect -42440 -4409 -40660 -2298
rect 110 2298 1890 4233
rect 110 -2298 142 2298
rect 1858 -2298 1890 2298
rect 110 -4244 1890 -2298
rect -42531 -4410 -40660 -4409
rect -42531 -4543 -40757 -4410
rect 104 -4482 1980 -4244
rect -42531 -4760 -42485 -4543
rect -42531 -4794 -42525 -4760
rect -42491 -4794 -42485 -4760
rect -42531 -4832 -42485 -4794
rect -42531 -4866 -42525 -4832
rect -42491 -4866 -42485 -4832
rect -42531 -4904 -42485 -4866
rect -42531 -4938 -42525 -4904
rect -42491 -4938 -42485 -4904
rect -42531 -4976 -42485 -4938
rect -42531 -5010 -42525 -4976
rect -42491 -5010 -42485 -4976
rect -42531 -5048 -42485 -5010
rect -42531 -5082 -42525 -5048
rect -42491 -5082 -42485 -5048
rect -42531 -5120 -42485 -5082
rect -42531 -5154 -42525 -5120
rect -42491 -5154 -42485 -5120
rect -42531 -5192 -42485 -5154
rect -42531 -5226 -42525 -5192
rect -42491 -5226 -42485 -5192
rect -42531 -5264 -42485 -5226
rect -42531 -5298 -42525 -5264
rect -42491 -5298 -42485 -5264
rect -42531 -5336 -42485 -5298
rect -42531 -5370 -42525 -5336
rect -42491 -5370 -42485 -5336
rect -42531 -5408 -42485 -5370
rect -42531 -5442 -42525 -5408
rect -42491 -5442 -42485 -5408
rect -42531 -5480 -42485 -5442
rect -42531 -5514 -42525 -5480
rect -42491 -5514 -42485 -5480
rect -42531 -5537 -42485 -5514
rect -42435 -4760 -42389 -4737
rect -42435 -4794 -42429 -4760
rect -42395 -4794 -42389 -4760
rect -42435 -4832 -42389 -4794
rect -42435 -4866 -42429 -4832
rect -42395 -4866 -42389 -4832
rect -42435 -4904 -42389 -4866
rect -42435 -4938 -42429 -4904
rect -42395 -4938 -42389 -4904
rect -42435 -4976 -42389 -4938
rect -42435 -5010 -42429 -4976
rect -42395 -5010 -42389 -4976
rect -42435 -5048 -42389 -5010
rect -42435 -5082 -42429 -5048
rect -42395 -5082 -42389 -5048
rect -42435 -5120 -42389 -5082
rect -42435 -5154 -42429 -5120
rect -42395 -5154 -42389 -5120
rect -42435 -5192 -42389 -5154
rect -42435 -5226 -42429 -5192
rect -42395 -5226 -42389 -5192
rect -42435 -5264 -42389 -5226
rect -42435 -5298 -42429 -5264
rect -42395 -5298 -42389 -5264
rect -42435 -5336 -42389 -5298
rect -42435 -5370 -42429 -5336
rect -42395 -5370 -42389 -5336
rect -42435 -5408 -42389 -5370
rect -42435 -5442 -42429 -5408
rect -42395 -5442 -42389 -5408
rect -42435 -5480 -42389 -5442
rect -42435 -5514 -42429 -5480
rect -42395 -5514 -42389 -5480
rect -42435 -5800 -42389 -5514
rect -42339 -4760 -42293 -4543
rect -42339 -4794 -42333 -4760
rect -42299 -4794 -42293 -4760
rect -42339 -4832 -42293 -4794
rect -42339 -4866 -42333 -4832
rect -42299 -4866 -42293 -4832
rect -42339 -4904 -42293 -4866
rect -42339 -4938 -42333 -4904
rect -42299 -4938 -42293 -4904
rect -42339 -4976 -42293 -4938
rect -42339 -5010 -42333 -4976
rect -42299 -5010 -42293 -4976
rect -42339 -5048 -42293 -5010
rect -42339 -5082 -42333 -5048
rect -42299 -5082 -42293 -5048
rect -42339 -5120 -42293 -5082
rect -42339 -5154 -42333 -5120
rect -42299 -5154 -42293 -5120
rect -42339 -5192 -42293 -5154
rect -42339 -5226 -42333 -5192
rect -42299 -5226 -42293 -5192
rect -42339 -5264 -42293 -5226
rect -42339 -5298 -42333 -5264
rect -42299 -5298 -42293 -5264
rect -42339 -5336 -42293 -5298
rect -42339 -5370 -42333 -5336
rect -42299 -5370 -42293 -5336
rect -42339 -5408 -42293 -5370
rect -42339 -5442 -42333 -5408
rect -42299 -5442 -42293 -5408
rect -42339 -5480 -42293 -5442
rect -42339 -5514 -42333 -5480
rect -42299 -5514 -42293 -5480
rect -42339 -5537 -42293 -5514
rect -42243 -4760 -42197 -4737
rect -42243 -4794 -42237 -4760
rect -42203 -4794 -42197 -4760
rect -42243 -4832 -42197 -4794
rect -42243 -4866 -42237 -4832
rect -42203 -4866 -42197 -4832
rect -42243 -4904 -42197 -4866
rect -42243 -4938 -42237 -4904
rect -42203 -4938 -42197 -4904
rect -42243 -4976 -42197 -4938
rect -42243 -5010 -42237 -4976
rect -42203 -5010 -42197 -4976
rect -42243 -5048 -42197 -5010
rect -42243 -5082 -42237 -5048
rect -42203 -5082 -42197 -5048
rect -42243 -5120 -42197 -5082
rect -42243 -5154 -42237 -5120
rect -42203 -5154 -42197 -5120
rect -42243 -5192 -42197 -5154
rect -42243 -5226 -42237 -5192
rect -42203 -5226 -42197 -5192
rect -42243 -5264 -42197 -5226
rect -42243 -5298 -42237 -5264
rect -42203 -5298 -42197 -5264
rect -42243 -5336 -42197 -5298
rect -42243 -5370 -42237 -5336
rect -42203 -5370 -42197 -5336
rect -42243 -5408 -42197 -5370
rect -42243 -5442 -42237 -5408
rect -42203 -5442 -42197 -5408
rect -42243 -5480 -42197 -5442
rect -42243 -5514 -42237 -5480
rect -42203 -5514 -42197 -5480
rect -42243 -5800 -42197 -5514
rect -42147 -4760 -42101 -4543
rect -42147 -4794 -42141 -4760
rect -42107 -4794 -42101 -4760
rect -42147 -4832 -42101 -4794
rect -42147 -4866 -42141 -4832
rect -42107 -4866 -42101 -4832
rect -42147 -4904 -42101 -4866
rect -42147 -4938 -42141 -4904
rect -42107 -4938 -42101 -4904
rect -42147 -4976 -42101 -4938
rect -42147 -5010 -42141 -4976
rect -42107 -5010 -42101 -4976
rect -42147 -5048 -42101 -5010
rect -42147 -5082 -42141 -5048
rect -42107 -5082 -42101 -5048
rect -42147 -5120 -42101 -5082
rect -42147 -5154 -42141 -5120
rect -42107 -5154 -42101 -5120
rect -42147 -5192 -42101 -5154
rect -42147 -5226 -42141 -5192
rect -42107 -5226 -42101 -5192
rect -42147 -5264 -42101 -5226
rect -42147 -5298 -42141 -5264
rect -42107 -5298 -42101 -5264
rect -42147 -5336 -42101 -5298
rect -42147 -5370 -42141 -5336
rect -42107 -5370 -42101 -5336
rect -42147 -5408 -42101 -5370
rect -42147 -5442 -42141 -5408
rect -42107 -5442 -42101 -5408
rect -42147 -5480 -42101 -5442
rect -42147 -5514 -42141 -5480
rect -42107 -5514 -42101 -5480
rect -42147 -5537 -42101 -5514
rect -42051 -4760 -42005 -4737
rect -42051 -4794 -42045 -4760
rect -42011 -4794 -42005 -4760
rect -42051 -4832 -42005 -4794
rect -42051 -4866 -42045 -4832
rect -42011 -4866 -42005 -4832
rect -42051 -4904 -42005 -4866
rect -42051 -4938 -42045 -4904
rect -42011 -4938 -42005 -4904
rect -42051 -4976 -42005 -4938
rect -42051 -5010 -42045 -4976
rect -42011 -5010 -42005 -4976
rect -42051 -5048 -42005 -5010
rect -42051 -5082 -42045 -5048
rect -42011 -5082 -42005 -5048
rect -42051 -5120 -42005 -5082
rect -42051 -5154 -42045 -5120
rect -42011 -5154 -42005 -5120
rect -42051 -5192 -42005 -5154
rect -42051 -5226 -42045 -5192
rect -42011 -5226 -42005 -5192
rect -42051 -5264 -42005 -5226
rect -42051 -5298 -42045 -5264
rect -42011 -5298 -42005 -5264
rect -42051 -5336 -42005 -5298
rect -42051 -5370 -42045 -5336
rect -42011 -5370 -42005 -5336
rect -42051 -5408 -42005 -5370
rect -42051 -5442 -42045 -5408
rect -42011 -5442 -42005 -5408
rect -42051 -5480 -42005 -5442
rect -42051 -5514 -42045 -5480
rect -42011 -5514 -42005 -5480
rect -42051 -5800 -42005 -5514
rect -41955 -4760 -41909 -4543
rect -41955 -4794 -41949 -4760
rect -41915 -4794 -41909 -4760
rect -41955 -4832 -41909 -4794
rect -41955 -4866 -41949 -4832
rect -41915 -4866 -41909 -4832
rect -41955 -4904 -41909 -4866
rect -41955 -4938 -41949 -4904
rect -41915 -4938 -41909 -4904
rect -41955 -4976 -41909 -4938
rect -41955 -5010 -41949 -4976
rect -41915 -5010 -41909 -4976
rect -41955 -5048 -41909 -5010
rect -41955 -5082 -41949 -5048
rect -41915 -5082 -41909 -5048
rect -41955 -5120 -41909 -5082
rect -41955 -5154 -41949 -5120
rect -41915 -5154 -41909 -5120
rect -41955 -5192 -41909 -5154
rect -41955 -5226 -41949 -5192
rect -41915 -5226 -41909 -5192
rect -41955 -5264 -41909 -5226
rect -41955 -5298 -41949 -5264
rect -41915 -5298 -41909 -5264
rect -41955 -5336 -41909 -5298
rect -41955 -5370 -41949 -5336
rect -41915 -5370 -41909 -5336
rect -41955 -5408 -41909 -5370
rect -41955 -5442 -41949 -5408
rect -41915 -5442 -41909 -5408
rect -41955 -5480 -41909 -5442
rect -41955 -5514 -41949 -5480
rect -41915 -5514 -41909 -5480
rect -41955 -5537 -41909 -5514
rect -41859 -4760 -41813 -4737
rect -41859 -4794 -41853 -4760
rect -41819 -4794 -41813 -4760
rect -41859 -4832 -41813 -4794
rect -41859 -4866 -41853 -4832
rect -41819 -4866 -41813 -4832
rect -41859 -4904 -41813 -4866
rect -41859 -4938 -41853 -4904
rect -41819 -4938 -41813 -4904
rect -41859 -4976 -41813 -4938
rect -41859 -5010 -41853 -4976
rect -41819 -5010 -41813 -4976
rect -41859 -5048 -41813 -5010
rect -41859 -5082 -41853 -5048
rect -41819 -5082 -41813 -5048
rect -41859 -5120 -41813 -5082
rect -41859 -5154 -41853 -5120
rect -41819 -5154 -41813 -5120
rect -41859 -5192 -41813 -5154
rect -41859 -5226 -41853 -5192
rect -41819 -5226 -41813 -5192
rect -41859 -5264 -41813 -5226
rect -41859 -5298 -41853 -5264
rect -41819 -5298 -41813 -5264
rect -41859 -5336 -41813 -5298
rect -41859 -5370 -41853 -5336
rect -41819 -5370 -41813 -5336
rect -41859 -5408 -41813 -5370
rect -41859 -5442 -41853 -5408
rect -41819 -5442 -41813 -5408
rect -41859 -5480 -41813 -5442
rect -41859 -5514 -41853 -5480
rect -41819 -5514 -41813 -5480
rect -41859 -5800 -41813 -5514
rect -41763 -4760 -41717 -4543
rect -41763 -4794 -41757 -4760
rect -41723 -4794 -41717 -4760
rect -41763 -4832 -41717 -4794
rect -41763 -4866 -41757 -4832
rect -41723 -4866 -41717 -4832
rect -41763 -4904 -41717 -4866
rect -41763 -4938 -41757 -4904
rect -41723 -4938 -41717 -4904
rect -41763 -4976 -41717 -4938
rect -41763 -5010 -41757 -4976
rect -41723 -5010 -41717 -4976
rect -41763 -5048 -41717 -5010
rect -41763 -5082 -41757 -5048
rect -41723 -5082 -41717 -5048
rect -41763 -5120 -41717 -5082
rect -41763 -5154 -41757 -5120
rect -41723 -5154 -41717 -5120
rect -41763 -5192 -41717 -5154
rect -41763 -5226 -41757 -5192
rect -41723 -5226 -41717 -5192
rect -41763 -5264 -41717 -5226
rect -41763 -5298 -41757 -5264
rect -41723 -5298 -41717 -5264
rect -41763 -5336 -41717 -5298
rect -41763 -5370 -41757 -5336
rect -41723 -5370 -41717 -5336
rect -41763 -5408 -41717 -5370
rect -41763 -5442 -41757 -5408
rect -41723 -5442 -41717 -5408
rect -41763 -5480 -41717 -5442
rect -41763 -5514 -41757 -5480
rect -41723 -5514 -41717 -5480
rect -41763 -5537 -41717 -5514
rect -41667 -4760 -41621 -4737
rect -41667 -4794 -41661 -4760
rect -41627 -4794 -41621 -4760
rect -41667 -4832 -41621 -4794
rect -41667 -4866 -41661 -4832
rect -41627 -4866 -41621 -4832
rect -41667 -4904 -41621 -4866
rect -41667 -4938 -41661 -4904
rect -41627 -4938 -41621 -4904
rect -41667 -4976 -41621 -4938
rect -41667 -5010 -41661 -4976
rect -41627 -5010 -41621 -4976
rect -41667 -5048 -41621 -5010
rect -41667 -5082 -41661 -5048
rect -41627 -5082 -41621 -5048
rect -41667 -5120 -41621 -5082
rect -41667 -5154 -41661 -5120
rect -41627 -5154 -41621 -5120
rect -41667 -5192 -41621 -5154
rect -41667 -5226 -41661 -5192
rect -41627 -5226 -41621 -5192
rect -41667 -5264 -41621 -5226
rect -41667 -5298 -41661 -5264
rect -41627 -5298 -41621 -5264
rect -41667 -5336 -41621 -5298
rect -41667 -5370 -41661 -5336
rect -41627 -5370 -41621 -5336
rect -41667 -5408 -41621 -5370
rect -41667 -5442 -41661 -5408
rect -41627 -5442 -41621 -5408
rect -41667 -5480 -41621 -5442
rect -41667 -5514 -41661 -5480
rect -41627 -5514 -41621 -5480
rect -41667 -5800 -41621 -5514
rect -41571 -4760 -41525 -4543
rect -41571 -4794 -41565 -4760
rect -41531 -4794 -41525 -4760
rect -41571 -4832 -41525 -4794
rect -41571 -4866 -41565 -4832
rect -41531 -4866 -41525 -4832
rect -41571 -4904 -41525 -4866
rect -41571 -4938 -41565 -4904
rect -41531 -4938 -41525 -4904
rect -41571 -4976 -41525 -4938
rect -41571 -5010 -41565 -4976
rect -41531 -5010 -41525 -4976
rect -41571 -5048 -41525 -5010
rect -41571 -5082 -41565 -5048
rect -41531 -5082 -41525 -5048
rect -41571 -5120 -41525 -5082
rect -41571 -5154 -41565 -5120
rect -41531 -5154 -41525 -5120
rect -41571 -5192 -41525 -5154
rect -41571 -5226 -41565 -5192
rect -41531 -5226 -41525 -5192
rect -41571 -5264 -41525 -5226
rect -41571 -5298 -41565 -5264
rect -41531 -5298 -41525 -5264
rect -41571 -5336 -41525 -5298
rect -41571 -5370 -41565 -5336
rect -41531 -5370 -41525 -5336
rect -41571 -5408 -41525 -5370
rect -41571 -5442 -41565 -5408
rect -41531 -5442 -41525 -5408
rect -41571 -5480 -41525 -5442
rect -41571 -5514 -41565 -5480
rect -41531 -5514 -41525 -5480
rect -41571 -5537 -41525 -5514
rect -41475 -4760 -41429 -4737
rect -41475 -4794 -41469 -4760
rect -41435 -4794 -41429 -4760
rect -41475 -4832 -41429 -4794
rect -41475 -4866 -41469 -4832
rect -41435 -4866 -41429 -4832
rect -41475 -4904 -41429 -4866
rect -41475 -4938 -41469 -4904
rect -41435 -4938 -41429 -4904
rect -41475 -4976 -41429 -4938
rect -41475 -5010 -41469 -4976
rect -41435 -5010 -41429 -4976
rect -41475 -5048 -41429 -5010
rect -41475 -5082 -41469 -5048
rect -41435 -5082 -41429 -5048
rect -41475 -5120 -41429 -5082
rect -41475 -5154 -41469 -5120
rect -41435 -5154 -41429 -5120
rect -41475 -5192 -41429 -5154
rect -41475 -5226 -41469 -5192
rect -41435 -5226 -41429 -5192
rect -41475 -5264 -41429 -5226
rect -41475 -5298 -41469 -5264
rect -41435 -5298 -41429 -5264
rect -41475 -5336 -41429 -5298
rect -41475 -5370 -41469 -5336
rect -41435 -5370 -41429 -5336
rect -41475 -5408 -41429 -5370
rect -41475 -5442 -41469 -5408
rect -41435 -5442 -41429 -5408
rect -41475 -5480 -41429 -5442
rect -41475 -5514 -41469 -5480
rect -41435 -5514 -41429 -5480
rect -41475 -5800 -41429 -5514
rect -41379 -4760 -41333 -4543
rect -41379 -4794 -41373 -4760
rect -41339 -4794 -41333 -4760
rect -41379 -4832 -41333 -4794
rect -41379 -4866 -41373 -4832
rect -41339 -4866 -41333 -4832
rect -41379 -4904 -41333 -4866
rect -41379 -4938 -41373 -4904
rect -41339 -4938 -41333 -4904
rect -41379 -4976 -41333 -4938
rect -41379 -5010 -41373 -4976
rect -41339 -5010 -41333 -4976
rect -41379 -5048 -41333 -5010
rect -41379 -5082 -41373 -5048
rect -41339 -5082 -41333 -5048
rect -41379 -5120 -41333 -5082
rect -41379 -5154 -41373 -5120
rect -41339 -5154 -41333 -5120
rect -41379 -5192 -41333 -5154
rect -41379 -5226 -41373 -5192
rect -41339 -5226 -41333 -5192
rect -41379 -5264 -41333 -5226
rect -41379 -5298 -41373 -5264
rect -41339 -5298 -41333 -5264
rect -41379 -5336 -41333 -5298
rect -41379 -5370 -41373 -5336
rect -41339 -5370 -41333 -5336
rect -41379 -5408 -41333 -5370
rect -41379 -5442 -41373 -5408
rect -41339 -5442 -41333 -5408
rect -41379 -5480 -41333 -5442
rect -41379 -5514 -41373 -5480
rect -41339 -5514 -41333 -5480
rect -41379 -5537 -41333 -5514
rect -41283 -4760 -41237 -4737
rect -41283 -4794 -41277 -4760
rect -41243 -4794 -41237 -4760
rect -41283 -4832 -41237 -4794
rect -41283 -4866 -41277 -4832
rect -41243 -4866 -41237 -4832
rect -41283 -4904 -41237 -4866
rect -41283 -4938 -41277 -4904
rect -41243 -4938 -41237 -4904
rect -41283 -4976 -41237 -4938
rect -41283 -5010 -41277 -4976
rect -41243 -5010 -41237 -4976
rect -41283 -5048 -41237 -5010
rect -41283 -5082 -41277 -5048
rect -41243 -5082 -41237 -5048
rect -41283 -5120 -41237 -5082
rect -41283 -5154 -41277 -5120
rect -41243 -5154 -41237 -5120
rect -41283 -5192 -41237 -5154
rect -41283 -5226 -41277 -5192
rect -41243 -5226 -41237 -5192
rect -41283 -5264 -41237 -5226
rect -41283 -5298 -41277 -5264
rect -41243 -5298 -41237 -5264
rect -41283 -5336 -41237 -5298
rect -41283 -5370 -41277 -5336
rect -41243 -5370 -41237 -5336
rect -41283 -5408 -41237 -5370
rect -41283 -5442 -41277 -5408
rect -41243 -5442 -41237 -5408
rect -41283 -5480 -41237 -5442
rect -41283 -5514 -41277 -5480
rect -41243 -5514 -41237 -5480
rect -41283 -5800 -41237 -5514
rect -41187 -4760 -41141 -4543
rect -41187 -4794 -41181 -4760
rect -41147 -4794 -41141 -4760
rect -41187 -4832 -41141 -4794
rect -41187 -4866 -41181 -4832
rect -41147 -4866 -41141 -4832
rect -41187 -4904 -41141 -4866
rect -41187 -4938 -41181 -4904
rect -41147 -4938 -41141 -4904
rect -41187 -4976 -41141 -4938
rect -41187 -5010 -41181 -4976
rect -41147 -5010 -41141 -4976
rect -41187 -5048 -41141 -5010
rect -41187 -5082 -41181 -5048
rect -41147 -5082 -41141 -5048
rect -41187 -5120 -41141 -5082
rect -41187 -5154 -41181 -5120
rect -41147 -5154 -41141 -5120
rect -41187 -5192 -41141 -5154
rect -41187 -5226 -41181 -5192
rect -41147 -5226 -41141 -5192
rect -41187 -5264 -41141 -5226
rect -41187 -5298 -41181 -5264
rect -41147 -5298 -41141 -5264
rect -41187 -5336 -41141 -5298
rect -41187 -5370 -41181 -5336
rect -41147 -5370 -41141 -5336
rect -41187 -5408 -41141 -5370
rect -41187 -5442 -41181 -5408
rect -41147 -5442 -41141 -5408
rect -41187 -5480 -41141 -5442
rect -41187 -5514 -41181 -5480
rect -41147 -5514 -41141 -5480
rect -41187 -5537 -41141 -5514
rect -41091 -4760 -41045 -4737
rect -41091 -4794 -41085 -4760
rect -41051 -4794 -41045 -4760
rect -41091 -4832 -41045 -4794
rect -41091 -4866 -41085 -4832
rect -41051 -4866 -41045 -4832
rect -41091 -4904 -41045 -4866
rect -41091 -4938 -41085 -4904
rect -41051 -4938 -41045 -4904
rect -41091 -4976 -41045 -4938
rect -41091 -5010 -41085 -4976
rect -41051 -5010 -41045 -4976
rect -41091 -5048 -41045 -5010
rect -41091 -5082 -41085 -5048
rect -41051 -5082 -41045 -5048
rect -41091 -5120 -41045 -5082
rect -41091 -5154 -41085 -5120
rect -41051 -5154 -41045 -5120
rect -41091 -5192 -41045 -5154
rect -41091 -5226 -41085 -5192
rect -41051 -5226 -41045 -5192
rect -41091 -5264 -41045 -5226
rect -41091 -5298 -41085 -5264
rect -41051 -5298 -41045 -5264
rect -41091 -5336 -41045 -5298
rect -41091 -5370 -41085 -5336
rect -41051 -5370 -41045 -5336
rect -41091 -5408 -41045 -5370
rect -41091 -5442 -41085 -5408
rect -41051 -5442 -41045 -5408
rect -41091 -5480 -41045 -5442
rect -41091 -5514 -41085 -5480
rect -41051 -5514 -41045 -5480
rect -41091 -5800 -41045 -5514
rect -40995 -4760 -40949 -4543
rect -40995 -4794 -40989 -4760
rect -40955 -4794 -40949 -4760
rect -40995 -4832 -40949 -4794
rect -40995 -4866 -40989 -4832
rect -40955 -4866 -40949 -4832
rect -40995 -4904 -40949 -4866
rect -40995 -4938 -40989 -4904
rect -40955 -4938 -40949 -4904
rect -40995 -4976 -40949 -4938
rect -40995 -5010 -40989 -4976
rect -40955 -5010 -40949 -4976
rect -40995 -5048 -40949 -5010
rect -40995 -5082 -40989 -5048
rect -40955 -5082 -40949 -5048
rect -40995 -5120 -40949 -5082
rect -40995 -5154 -40989 -5120
rect -40955 -5154 -40949 -5120
rect -40995 -5192 -40949 -5154
rect -40995 -5226 -40989 -5192
rect -40955 -5226 -40949 -5192
rect -40995 -5264 -40949 -5226
rect -40995 -5298 -40989 -5264
rect -40955 -5298 -40949 -5264
rect -40995 -5336 -40949 -5298
rect -40995 -5370 -40989 -5336
rect -40955 -5370 -40949 -5336
rect -40995 -5408 -40949 -5370
rect -40995 -5442 -40989 -5408
rect -40955 -5442 -40949 -5408
rect -40995 -5480 -40949 -5442
rect -40995 -5514 -40989 -5480
rect -40955 -5514 -40949 -5480
rect -40995 -5537 -40949 -5514
rect -40899 -4760 -40853 -4737
rect -40899 -4794 -40893 -4760
rect -40859 -4794 -40853 -4760
rect -40899 -4832 -40853 -4794
rect -40899 -4866 -40893 -4832
rect -40859 -4866 -40853 -4832
rect -40899 -4904 -40853 -4866
rect -40899 -4938 -40893 -4904
rect -40859 -4938 -40853 -4904
rect -40899 -4976 -40853 -4938
rect -40899 -5010 -40893 -4976
rect -40859 -5010 -40853 -4976
rect -40899 -5048 -40853 -5010
rect -40899 -5082 -40893 -5048
rect -40859 -5082 -40853 -5048
rect -40899 -5120 -40853 -5082
rect -40899 -5154 -40893 -5120
rect -40859 -5154 -40853 -5120
rect -40899 -5192 -40853 -5154
rect -40899 -5226 -40893 -5192
rect -40859 -5226 -40853 -5192
rect -40899 -5264 -40853 -5226
rect -40899 -5298 -40893 -5264
rect -40859 -5298 -40853 -5264
rect -40899 -5336 -40853 -5298
rect -40899 -5370 -40893 -5336
rect -40859 -5370 -40853 -5336
rect -40899 -5408 -40853 -5370
rect -40899 -5442 -40893 -5408
rect -40859 -5442 -40853 -5408
rect -40899 -5480 -40853 -5442
rect -40899 -5514 -40893 -5480
rect -40859 -5514 -40853 -5480
rect -40899 -5800 -40853 -5514
rect -40803 -4760 -40757 -4543
rect 206 -4569 1980 -4482
rect -40803 -4794 -40797 -4760
rect -40763 -4794 -40757 -4760
rect -40803 -4832 -40757 -4794
rect -40803 -4866 -40797 -4832
rect -40763 -4866 -40757 -4832
rect -40803 -4904 -40757 -4866
rect -40803 -4938 -40797 -4904
rect -40763 -4938 -40757 -4904
rect -40803 -4976 -40757 -4938
rect -40803 -5010 -40797 -4976
rect -40763 -5010 -40757 -4976
rect -40803 -5048 -40757 -5010
rect -40803 -5082 -40797 -5048
rect -40763 -5082 -40757 -5048
rect -40803 -5120 -40757 -5082
rect -40803 -5154 -40797 -5120
rect -40763 -5154 -40757 -5120
rect -40803 -5192 -40757 -5154
rect -40803 -5226 -40797 -5192
rect -40763 -5226 -40757 -5192
rect -40803 -5264 -40757 -5226
rect -40803 -5298 -40797 -5264
rect -40763 -5298 -40757 -5264
rect -40803 -5336 -40757 -5298
rect -40803 -5370 -40797 -5336
rect -40763 -5370 -40757 -5336
rect -40803 -5408 -40757 -5370
rect -40803 -5442 -40797 -5408
rect -40763 -5442 -40757 -5408
rect -40803 -5480 -40757 -5442
rect -40803 -5514 -40797 -5480
rect -40763 -5514 -40757 -5480
rect -40803 -5537 -40757 -5514
rect -40707 -4760 -40661 -4737
rect -40707 -4794 -40701 -4760
rect -40667 -4794 -40661 -4760
rect -40707 -4832 -40661 -4794
rect -40707 -4866 -40701 -4832
rect -40667 -4866 -40661 -4832
rect -40707 -4904 -40661 -4866
rect -40707 -4938 -40701 -4904
rect -40667 -4938 -40661 -4904
rect -40707 -4976 -40661 -4938
rect -40707 -5010 -40701 -4976
rect -40667 -5010 -40661 -4976
rect -40707 -5048 -40661 -5010
rect -40707 -5082 -40701 -5048
rect -40667 -5082 -40661 -5048
rect -40707 -5120 -40661 -5082
rect -40707 -5154 -40701 -5120
rect -40667 -5154 -40661 -5120
rect -40707 -5192 -40661 -5154
rect -40707 -5226 -40701 -5192
rect -40667 -5226 -40661 -5192
rect -40707 -5264 -40661 -5226
rect -40707 -5298 -40701 -5264
rect -40667 -5298 -40661 -5264
rect -40707 -5336 -40661 -5298
rect -40707 -5370 -40701 -5336
rect -40667 -5370 -40661 -5336
rect -40707 -5408 -40661 -5370
rect -40707 -5442 -40701 -5408
rect -40667 -5442 -40661 -5408
rect -40707 -5480 -40661 -5442
rect -40707 -5514 -40701 -5480
rect -40667 -5514 -40661 -5480
rect -40707 -5800 -40661 -5514
rect -42435 -5934 -40661 -5800
rect 110 -4786 156 -4744
rect 110 -4820 116 -4786
rect 150 -4820 156 -4786
rect 110 -4858 156 -4820
rect 110 -4892 116 -4858
rect 150 -4892 156 -4858
rect 110 -4930 156 -4892
rect 110 -4964 116 -4930
rect 150 -4964 156 -4930
rect 110 -5002 156 -4964
rect 110 -5036 116 -5002
rect 150 -5036 156 -5002
rect 110 -5074 156 -5036
rect 110 -5108 116 -5074
rect 150 -5108 156 -5074
rect 110 -5146 156 -5108
rect 110 -5180 116 -5146
rect 150 -5180 156 -5146
rect 110 -5218 156 -5180
rect 110 -5252 116 -5218
rect 150 -5252 156 -5218
rect 110 -5290 156 -5252
rect 110 -5324 116 -5290
rect 150 -5324 156 -5290
rect 110 -5362 156 -5324
rect 110 -5396 116 -5362
rect 150 -5396 156 -5362
rect 110 -5434 156 -5396
rect 110 -5468 116 -5434
rect 150 -5468 156 -5434
rect 110 -5506 156 -5468
rect 110 -5540 116 -5506
rect 150 -5540 156 -5506
rect 110 -5790 156 -5540
rect 206 -4786 252 -4569
rect 206 -4820 212 -4786
rect 246 -4820 252 -4786
rect 206 -4858 252 -4820
rect 206 -4892 212 -4858
rect 246 -4892 252 -4858
rect 206 -4930 252 -4892
rect 206 -4964 212 -4930
rect 246 -4964 252 -4930
rect 206 -5002 252 -4964
rect 206 -5036 212 -5002
rect 246 -5036 252 -5002
rect 206 -5074 252 -5036
rect 206 -5108 212 -5074
rect 246 -5108 252 -5074
rect 206 -5146 252 -5108
rect 206 -5180 212 -5146
rect 246 -5180 252 -5146
rect 206 -5218 252 -5180
rect 206 -5252 212 -5218
rect 246 -5252 252 -5218
rect 206 -5290 252 -5252
rect 206 -5324 212 -5290
rect 246 -5324 252 -5290
rect 206 -5362 252 -5324
rect 206 -5396 212 -5362
rect 246 -5396 252 -5362
rect 206 -5434 252 -5396
rect 206 -5468 212 -5434
rect 246 -5468 252 -5434
rect 206 -5506 252 -5468
rect 206 -5540 212 -5506
rect 246 -5540 252 -5506
rect 206 -5563 252 -5540
rect 302 -4786 348 -4744
rect 302 -4820 308 -4786
rect 342 -4820 348 -4786
rect 302 -4858 348 -4820
rect 302 -4892 308 -4858
rect 342 -4892 348 -4858
rect 302 -4930 348 -4892
rect 302 -4964 308 -4930
rect 342 -4964 348 -4930
rect 302 -5002 348 -4964
rect 302 -5036 308 -5002
rect 342 -5036 348 -5002
rect 302 -5074 348 -5036
rect 302 -5108 308 -5074
rect 342 -5108 348 -5074
rect 302 -5146 348 -5108
rect 302 -5180 308 -5146
rect 342 -5180 348 -5146
rect 302 -5218 348 -5180
rect 302 -5252 308 -5218
rect 342 -5252 348 -5218
rect 302 -5290 348 -5252
rect 302 -5324 308 -5290
rect 342 -5324 348 -5290
rect 302 -5362 348 -5324
rect 302 -5396 308 -5362
rect 342 -5396 348 -5362
rect 302 -5434 348 -5396
rect 302 -5468 308 -5434
rect 342 -5468 348 -5434
rect 302 -5506 348 -5468
rect 302 -5540 308 -5506
rect 342 -5540 348 -5506
rect 302 -5790 348 -5540
rect 398 -4786 444 -4569
rect 398 -4820 404 -4786
rect 438 -4820 444 -4786
rect 398 -4858 444 -4820
rect 398 -4892 404 -4858
rect 438 -4892 444 -4858
rect 398 -4930 444 -4892
rect 398 -4964 404 -4930
rect 438 -4964 444 -4930
rect 398 -5002 444 -4964
rect 398 -5036 404 -5002
rect 438 -5036 444 -5002
rect 398 -5074 444 -5036
rect 398 -5108 404 -5074
rect 438 -5108 444 -5074
rect 398 -5146 444 -5108
rect 398 -5180 404 -5146
rect 438 -5180 444 -5146
rect 398 -5218 444 -5180
rect 398 -5252 404 -5218
rect 438 -5252 444 -5218
rect 398 -5290 444 -5252
rect 398 -5324 404 -5290
rect 438 -5324 444 -5290
rect 398 -5362 444 -5324
rect 398 -5396 404 -5362
rect 438 -5396 444 -5362
rect 398 -5434 444 -5396
rect 398 -5468 404 -5434
rect 438 -5468 444 -5434
rect 398 -5506 444 -5468
rect 398 -5540 404 -5506
rect 438 -5540 444 -5506
rect 398 -5563 444 -5540
rect 494 -4786 540 -4744
rect 494 -4820 500 -4786
rect 534 -4820 540 -4786
rect 494 -4858 540 -4820
rect 494 -4892 500 -4858
rect 534 -4892 540 -4858
rect 494 -4930 540 -4892
rect 494 -4964 500 -4930
rect 534 -4964 540 -4930
rect 494 -5002 540 -4964
rect 494 -5036 500 -5002
rect 534 -5036 540 -5002
rect 494 -5074 540 -5036
rect 494 -5108 500 -5074
rect 534 -5108 540 -5074
rect 494 -5146 540 -5108
rect 494 -5180 500 -5146
rect 534 -5180 540 -5146
rect 494 -5218 540 -5180
rect 494 -5252 500 -5218
rect 534 -5252 540 -5218
rect 494 -5290 540 -5252
rect 494 -5324 500 -5290
rect 534 -5324 540 -5290
rect 494 -5362 540 -5324
rect 494 -5396 500 -5362
rect 534 -5396 540 -5362
rect 494 -5434 540 -5396
rect 494 -5468 500 -5434
rect 534 -5468 540 -5434
rect 494 -5506 540 -5468
rect 494 -5540 500 -5506
rect 534 -5540 540 -5506
rect 494 -5790 540 -5540
rect 590 -4786 636 -4569
rect 590 -4820 596 -4786
rect 630 -4820 636 -4786
rect 590 -4858 636 -4820
rect 590 -4892 596 -4858
rect 630 -4892 636 -4858
rect 590 -4930 636 -4892
rect 590 -4964 596 -4930
rect 630 -4964 636 -4930
rect 590 -5002 636 -4964
rect 590 -5036 596 -5002
rect 630 -5036 636 -5002
rect 590 -5074 636 -5036
rect 590 -5108 596 -5074
rect 630 -5108 636 -5074
rect 590 -5146 636 -5108
rect 590 -5180 596 -5146
rect 630 -5180 636 -5146
rect 590 -5218 636 -5180
rect 590 -5252 596 -5218
rect 630 -5252 636 -5218
rect 590 -5290 636 -5252
rect 590 -5324 596 -5290
rect 630 -5324 636 -5290
rect 590 -5362 636 -5324
rect 590 -5396 596 -5362
rect 630 -5396 636 -5362
rect 590 -5434 636 -5396
rect 590 -5468 596 -5434
rect 630 -5468 636 -5434
rect 590 -5506 636 -5468
rect 590 -5540 596 -5506
rect 630 -5540 636 -5506
rect 590 -5563 636 -5540
rect 686 -4786 732 -4744
rect 686 -4820 692 -4786
rect 726 -4820 732 -4786
rect 686 -4858 732 -4820
rect 686 -4892 692 -4858
rect 726 -4892 732 -4858
rect 686 -4930 732 -4892
rect 686 -4964 692 -4930
rect 726 -4964 732 -4930
rect 686 -5002 732 -4964
rect 686 -5036 692 -5002
rect 726 -5036 732 -5002
rect 686 -5074 732 -5036
rect 686 -5108 692 -5074
rect 726 -5108 732 -5074
rect 686 -5146 732 -5108
rect 686 -5180 692 -5146
rect 726 -5180 732 -5146
rect 686 -5218 732 -5180
rect 686 -5252 692 -5218
rect 726 -5252 732 -5218
rect 686 -5290 732 -5252
rect 686 -5324 692 -5290
rect 726 -5324 732 -5290
rect 686 -5362 732 -5324
rect 686 -5396 692 -5362
rect 726 -5396 732 -5362
rect 686 -5434 732 -5396
rect 686 -5468 692 -5434
rect 726 -5468 732 -5434
rect 686 -5506 732 -5468
rect 686 -5540 692 -5506
rect 726 -5540 732 -5506
rect 686 -5790 732 -5540
rect 782 -4786 828 -4569
rect 782 -4820 788 -4786
rect 822 -4820 828 -4786
rect 782 -4858 828 -4820
rect 782 -4892 788 -4858
rect 822 -4892 828 -4858
rect 782 -4930 828 -4892
rect 782 -4964 788 -4930
rect 822 -4964 828 -4930
rect 782 -5002 828 -4964
rect 782 -5036 788 -5002
rect 822 -5036 828 -5002
rect 782 -5074 828 -5036
rect 782 -5108 788 -5074
rect 822 -5108 828 -5074
rect 782 -5146 828 -5108
rect 782 -5180 788 -5146
rect 822 -5180 828 -5146
rect 782 -5218 828 -5180
rect 782 -5252 788 -5218
rect 822 -5252 828 -5218
rect 782 -5290 828 -5252
rect 782 -5324 788 -5290
rect 822 -5324 828 -5290
rect 782 -5362 828 -5324
rect 782 -5396 788 -5362
rect 822 -5396 828 -5362
rect 782 -5434 828 -5396
rect 782 -5468 788 -5434
rect 822 -5468 828 -5434
rect 782 -5506 828 -5468
rect 782 -5540 788 -5506
rect 822 -5540 828 -5506
rect 782 -5563 828 -5540
rect 878 -4786 924 -4744
rect 878 -4820 884 -4786
rect 918 -4820 924 -4786
rect 878 -4858 924 -4820
rect 878 -4892 884 -4858
rect 918 -4892 924 -4858
rect 878 -4930 924 -4892
rect 878 -4964 884 -4930
rect 918 -4964 924 -4930
rect 878 -5002 924 -4964
rect 878 -5036 884 -5002
rect 918 -5036 924 -5002
rect 878 -5074 924 -5036
rect 878 -5108 884 -5074
rect 918 -5108 924 -5074
rect 878 -5146 924 -5108
rect 878 -5180 884 -5146
rect 918 -5180 924 -5146
rect 878 -5218 924 -5180
rect 878 -5252 884 -5218
rect 918 -5252 924 -5218
rect 878 -5290 924 -5252
rect 878 -5324 884 -5290
rect 918 -5324 924 -5290
rect 878 -5362 924 -5324
rect 878 -5396 884 -5362
rect 918 -5396 924 -5362
rect 878 -5434 924 -5396
rect 878 -5468 884 -5434
rect 918 -5468 924 -5434
rect 878 -5506 924 -5468
rect 878 -5540 884 -5506
rect 918 -5540 924 -5506
rect 878 -5790 924 -5540
rect 974 -4786 1020 -4569
rect 974 -4820 980 -4786
rect 1014 -4820 1020 -4786
rect 974 -4858 1020 -4820
rect 974 -4892 980 -4858
rect 1014 -4892 1020 -4858
rect 974 -4930 1020 -4892
rect 974 -4964 980 -4930
rect 1014 -4964 1020 -4930
rect 974 -5002 1020 -4964
rect 974 -5036 980 -5002
rect 1014 -5036 1020 -5002
rect 974 -5074 1020 -5036
rect 974 -5108 980 -5074
rect 1014 -5108 1020 -5074
rect 974 -5146 1020 -5108
rect 974 -5180 980 -5146
rect 1014 -5180 1020 -5146
rect 974 -5218 1020 -5180
rect 974 -5252 980 -5218
rect 1014 -5252 1020 -5218
rect 974 -5290 1020 -5252
rect 974 -5324 980 -5290
rect 1014 -5324 1020 -5290
rect 974 -5362 1020 -5324
rect 974 -5396 980 -5362
rect 1014 -5396 1020 -5362
rect 974 -5434 1020 -5396
rect 974 -5468 980 -5434
rect 1014 -5468 1020 -5434
rect 974 -5506 1020 -5468
rect 974 -5540 980 -5506
rect 1014 -5540 1020 -5506
rect 974 -5563 1020 -5540
rect 1070 -4786 1116 -4744
rect 1070 -4820 1076 -4786
rect 1110 -4820 1116 -4786
rect 1070 -4858 1116 -4820
rect 1070 -4892 1076 -4858
rect 1110 -4892 1116 -4858
rect 1070 -4930 1116 -4892
rect 1070 -4964 1076 -4930
rect 1110 -4964 1116 -4930
rect 1070 -5002 1116 -4964
rect 1070 -5036 1076 -5002
rect 1110 -5036 1116 -5002
rect 1070 -5074 1116 -5036
rect 1070 -5108 1076 -5074
rect 1110 -5108 1116 -5074
rect 1070 -5146 1116 -5108
rect 1070 -5180 1076 -5146
rect 1110 -5180 1116 -5146
rect 1070 -5218 1116 -5180
rect 1070 -5252 1076 -5218
rect 1110 -5252 1116 -5218
rect 1070 -5290 1116 -5252
rect 1070 -5324 1076 -5290
rect 1110 -5324 1116 -5290
rect 1070 -5362 1116 -5324
rect 1070 -5396 1076 -5362
rect 1110 -5396 1116 -5362
rect 1070 -5434 1116 -5396
rect 1070 -5468 1076 -5434
rect 1110 -5468 1116 -5434
rect 1070 -5506 1116 -5468
rect 1070 -5540 1076 -5506
rect 1110 -5540 1116 -5506
rect 1070 -5790 1116 -5540
rect 1166 -4786 1212 -4569
rect 1166 -4820 1172 -4786
rect 1206 -4820 1212 -4786
rect 1166 -4858 1212 -4820
rect 1166 -4892 1172 -4858
rect 1206 -4892 1212 -4858
rect 1166 -4930 1212 -4892
rect 1166 -4964 1172 -4930
rect 1206 -4964 1212 -4930
rect 1166 -5002 1212 -4964
rect 1166 -5036 1172 -5002
rect 1206 -5036 1212 -5002
rect 1166 -5074 1212 -5036
rect 1166 -5108 1172 -5074
rect 1206 -5108 1212 -5074
rect 1166 -5146 1212 -5108
rect 1166 -5180 1172 -5146
rect 1206 -5180 1212 -5146
rect 1166 -5218 1212 -5180
rect 1166 -5252 1172 -5218
rect 1206 -5252 1212 -5218
rect 1166 -5290 1212 -5252
rect 1166 -5324 1172 -5290
rect 1206 -5324 1212 -5290
rect 1166 -5362 1212 -5324
rect 1166 -5396 1172 -5362
rect 1206 -5396 1212 -5362
rect 1166 -5434 1212 -5396
rect 1166 -5468 1172 -5434
rect 1206 -5468 1212 -5434
rect 1166 -5506 1212 -5468
rect 1166 -5540 1172 -5506
rect 1206 -5540 1212 -5506
rect 1166 -5563 1212 -5540
rect 1262 -4786 1308 -4744
rect 1262 -4820 1268 -4786
rect 1302 -4820 1308 -4786
rect 1262 -4858 1308 -4820
rect 1262 -4892 1268 -4858
rect 1302 -4892 1308 -4858
rect 1262 -4930 1308 -4892
rect 1262 -4964 1268 -4930
rect 1302 -4964 1308 -4930
rect 1262 -5002 1308 -4964
rect 1262 -5036 1268 -5002
rect 1302 -5036 1308 -5002
rect 1262 -5074 1308 -5036
rect 1262 -5108 1268 -5074
rect 1302 -5108 1308 -5074
rect 1262 -5146 1308 -5108
rect 1262 -5180 1268 -5146
rect 1302 -5180 1308 -5146
rect 1262 -5218 1308 -5180
rect 1262 -5252 1268 -5218
rect 1302 -5252 1308 -5218
rect 1262 -5290 1308 -5252
rect 1262 -5324 1268 -5290
rect 1302 -5324 1308 -5290
rect 1262 -5362 1308 -5324
rect 1262 -5396 1268 -5362
rect 1302 -5396 1308 -5362
rect 1262 -5434 1308 -5396
rect 1262 -5468 1268 -5434
rect 1302 -5468 1308 -5434
rect 1262 -5506 1308 -5468
rect 1262 -5540 1268 -5506
rect 1302 -5540 1308 -5506
rect 1262 -5790 1308 -5540
rect 1358 -4786 1404 -4569
rect 1358 -4820 1364 -4786
rect 1398 -4820 1404 -4786
rect 1358 -4858 1404 -4820
rect 1358 -4892 1364 -4858
rect 1398 -4892 1404 -4858
rect 1358 -4930 1404 -4892
rect 1358 -4964 1364 -4930
rect 1398 -4964 1404 -4930
rect 1358 -5002 1404 -4964
rect 1358 -5036 1364 -5002
rect 1398 -5036 1404 -5002
rect 1358 -5074 1404 -5036
rect 1358 -5108 1364 -5074
rect 1398 -5108 1404 -5074
rect 1358 -5146 1404 -5108
rect 1358 -5180 1364 -5146
rect 1398 -5180 1404 -5146
rect 1358 -5218 1404 -5180
rect 1358 -5252 1364 -5218
rect 1398 -5252 1404 -5218
rect 1358 -5290 1404 -5252
rect 1358 -5324 1364 -5290
rect 1398 -5324 1404 -5290
rect 1358 -5362 1404 -5324
rect 1358 -5396 1364 -5362
rect 1398 -5396 1404 -5362
rect 1358 -5434 1404 -5396
rect 1358 -5468 1364 -5434
rect 1398 -5468 1404 -5434
rect 1358 -5506 1404 -5468
rect 1358 -5540 1364 -5506
rect 1398 -5540 1404 -5506
rect 1358 -5563 1404 -5540
rect 1454 -4786 1500 -4744
rect 1454 -4820 1460 -4786
rect 1494 -4820 1500 -4786
rect 1454 -4858 1500 -4820
rect 1454 -4892 1460 -4858
rect 1494 -4892 1500 -4858
rect 1454 -4930 1500 -4892
rect 1454 -4964 1460 -4930
rect 1494 -4964 1500 -4930
rect 1454 -5002 1500 -4964
rect 1454 -5036 1460 -5002
rect 1494 -5036 1500 -5002
rect 1454 -5074 1500 -5036
rect 1454 -5108 1460 -5074
rect 1494 -5108 1500 -5074
rect 1454 -5146 1500 -5108
rect 1454 -5180 1460 -5146
rect 1494 -5180 1500 -5146
rect 1454 -5218 1500 -5180
rect 1454 -5252 1460 -5218
rect 1494 -5252 1500 -5218
rect 1454 -5290 1500 -5252
rect 1454 -5324 1460 -5290
rect 1494 -5324 1500 -5290
rect 1454 -5362 1500 -5324
rect 1454 -5396 1460 -5362
rect 1494 -5396 1500 -5362
rect 1454 -5434 1500 -5396
rect 1454 -5468 1460 -5434
rect 1494 -5468 1500 -5434
rect 1454 -5506 1500 -5468
rect 1454 -5540 1460 -5506
rect 1494 -5540 1500 -5506
rect 1454 -5790 1500 -5540
rect 1550 -4786 1596 -4569
rect 1550 -4820 1556 -4786
rect 1590 -4820 1596 -4786
rect 1550 -4858 1596 -4820
rect 1550 -4892 1556 -4858
rect 1590 -4892 1596 -4858
rect 1550 -4930 1596 -4892
rect 1550 -4964 1556 -4930
rect 1590 -4964 1596 -4930
rect 1550 -5002 1596 -4964
rect 1550 -5036 1556 -5002
rect 1590 -5036 1596 -5002
rect 1550 -5074 1596 -5036
rect 1550 -5108 1556 -5074
rect 1590 -5108 1596 -5074
rect 1550 -5146 1596 -5108
rect 1550 -5180 1556 -5146
rect 1590 -5180 1596 -5146
rect 1550 -5218 1596 -5180
rect 1550 -5252 1556 -5218
rect 1590 -5252 1596 -5218
rect 1550 -5290 1596 -5252
rect 1550 -5324 1556 -5290
rect 1590 -5324 1596 -5290
rect 1550 -5362 1596 -5324
rect 1550 -5396 1556 -5362
rect 1590 -5396 1596 -5362
rect 1550 -5434 1596 -5396
rect 1550 -5468 1556 -5434
rect 1590 -5468 1596 -5434
rect 1550 -5506 1596 -5468
rect 1550 -5540 1556 -5506
rect 1590 -5540 1596 -5506
rect 1550 -5563 1596 -5540
rect 1646 -4786 1692 -4744
rect 1646 -4820 1652 -4786
rect 1686 -4820 1692 -4786
rect 1646 -4858 1692 -4820
rect 1646 -4892 1652 -4858
rect 1686 -4892 1692 -4858
rect 1646 -4930 1692 -4892
rect 1646 -4964 1652 -4930
rect 1686 -4964 1692 -4930
rect 1646 -5002 1692 -4964
rect 1646 -5036 1652 -5002
rect 1686 -5036 1692 -5002
rect 1646 -5074 1692 -5036
rect 1646 -5108 1652 -5074
rect 1686 -5108 1692 -5074
rect 1646 -5146 1692 -5108
rect 1646 -5180 1652 -5146
rect 1686 -5180 1692 -5146
rect 1646 -5218 1692 -5180
rect 1646 -5252 1652 -5218
rect 1686 -5252 1692 -5218
rect 1646 -5290 1692 -5252
rect 1646 -5324 1652 -5290
rect 1686 -5324 1692 -5290
rect 1646 -5362 1692 -5324
rect 1646 -5396 1652 -5362
rect 1686 -5396 1692 -5362
rect 1646 -5434 1692 -5396
rect 1646 -5468 1652 -5434
rect 1686 -5468 1692 -5434
rect 1646 -5506 1692 -5468
rect 1646 -5540 1652 -5506
rect 1686 -5540 1692 -5506
rect 1646 -5790 1692 -5540
rect 1742 -4786 1788 -4569
rect 1742 -4820 1748 -4786
rect 1782 -4820 1788 -4786
rect 1742 -4858 1788 -4820
rect 1742 -4892 1748 -4858
rect 1782 -4892 1788 -4858
rect 1742 -4930 1788 -4892
rect 1742 -4964 1748 -4930
rect 1782 -4964 1788 -4930
rect 1742 -5002 1788 -4964
rect 1742 -5036 1748 -5002
rect 1782 -5036 1788 -5002
rect 1742 -5074 1788 -5036
rect 1742 -5108 1748 -5074
rect 1782 -5108 1788 -5074
rect 1742 -5146 1788 -5108
rect 1742 -5180 1748 -5146
rect 1782 -5180 1788 -5146
rect 1742 -5218 1788 -5180
rect 1742 -5252 1748 -5218
rect 1782 -5252 1788 -5218
rect 1742 -5290 1788 -5252
rect 1742 -5324 1748 -5290
rect 1782 -5324 1788 -5290
rect 1742 -5362 1788 -5324
rect 1742 -5396 1748 -5362
rect 1782 -5396 1788 -5362
rect 1742 -5434 1788 -5396
rect 1742 -5468 1748 -5434
rect 1782 -5468 1788 -5434
rect 1742 -5506 1788 -5468
rect 1742 -5540 1748 -5506
rect 1782 -5540 1788 -5506
rect 1742 -5563 1788 -5540
rect 1838 -4786 1884 -4744
rect 1838 -4820 1844 -4786
rect 1878 -4820 1884 -4786
rect 1838 -4858 1884 -4820
rect 1838 -4892 1844 -4858
rect 1878 -4892 1884 -4858
rect 1838 -4930 1884 -4892
rect 1838 -4964 1844 -4930
rect 1878 -4964 1884 -4930
rect 1838 -5002 1884 -4964
rect 1838 -5036 1844 -5002
rect 1878 -5036 1884 -5002
rect 1838 -5074 1884 -5036
rect 1838 -5108 1844 -5074
rect 1878 -5108 1884 -5074
rect 1838 -5146 1884 -5108
rect 1838 -5180 1844 -5146
rect 1878 -5180 1884 -5146
rect 1838 -5218 1884 -5180
rect 1838 -5252 1844 -5218
rect 1878 -5252 1884 -5218
rect 1838 -5290 1884 -5252
rect 1838 -5324 1844 -5290
rect 1878 -5324 1884 -5290
rect 1838 -5362 1884 -5324
rect 1838 -5396 1844 -5362
rect 1878 -5396 1884 -5362
rect 1838 -5434 1884 -5396
rect 1838 -5468 1844 -5434
rect 1878 -5468 1884 -5434
rect 1838 -5506 1884 -5468
rect 1838 -5540 1844 -5506
rect 1878 -5540 1884 -5506
rect 1838 -5790 1884 -5540
rect 1934 -4786 1980 -4569
rect 1934 -4820 1940 -4786
rect 1974 -4820 1980 -4786
rect 1934 -4858 1980 -4820
rect 1934 -4892 1940 -4858
rect 1974 -4892 1980 -4858
rect 1934 -4930 1980 -4892
rect 1934 -4964 1940 -4930
rect 1974 -4964 1980 -4930
rect 1934 -5002 1980 -4964
rect 1934 -5036 1940 -5002
rect 1974 -5036 1980 -5002
rect 1934 -5074 1980 -5036
rect 1934 -5108 1940 -5074
rect 1974 -5108 1980 -5074
rect 1934 -5146 1980 -5108
rect 1934 -5180 1940 -5146
rect 1974 -5180 1980 -5146
rect 1934 -5218 1980 -5180
rect 1934 -5252 1940 -5218
rect 1974 -5252 1980 -5218
rect 1934 -5290 1980 -5252
rect 1934 -5324 1940 -5290
rect 1974 -5324 1980 -5290
rect 1934 -5362 1980 -5324
rect 1934 -5396 1940 -5362
rect 1974 -5396 1980 -5362
rect 1934 -5434 1980 -5396
rect 1934 -5468 1940 -5434
rect 1974 -5468 1980 -5434
rect 1934 -5506 1980 -5468
rect 1934 -5540 1940 -5506
rect 1974 -5540 1980 -5506
rect 1934 -5563 1980 -5540
rect -42440 -7880 -40660 -5934
rect -42440 -13820 -42408 -7880
rect -40692 -13820 -40660 -7880
rect -42440 -13850 -40660 -13820
rect 110 -7880 1890 -5790
rect 110 -13820 142 -7880
rect 1858 -13820 1890 -7880
rect 110 -13850 1890 -13820
rect 2605 -13850 2675 13850
rect 3265 -13850 3335 13850
rect 3925 -13850 3995 13850
rect 4585 -13850 4655 13850
rect 5245 -13850 5315 13850
rect 5905 -13850 5975 13850
rect 6565 -13850 6635 13850
rect 7225 -13850 7295 13850
rect 7885 -13850 7955 13850
rect 8545 -13850 8615 13850
rect 9205 -13850 9275 13850
rect 9865 -13850 9935 13850
rect 10525 -13850 10595 13850
rect 11185 -13850 11255 13850
rect 11845 -13850 11915 13850
rect 12505 -13850 12575 13850
rect 13165 -13850 13235 13850
rect 13825 -13850 13895 13850
rect 14485 -13850 14555 13850
rect 15145 -13850 15215 13850
rect 15805 -13850 15875 13850
rect 16465 -13850 16535 13850
rect 20275 7600 32275 16046
rect 21575 -7600 23075 7600
rect 23875 -7600 25375 7600
rect 26175 -7600 27675 7600
rect 28475 -7600 29975 7600
rect 30775 -7600 32275 7600
rect -34125 -14320 -6425 -14250
rect -34125 -14980 -6425 -14910
rect -34125 -15640 -6425 -15570
rect -72825 -25954 -72776 -16046
rect -60884 -25954 -60825 -16046
rect 20275 -16046 32275 -7600
rect -34125 -16300 -6425 -16230
rect -34125 -16960 -6425 -16890
rect -34125 -17620 -6425 -17550
rect -34125 -18280 -6425 -18210
rect -34125 -18940 -6425 -18870
rect -34125 -19600 -6425 -19530
rect -34125 -20260 -6425 -20190
rect -34125 -20920 -6425 -20850
rect -34125 -21580 -6425 -21510
rect -34125 -22240 -6425 -22170
rect -34125 -22900 -6425 -22830
rect -34125 -23560 -6425 -23490
rect -34125 -24220 -6425 -24150
rect -34125 -24880 -6425 -24810
rect -34125 -25540 -6425 -25470
rect -72825 -26000 -60825 -25954
rect 20275 -25954 20324 -16046
rect 32216 -25954 32275 -16046
rect 20275 -26000 32275 -25954
rect -34125 -26200 -6425 -26130
rect -34125 -26860 -6425 -26790
rect -74485 -28556 -74165 -28550
rect -74485 -28864 -74479 -28556
rect -74171 -28864 -74165 -28556
rect -74485 -28890 -74165 -28864
rect -73485 -28556 -73165 -28550
rect -73485 -28864 -73479 -28556
rect -73171 -28864 -73165 -28556
rect -73485 -28890 -73165 -28864
rect -72485 -28556 -72165 -28550
rect -72485 -28864 -72479 -28556
rect -72171 -28864 -72165 -28556
rect -72485 -28890 -72165 -28864
rect -71485 -28556 -71165 -28550
rect -71485 -28864 -71479 -28556
rect -71171 -28864 -71165 -28556
rect -71485 -28890 -71165 -28864
rect -70485 -28556 -70165 -28550
rect -70485 -28864 -70479 -28556
rect -70171 -28864 -70165 -28556
rect -70485 -28890 -70165 -28864
rect -69485 -28556 -69165 -28550
rect -69485 -28864 -69479 -28556
rect -69171 -28864 -69165 -28556
rect -69485 -28890 -69165 -28864
rect -68485 -28556 -68165 -28550
rect -68485 -28864 -68479 -28556
rect -68171 -28864 -68165 -28556
rect -68485 -28890 -68165 -28864
rect -67485 -28556 -67165 -28550
rect -67485 -28864 -67479 -28556
rect -67171 -28864 -67165 -28556
rect -67485 -28890 -67165 -28864
rect -66485 -28556 -66165 -28550
rect -66485 -28864 -66479 -28556
rect -66171 -28864 -66165 -28556
rect -66485 -28890 -66165 -28864
rect -65485 -28556 -65165 -28550
rect -65485 -28864 -65479 -28556
rect -65171 -28864 -65165 -28556
rect -65485 -28890 -65165 -28864
rect -64485 -28556 -64165 -28550
rect -64485 -28864 -64479 -28556
rect -64171 -28864 -64165 -28556
rect -64485 -28890 -64165 -28864
rect -63485 -28556 -63165 -28550
rect -63485 -28864 -63479 -28556
rect -63171 -28864 -63165 -28556
rect -63485 -28890 -63165 -28864
rect -62485 -28556 -62165 -28550
rect -62485 -28864 -62479 -28556
rect -62171 -28864 -62165 -28556
rect -62485 -28890 -62165 -28864
rect -61485 -28556 -61165 -28550
rect -61485 -28864 -61479 -28556
rect -61171 -28864 -61165 -28556
rect -61485 -28890 -61165 -28864
rect -60485 -28556 -60165 -28550
rect -60485 -28864 -60479 -28556
rect -60171 -28864 -60165 -28556
rect -60485 -28890 -60165 -28864
rect -59485 -28556 -59165 -28550
rect -59485 -28864 -59479 -28556
rect -59171 -28864 -59165 -28556
rect -59485 -28890 -59165 -28864
rect -58485 -28556 -58165 -28550
rect -58485 -28864 -58479 -28556
rect -58171 -28864 -58165 -28556
rect -58485 -28890 -58165 -28864
rect -57485 -28556 -57165 -28550
rect -57485 -28864 -57479 -28556
rect -57171 -28864 -57165 -28556
rect -57485 -28890 -57165 -28864
rect -56485 -28556 -56165 -28550
rect -56485 -28864 -56479 -28556
rect -56171 -28864 -56165 -28556
rect -56485 -28890 -56165 -28864
rect -55485 -28556 -55165 -28550
rect -55485 -28864 -55479 -28556
rect -55171 -28864 -55165 -28556
rect -55485 -28890 -55165 -28864
rect -54485 -28556 -54165 -28550
rect -54485 -28864 -54479 -28556
rect -54171 -28864 -54165 -28556
rect -54485 -28890 -54165 -28864
rect -53485 -28556 -53165 -28550
rect -53485 -28864 -53479 -28556
rect -53171 -28864 -53165 -28556
rect -53485 -28890 -53165 -28864
rect -52485 -28556 -52165 -28550
rect -52485 -28864 -52479 -28556
rect -52171 -28864 -52165 -28556
rect -52485 -28890 -52165 -28864
rect -51485 -28556 -51165 -28550
rect -51485 -28864 -51479 -28556
rect -51171 -28864 -51165 -28556
rect -51485 -28890 -51165 -28864
rect -50485 -28556 -50165 -28550
rect -50485 -28864 -50479 -28556
rect -50171 -28864 -50165 -28556
rect -50485 -28890 -50165 -28864
rect -49485 -28556 -49165 -28550
rect -49485 -28864 -49479 -28556
rect -49171 -28864 -49165 -28556
rect -49485 -28890 -49165 -28864
rect 8615 -28556 8935 -28550
rect 8615 -28864 8621 -28556
rect 8929 -28864 8935 -28556
rect 8615 -28890 8935 -28864
rect 9615 -28556 9935 -28550
rect 9615 -28864 9621 -28556
rect 9929 -28864 9935 -28556
rect 9615 -28890 9935 -28864
rect 10615 -28556 10935 -28550
rect 10615 -28864 10621 -28556
rect 10929 -28864 10935 -28556
rect 10615 -28890 10935 -28864
rect 11615 -28556 11935 -28550
rect 11615 -28864 11621 -28556
rect 11929 -28864 11935 -28556
rect 11615 -28890 11935 -28864
rect 12615 -28556 12935 -28550
rect 12615 -28864 12621 -28556
rect 12929 -28864 12935 -28556
rect 12615 -28890 12935 -28864
rect 13615 -28556 13935 -28550
rect 13615 -28864 13621 -28556
rect 13929 -28864 13935 -28556
rect 13615 -28890 13935 -28864
rect 14615 -28556 14935 -28550
rect 14615 -28864 14621 -28556
rect 14929 -28864 14935 -28556
rect 14615 -28890 14935 -28864
rect 15615 -28556 15935 -28550
rect 15615 -28864 15621 -28556
rect 15929 -28864 15935 -28556
rect 15615 -28890 15935 -28864
rect 16615 -28556 16935 -28550
rect 16615 -28864 16621 -28556
rect 16929 -28864 16935 -28556
rect 16615 -28890 16935 -28864
rect 17615 -28556 17935 -28550
rect 17615 -28864 17621 -28556
rect 17929 -28864 17935 -28556
rect 17615 -28890 17935 -28864
rect 18615 -28556 18935 -28550
rect 18615 -28864 18621 -28556
rect 18929 -28864 18935 -28556
rect 18615 -28890 18935 -28864
rect 19615 -28556 19935 -28550
rect 19615 -28864 19621 -28556
rect 19929 -28864 19935 -28556
rect 19615 -28890 19935 -28864
rect 20615 -28556 20935 -28550
rect 20615 -28864 20621 -28556
rect 20929 -28864 20935 -28556
rect 20615 -28890 20935 -28864
rect 21615 -28556 21935 -28550
rect 21615 -28864 21621 -28556
rect 21929 -28864 21935 -28556
rect 21615 -28890 21935 -28864
rect 22615 -28556 22935 -28550
rect 22615 -28864 22621 -28556
rect 22929 -28864 22935 -28556
rect 22615 -28890 22935 -28864
rect 23615 -28556 23935 -28550
rect 23615 -28864 23621 -28556
rect 23929 -28864 23935 -28556
rect 23615 -28890 23935 -28864
rect 24615 -28556 24935 -28550
rect 24615 -28864 24621 -28556
rect 24929 -28864 24935 -28556
rect 24615 -28890 24935 -28864
rect 25615 -28556 25935 -28550
rect 25615 -28864 25621 -28556
rect 25929 -28864 25935 -28556
rect 25615 -28890 25935 -28864
rect 26615 -28556 26935 -28550
rect 26615 -28864 26621 -28556
rect 26929 -28864 26935 -28556
rect 26615 -28890 26935 -28864
rect 27615 -28556 27935 -28550
rect 27615 -28864 27621 -28556
rect 27929 -28864 27935 -28556
rect 27615 -28890 27935 -28864
rect 28615 -28556 28935 -28550
rect 28615 -28864 28621 -28556
rect 28929 -28864 28935 -28556
rect 28615 -28890 28935 -28864
rect 29615 -28556 29935 -28550
rect 29615 -28864 29621 -28556
rect 29929 -28864 29935 -28556
rect 29615 -28890 29935 -28864
rect 30615 -28556 30935 -28550
rect 30615 -28864 30621 -28556
rect 30929 -28864 30935 -28556
rect 30615 -28890 30935 -28864
rect 31615 -28556 31935 -28550
rect 31615 -28864 31621 -28556
rect 31929 -28864 31935 -28556
rect 31615 -28890 31935 -28864
rect 32615 -28556 32935 -28550
rect 32615 -28864 32621 -28556
rect 32929 -28864 32935 -28556
rect 32615 -28890 32935 -28864
rect 33615 -28556 33935 -28550
rect 33615 -28864 33621 -28556
rect 33929 -28864 33935 -28556
rect 33615 -28890 33935 -28864
rect -74825 -28896 -48825 -28890
rect -74825 -29204 -74819 -28896
rect -74511 -28928 -74139 -28896
rect -74511 -29172 -74447 -28928
rect -74203 -29172 -74139 -28928
rect -74511 -29204 -74139 -29172
rect -73511 -28928 -73139 -28896
rect -73511 -29172 -73447 -28928
rect -73203 -29172 -73139 -28928
rect -73511 -29204 -73139 -29172
rect -72511 -28928 -72139 -28896
rect -72511 -29172 -72447 -28928
rect -72203 -29172 -72139 -28928
rect -72511 -29204 -72139 -29172
rect -71511 -28928 -71139 -28896
rect -71511 -29172 -71447 -28928
rect -71203 -29172 -71139 -28928
rect -71511 -29204 -71139 -29172
rect -70511 -28928 -70139 -28896
rect -70511 -29172 -70447 -28928
rect -70203 -29172 -70139 -28928
rect -70511 -29204 -70139 -29172
rect -69511 -28928 -69139 -28896
rect -69511 -29172 -69447 -28928
rect -69203 -29172 -69139 -28928
rect -69511 -29204 -69139 -29172
rect -68511 -28928 -68139 -28896
rect -68511 -29172 -68447 -28928
rect -68203 -29172 -68139 -28928
rect -68511 -29204 -68139 -29172
rect -67511 -28928 -67139 -28896
rect -67511 -29172 -67447 -28928
rect -67203 -29172 -67139 -28928
rect -67511 -29204 -67139 -29172
rect -66511 -28928 -66139 -28896
rect -66511 -29172 -66447 -28928
rect -66203 -29172 -66139 -28928
rect -66511 -29204 -66139 -29172
rect -65511 -28928 -65139 -28896
rect -65511 -29172 -65447 -28928
rect -65203 -29172 -65139 -28928
rect -65511 -29204 -65139 -29172
rect -64511 -28928 -64139 -28896
rect -64511 -29172 -64447 -28928
rect -64203 -29172 -64139 -28928
rect -64511 -29204 -64139 -29172
rect -63511 -28928 -63139 -28896
rect -63511 -29172 -63447 -28928
rect -63203 -29172 -63139 -28928
rect -63511 -29204 -63139 -29172
rect -62511 -28928 -62139 -28896
rect -62511 -29172 -62447 -28928
rect -62203 -29172 -62139 -28928
rect -62511 -29204 -62139 -29172
rect -61511 -28928 -61139 -28896
rect -61511 -29172 -61447 -28928
rect -61203 -29172 -61139 -28928
rect -61511 -29204 -61139 -29172
rect -60511 -28928 -60139 -28896
rect -60511 -29172 -60447 -28928
rect -60203 -29172 -60139 -28928
rect -60511 -29204 -60139 -29172
rect -59511 -28928 -59139 -28896
rect -59511 -29172 -59447 -28928
rect -59203 -29172 -59139 -28928
rect -59511 -29204 -59139 -29172
rect -58511 -28928 -58139 -28896
rect -58511 -29172 -58447 -28928
rect -58203 -29172 -58139 -28928
rect -58511 -29204 -58139 -29172
rect -57511 -28928 -57139 -28896
rect -57511 -29172 -57447 -28928
rect -57203 -29172 -57139 -28928
rect -57511 -29204 -57139 -29172
rect -56511 -28928 -56139 -28896
rect -56511 -29172 -56447 -28928
rect -56203 -29172 -56139 -28928
rect -56511 -29204 -56139 -29172
rect -55511 -28928 -55139 -28896
rect -55511 -29172 -55447 -28928
rect -55203 -29172 -55139 -28928
rect -55511 -29204 -55139 -29172
rect -54511 -28928 -54139 -28896
rect -54511 -29172 -54447 -28928
rect -54203 -29172 -54139 -28928
rect -54511 -29204 -54139 -29172
rect -53511 -28928 -53139 -28896
rect -53511 -29172 -53447 -28928
rect -53203 -29172 -53139 -28928
rect -53511 -29204 -53139 -29172
rect -52511 -28928 -52139 -28896
rect -52511 -29172 -52447 -28928
rect -52203 -29172 -52139 -28928
rect -52511 -29204 -52139 -29172
rect -51511 -28928 -51139 -28896
rect -51511 -29172 -51447 -28928
rect -51203 -29172 -51139 -28928
rect -51511 -29204 -51139 -29172
rect -50511 -28928 -50139 -28896
rect -50511 -29172 -50447 -28928
rect -50203 -29172 -50139 -28928
rect -50511 -29204 -50139 -29172
rect -49511 -28928 -49139 -28896
rect -49511 -29172 -49447 -28928
rect -49203 -29172 -49139 -28928
rect -49511 -29204 -49139 -29172
rect -48831 -29204 -48825 -28896
rect -74825 -29210 -48825 -29204
rect 8275 -28896 34275 -28890
rect 8275 -29204 8281 -28896
rect 8589 -28928 8961 -28896
rect 8589 -29172 8653 -28928
rect 8897 -29172 8961 -28928
rect 8589 -29204 8961 -29172
rect 9589 -28928 9961 -28896
rect 9589 -29172 9653 -28928
rect 9897 -29172 9961 -28928
rect 9589 -29204 9961 -29172
rect 10589 -28928 10961 -28896
rect 10589 -29172 10653 -28928
rect 10897 -29172 10961 -28928
rect 10589 -29204 10961 -29172
rect 11589 -28928 11961 -28896
rect 11589 -29172 11653 -28928
rect 11897 -29172 11961 -28928
rect 11589 -29204 11961 -29172
rect 12589 -28928 12961 -28896
rect 12589 -29172 12653 -28928
rect 12897 -29172 12961 -28928
rect 12589 -29204 12961 -29172
rect 13589 -28928 13961 -28896
rect 13589 -29172 13653 -28928
rect 13897 -29172 13961 -28928
rect 13589 -29204 13961 -29172
rect 14589 -28928 14961 -28896
rect 14589 -29172 14653 -28928
rect 14897 -29172 14961 -28928
rect 14589 -29204 14961 -29172
rect 15589 -28928 15961 -28896
rect 15589 -29172 15653 -28928
rect 15897 -29172 15961 -28928
rect 15589 -29204 15961 -29172
rect 16589 -28928 16961 -28896
rect 16589 -29172 16653 -28928
rect 16897 -29172 16961 -28928
rect 16589 -29204 16961 -29172
rect 17589 -28928 17961 -28896
rect 17589 -29172 17653 -28928
rect 17897 -29172 17961 -28928
rect 17589 -29204 17961 -29172
rect 18589 -28928 18961 -28896
rect 18589 -29172 18653 -28928
rect 18897 -29172 18961 -28928
rect 18589 -29204 18961 -29172
rect 19589 -28928 19961 -28896
rect 19589 -29172 19653 -28928
rect 19897 -29172 19961 -28928
rect 19589 -29204 19961 -29172
rect 20589 -28928 20961 -28896
rect 20589 -29172 20653 -28928
rect 20897 -29172 20961 -28928
rect 20589 -29204 20961 -29172
rect 21589 -28928 21961 -28896
rect 21589 -29172 21653 -28928
rect 21897 -29172 21961 -28928
rect 21589 -29204 21961 -29172
rect 22589 -28928 22961 -28896
rect 22589 -29172 22653 -28928
rect 22897 -29172 22961 -28928
rect 22589 -29204 22961 -29172
rect 23589 -28928 23961 -28896
rect 23589 -29172 23653 -28928
rect 23897 -29172 23961 -28928
rect 23589 -29204 23961 -29172
rect 24589 -28928 24961 -28896
rect 24589 -29172 24653 -28928
rect 24897 -29172 24961 -28928
rect 24589 -29204 24961 -29172
rect 25589 -28928 25961 -28896
rect 25589 -29172 25653 -28928
rect 25897 -29172 25961 -28928
rect 25589 -29204 25961 -29172
rect 26589 -28928 26961 -28896
rect 26589 -29172 26653 -28928
rect 26897 -29172 26961 -28928
rect 26589 -29204 26961 -29172
rect 27589 -28928 27961 -28896
rect 27589 -29172 27653 -28928
rect 27897 -29172 27961 -28928
rect 27589 -29204 27961 -29172
rect 28589 -28928 28961 -28896
rect 28589 -29172 28653 -28928
rect 28897 -29172 28961 -28928
rect 28589 -29204 28961 -29172
rect 29589 -28928 29961 -28896
rect 29589 -29172 29653 -28928
rect 29897 -29172 29961 -28928
rect 29589 -29204 29961 -29172
rect 30589 -28928 30961 -28896
rect 30589 -29172 30653 -28928
rect 30897 -29172 30961 -28928
rect 30589 -29204 30961 -29172
rect 31589 -28928 31961 -28896
rect 31589 -29172 31653 -28928
rect 31897 -29172 31961 -28928
rect 31589 -29204 31961 -29172
rect 32589 -28928 32961 -28896
rect 32589 -29172 32653 -28928
rect 32897 -29172 32961 -28928
rect 32589 -29204 32961 -29172
rect 33589 -28928 33961 -28896
rect 33589 -29172 33653 -28928
rect 33897 -29172 33961 -28928
rect 33589 -29204 33961 -29172
rect 34269 -29204 34275 -28896
rect 8275 -29210 34275 -29204
rect -74485 -29236 -74165 -29210
rect -74485 -29864 -74479 -29236
rect -74171 -29864 -74165 -29236
rect -74485 -29890 -74165 -29864
rect -73485 -29236 -73165 -29210
rect -73485 -29864 -73479 -29236
rect -73171 -29864 -73165 -29236
rect -73485 -29890 -73165 -29864
rect -72485 -29236 -72165 -29210
rect -72485 -29864 -72479 -29236
rect -72171 -29864 -72165 -29236
rect -72485 -29890 -72165 -29864
rect -71485 -29236 -71165 -29210
rect -71485 -29864 -71479 -29236
rect -71171 -29864 -71165 -29236
rect -71485 -29890 -71165 -29864
rect -70485 -29236 -70165 -29210
rect -70485 -29864 -70479 -29236
rect -70171 -29864 -70165 -29236
rect -70485 -29890 -70165 -29864
rect -69485 -29236 -69165 -29210
rect -69485 -29864 -69479 -29236
rect -69171 -29864 -69165 -29236
rect -69485 -29890 -69165 -29864
rect -68485 -29236 -68165 -29210
rect -68485 -29864 -68479 -29236
rect -68171 -29864 -68165 -29236
rect -68485 -29890 -68165 -29864
rect -67485 -29236 -67165 -29210
rect -67485 -29864 -67479 -29236
rect -67171 -29864 -67165 -29236
rect -67485 -29890 -67165 -29864
rect -66485 -29236 -66165 -29210
rect -66485 -29864 -66479 -29236
rect -66171 -29864 -66165 -29236
rect -66485 -29890 -66165 -29864
rect -65485 -29236 -65165 -29210
rect -65485 -29864 -65479 -29236
rect -65171 -29864 -65165 -29236
rect -65485 -29890 -65165 -29864
rect -64485 -29236 -64165 -29210
rect -64485 -29864 -64479 -29236
rect -64171 -29864 -64165 -29236
rect -64485 -29890 -64165 -29864
rect -63485 -29236 -63165 -29210
rect -63485 -29864 -63479 -29236
rect -63171 -29864 -63165 -29236
rect -63485 -29890 -63165 -29864
rect -62485 -29236 -62165 -29210
rect -62485 -29864 -62479 -29236
rect -62171 -29864 -62165 -29236
rect -62485 -29890 -62165 -29864
rect -61485 -29236 -61165 -29210
rect -61485 -29864 -61479 -29236
rect -61171 -29864 -61165 -29236
rect -61485 -29890 -61165 -29864
rect -60485 -29236 -60165 -29210
rect -60485 -29864 -60479 -29236
rect -60171 -29864 -60165 -29236
rect -60485 -29890 -60165 -29864
rect -59485 -29236 -59165 -29210
rect -59485 -29864 -59479 -29236
rect -59171 -29864 -59165 -29236
rect -59485 -29890 -59165 -29864
rect -58485 -29236 -58165 -29210
rect -58485 -29864 -58479 -29236
rect -58171 -29864 -58165 -29236
rect -58485 -29890 -58165 -29864
rect -57485 -29236 -57165 -29210
rect -57485 -29864 -57479 -29236
rect -57171 -29864 -57165 -29236
rect -57485 -29890 -57165 -29864
rect -56485 -29236 -56165 -29210
rect -56485 -29864 -56479 -29236
rect -56171 -29864 -56165 -29236
rect -56485 -29890 -56165 -29864
rect -55485 -29236 -55165 -29210
rect -55485 -29864 -55479 -29236
rect -55171 -29864 -55165 -29236
rect -55485 -29890 -55165 -29864
rect -54485 -29236 -54165 -29210
rect -54485 -29864 -54479 -29236
rect -54171 -29864 -54165 -29236
rect -54485 -29890 -54165 -29864
rect -53485 -29236 -53165 -29210
rect -53485 -29864 -53479 -29236
rect -53171 -29864 -53165 -29236
rect -53485 -29890 -53165 -29864
rect -52485 -29236 -52165 -29210
rect -52485 -29864 -52479 -29236
rect -52171 -29864 -52165 -29236
rect -52485 -29890 -52165 -29864
rect -51485 -29236 -51165 -29210
rect -51485 -29864 -51479 -29236
rect -51171 -29864 -51165 -29236
rect -51485 -29890 -51165 -29864
rect -50485 -29236 -50165 -29210
rect -50485 -29864 -50479 -29236
rect -50171 -29864 -50165 -29236
rect -50485 -29890 -50165 -29864
rect -49485 -29236 -49165 -29210
rect -49485 -29864 -49479 -29236
rect -49171 -29864 -49165 -29236
rect -49485 -29890 -49165 -29864
rect 8615 -29236 8935 -29210
rect 8615 -29864 8621 -29236
rect 8929 -29864 8935 -29236
rect 8615 -29890 8935 -29864
rect 9615 -29236 9935 -29210
rect 9615 -29864 9621 -29236
rect 9929 -29864 9935 -29236
rect 9615 -29890 9935 -29864
rect 10615 -29236 10935 -29210
rect 10615 -29864 10621 -29236
rect 10929 -29864 10935 -29236
rect 10615 -29890 10935 -29864
rect 11615 -29236 11935 -29210
rect 11615 -29864 11621 -29236
rect 11929 -29864 11935 -29236
rect 11615 -29890 11935 -29864
rect 12615 -29236 12935 -29210
rect 12615 -29864 12621 -29236
rect 12929 -29864 12935 -29236
rect 12615 -29890 12935 -29864
rect 13615 -29236 13935 -29210
rect 13615 -29864 13621 -29236
rect 13929 -29864 13935 -29236
rect 13615 -29890 13935 -29864
rect 14615 -29236 14935 -29210
rect 14615 -29864 14621 -29236
rect 14929 -29864 14935 -29236
rect 14615 -29890 14935 -29864
rect 15615 -29236 15935 -29210
rect 15615 -29864 15621 -29236
rect 15929 -29864 15935 -29236
rect 15615 -29890 15935 -29864
rect 16615 -29236 16935 -29210
rect 16615 -29864 16621 -29236
rect 16929 -29864 16935 -29236
rect 16615 -29890 16935 -29864
rect 17615 -29236 17935 -29210
rect 17615 -29864 17621 -29236
rect 17929 -29864 17935 -29236
rect 17615 -29890 17935 -29864
rect 18615 -29236 18935 -29210
rect 18615 -29864 18621 -29236
rect 18929 -29864 18935 -29236
rect 18615 -29890 18935 -29864
rect 19615 -29236 19935 -29210
rect 19615 -29864 19621 -29236
rect 19929 -29864 19935 -29236
rect 19615 -29890 19935 -29864
rect 20615 -29236 20935 -29210
rect 20615 -29864 20621 -29236
rect 20929 -29864 20935 -29236
rect 20615 -29890 20935 -29864
rect 21615 -29236 21935 -29210
rect 21615 -29864 21621 -29236
rect 21929 -29864 21935 -29236
rect 21615 -29890 21935 -29864
rect 22615 -29236 22935 -29210
rect 22615 -29864 22621 -29236
rect 22929 -29864 22935 -29236
rect 22615 -29890 22935 -29864
rect 23615 -29236 23935 -29210
rect 23615 -29864 23621 -29236
rect 23929 -29864 23935 -29236
rect 23615 -29890 23935 -29864
rect 24615 -29236 24935 -29210
rect 24615 -29864 24621 -29236
rect 24929 -29864 24935 -29236
rect 24615 -29890 24935 -29864
rect 25615 -29236 25935 -29210
rect 25615 -29864 25621 -29236
rect 25929 -29864 25935 -29236
rect 25615 -29890 25935 -29864
rect 26615 -29236 26935 -29210
rect 26615 -29864 26621 -29236
rect 26929 -29864 26935 -29236
rect 26615 -29890 26935 -29864
rect 27615 -29236 27935 -29210
rect 27615 -29864 27621 -29236
rect 27929 -29864 27935 -29236
rect 27615 -29890 27935 -29864
rect 28615 -29236 28935 -29210
rect 28615 -29864 28621 -29236
rect 28929 -29864 28935 -29236
rect 28615 -29890 28935 -29864
rect 29615 -29236 29935 -29210
rect 29615 -29864 29621 -29236
rect 29929 -29864 29935 -29236
rect 29615 -29890 29935 -29864
rect 30615 -29236 30935 -29210
rect 30615 -29864 30621 -29236
rect 30929 -29864 30935 -29236
rect 30615 -29890 30935 -29864
rect 31615 -29236 31935 -29210
rect 31615 -29864 31621 -29236
rect 31929 -29864 31935 -29236
rect 31615 -29890 31935 -29864
rect 32615 -29236 32935 -29210
rect 32615 -29864 32621 -29236
rect 32929 -29864 32935 -29236
rect 32615 -29890 32935 -29864
rect 33615 -29236 33935 -29210
rect 33615 -29864 33621 -29236
rect 33929 -29864 33935 -29236
rect 33615 -29890 33935 -29864
rect -74825 -29896 -48825 -29890
rect -74825 -30204 -74819 -29896
rect -74511 -29928 -74139 -29896
rect -74511 -30172 -74447 -29928
rect -74203 -30172 -74139 -29928
rect -74511 -30204 -74139 -30172
rect -73511 -29928 -73139 -29896
rect -73511 -30172 -73447 -29928
rect -73203 -30172 -73139 -29928
rect -73511 -30204 -73139 -30172
rect -72511 -29928 -72139 -29896
rect -72511 -30172 -72447 -29928
rect -72203 -30172 -72139 -29928
rect -72511 -30204 -72139 -30172
rect -71511 -29928 -71139 -29896
rect -71511 -30172 -71447 -29928
rect -71203 -30172 -71139 -29928
rect -71511 -30204 -71139 -30172
rect -70511 -29928 -70139 -29896
rect -70511 -30172 -70447 -29928
rect -70203 -30172 -70139 -29928
rect -70511 -30204 -70139 -30172
rect -69511 -29928 -69139 -29896
rect -69511 -30172 -69447 -29928
rect -69203 -30172 -69139 -29928
rect -69511 -30204 -69139 -30172
rect -68511 -29928 -68139 -29896
rect -68511 -30172 -68447 -29928
rect -68203 -30172 -68139 -29928
rect -68511 -30204 -68139 -30172
rect -67511 -29928 -67139 -29896
rect -67511 -30172 -67447 -29928
rect -67203 -30172 -67139 -29928
rect -67511 -30204 -67139 -30172
rect -66511 -29928 -66139 -29896
rect -66511 -30172 -66447 -29928
rect -66203 -30172 -66139 -29928
rect -66511 -30204 -66139 -30172
rect -65511 -29928 -65139 -29896
rect -65511 -30172 -65447 -29928
rect -65203 -30172 -65139 -29928
rect -65511 -30204 -65139 -30172
rect -64511 -29928 -64139 -29896
rect -64511 -30172 -64447 -29928
rect -64203 -30172 -64139 -29928
rect -64511 -30204 -64139 -30172
rect -63511 -29928 -63139 -29896
rect -63511 -30172 -63447 -29928
rect -63203 -30172 -63139 -29928
rect -63511 -30204 -63139 -30172
rect -62511 -29928 -62139 -29896
rect -62511 -30172 -62447 -29928
rect -62203 -30172 -62139 -29928
rect -62511 -30204 -62139 -30172
rect -61511 -29928 -61139 -29896
rect -61511 -30172 -61447 -29928
rect -61203 -30172 -61139 -29928
rect -61511 -30204 -61139 -30172
rect -60511 -29928 -60139 -29896
rect -60511 -30172 -60447 -29928
rect -60203 -30172 -60139 -29928
rect -60511 -30204 -60139 -30172
rect -59511 -29928 -59139 -29896
rect -59511 -30172 -59447 -29928
rect -59203 -30172 -59139 -29928
rect -59511 -30204 -59139 -30172
rect -58511 -29928 -58139 -29896
rect -58511 -30172 -58447 -29928
rect -58203 -30172 -58139 -29928
rect -58511 -30204 -58139 -30172
rect -57511 -29928 -57139 -29896
rect -57511 -30172 -57447 -29928
rect -57203 -30172 -57139 -29928
rect -57511 -30204 -57139 -30172
rect -56511 -29928 -56139 -29896
rect -56511 -30172 -56447 -29928
rect -56203 -30172 -56139 -29928
rect -56511 -30204 -56139 -30172
rect -55511 -29928 -55139 -29896
rect -55511 -30172 -55447 -29928
rect -55203 -30172 -55139 -29928
rect -55511 -30204 -55139 -30172
rect -54511 -29928 -54139 -29896
rect -54511 -30172 -54447 -29928
rect -54203 -30172 -54139 -29928
rect -54511 -30204 -54139 -30172
rect -53511 -29928 -53139 -29896
rect -53511 -30172 -53447 -29928
rect -53203 -30172 -53139 -29928
rect -53511 -30204 -53139 -30172
rect -52511 -29928 -52139 -29896
rect -52511 -30172 -52447 -29928
rect -52203 -30172 -52139 -29928
rect -52511 -30204 -52139 -30172
rect -51511 -29928 -51139 -29896
rect -51511 -30172 -51447 -29928
rect -51203 -30172 -51139 -29928
rect -51511 -30204 -51139 -30172
rect -50511 -29928 -50139 -29896
rect -50511 -30172 -50447 -29928
rect -50203 -30172 -50139 -29928
rect -50511 -30204 -50139 -30172
rect -49511 -29928 -49139 -29896
rect -49511 -30172 -49447 -29928
rect -49203 -30172 -49139 -29928
rect -49511 -30204 -49139 -30172
rect -48831 -30204 -48825 -29896
rect -74825 -30210 -48825 -30204
rect 8275 -29896 34275 -29890
rect 8275 -30204 8281 -29896
rect 8589 -29928 8961 -29896
rect 8589 -30172 8653 -29928
rect 8897 -30172 8961 -29928
rect 8589 -30204 8961 -30172
rect 9589 -29928 9961 -29896
rect 9589 -30172 9653 -29928
rect 9897 -30172 9961 -29928
rect 9589 -30204 9961 -30172
rect 10589 -29928 10961 -29896
rect 10589 -30172 10653 -29928
rect 10897 -30172 10961 -29928
rect 10589 -30204 10961 -30172
rect 11589 -29928 11961 -29896
rect 11589 -30172 11653 -29928
rect 11897 -30172 11961 -29928
rect 11589 -30204 11961 -30172
rect 12589 -29928 12961 -29896
rect 12589 -30172 12653 -29928
rect 12897 -30172 12961 -29928
rect 12589 -30204 12961 -30172
rect 13589 -29928 13961 -29896
rect 13589 -30172 13653 -29928
rect 13897 -30172 13961 -29928
rect 13589 -30204 13961 -30172
rect 14589 -29928 14961 -29896
rect 14589 -30172 14653 -29928
rect 14897 -30172 14961 -29928
rect 14589 -30204 14961 -30172
rect 15589 -29928 15961 -29896
rect 15589 -30172 15653 -29928
rect 15897 -30172 15961 -29928
rect 15589 -30204 15961 -30172
rect 16589 -29928 16961 -29896
rect 16589 -30172 16653 -29928
rect 16897 -30172 16961 -29928
rect 16589 -30204 16961 -30172
rect 17589 -29928 17961 -29896
rect 17589 -30172 17653 -29928
rect 17897 -30172 17961 -29928
rect 17589 -30204 17961 -30172
rect 18589 -29928 18961 -29896
rect 18589 -30172 18653 -29928
rect 18897 -30172 18961 -29928
rect 18589 -30204 18961 -30172
rect 19589 -29928 19961 -29896
rect 19589 -30172 19653 -29928
rect 19897 -30172 19961 -29928
rect 19589 -30204 19961 -30172
rect 20589 -29928 20961 -29896
rect 20589 -30172 20653 -29928
rect 20897 -30172 20961 -29928
rect 20589 -30204 20961 -30172
rect 21589 -29928 21961 -29896
rect 21589 -30172 21653 -29928
rect 21897 -30172 21961 -29928
rect 21589 -30204 21961 -30172
rect 22589 -29928 22961 -29896
rect 22589 -30172 22653 -29928
rect 22897 -30172 22961 -29928
rect 22589 -30204 22961 -30172
rect 23589 -29928 23961 -29896
rect 23589 -30172 23653 -29928
rect 23897 -30172 23961 -29928
rect 23589 -30204 23961 -30172
rect 24589 -29928 24961 -29896
rect 24589 -30172 24653 -29928
rect 24897 -30172 24961 -29928
rect 24589 -30204 24961 -30172
rect 25589 -29928 25961 -29896
rect 25589 -30172 25653 -29928
rect 25897 -30172 25961 -29928
rect 25589 -30204 25961 -30172
rect 26589 -29928 26961 -29896
rect 26589 -30172 26653 -29928
rect 26897 -30172 26961 -29928
rect 26589 -30204 26961 -30172
rect 27589 -29928 27961 -29896
rect 27589 -30172 27653 -29928
rect 27897 -30172 27961 -29928
rect 27589 -30204 27961 -30172
rect 28589 -29928 28961 -29896
rect 28589 -30172 28653 -29928
rect 28897 -30172 28961 -29928
rect 28589 -30204 28961 -30172
rect 29589 -29928 29961 -29896
rect 29589 -30172 29653 -29928
rect 29897 -30172 29961 -29928
rect 29589 -30204 29961 -30172
rect 30589 -29928 30961 -29896
rect 30589 -30172 30653 -29928
rect 30897 -30172 30961 -29928
rect 30589 -30204 30961 -30172
rect 31589 -29928 31961 -29896
rect 31589 -30172 31653 -29928
rect 31897 -30172 31961 -29928
rect 31589 -30204 31961 -30172
rect 32589 -29928 32961 -29896
rect 32589 -30172 32653 -29928
rect 32897 -30172 32961 -29928
rect 32589 -30204 32961 -30172
rect 33589 -29928 33961 -29896
rect 33589 -30172 33653 -29928
rect 33897 -30172 33961 -29928
rect 33589 -30204 33961 -30172
rect 34269 -30204 34275 -29896
rect 8275 -30210 34275 -30204
rect -74485 -30236 -74165 -30210
rect -74485 -30864 -74479 -30236
rect -74171 -30864 -74165 -30236
rect -74485 -30890 -74165 -30864
rect -73485 -30236 -73165 -30210
rect -73485 -30864 -73479 -30236
rect -73171 -30864 -73165 -30236
rect -73485 -30890 -73165 -30864
rect -72485 -30236 -72165 -30210
rect -72485 -30864 -72479 -30236
rect -72171 -30864 -72165 -30236
rect -72485 -30890 -72165 -30864
rect -71485 -30236 -71165 -30210
rect -71485 -30864 -71479 -30236
rect -71171 -30864 -71165 -30236
rect -71485 -30890 -71165 -30864
rect -70485 -30236 -70165 -30210
rect -70485 -30864 -70479 -30236
rect -70171 -30864 -70165 -30236
rect -70485 -30890 -70165 -30864
rect -69485 -30236 -69165 -30210
rect -69485 -30864 -69479 -30236
rect -69171 -30864 -69165 -30236
rect -69485 -30890 -69165 -30864
rect -68485 -30236 -68165 -30210
rect -68485 -30864 -68479 -30236
rect -68171 -30864 -68165 -30236
rect -68485 -30890 -68165 -30864
rect -67485 -30236 -67165 -30210
rect -67485 -30864 -67479 -30236
rect -67171 -30864 -67165 -30236
rect -67485 -30890 -67165 -30864
rect -66485 -30236 -66165 -30210
rect -66485 -30864 -66479 -30236
rect -66171 -30864 -66165 -30236
rect -66485 -30890 -66165 -30864
rect -65485 -30236 -65165 -30210
rect -65485 -30864 -65479 -30236
rect -65171 -30864 -65165 -30236
rect -65485 -30890 -65165 -30864
rect -64485 -30236 -64165 -30210
rect -64485 -30864 -64479 -30236
rect -64171 -30864 -64165 -30236
rect -64485 -30890 -64165 -30864
rect -63485 -30236 -63165 -30210
rect -63485 -30864 -63479 -30236
rect -63171 -30864 -63165 -30236
rect -63485 -30890 -63165 -30864
rect -62485 -30236 -62165 -30210
rect -62485 -30864 -62479 -30236
rect -62171 -30864 -62165 -30236
rect -62485 -30890 -62165 -30864
rect -61485 -30236 -61165 -30210
rect -61485 -30864 -61479 -30236
rect -61171 -30864 -61165 -30236
rect -61485 -30890 -61165 -30864
rect -60485 -30236 -60165 -30210
rect -60485 -30864 -60479 -30236
rect -60171 -30864 -60165 -30236
rect -60485 -30890 -60165 -30864
rect -59485 -30236 -59165 -30210
rect -59485 -30864 -59479 -30236
rect -59171 -30864 -59165 -30236
rect -59485 -30890 -59165 -30864
rect -58485 -30236 -58165 -30210
rect -58485 -30864 -58479 -30236
rect -58171 -30864 -58165 -30236
rect -58485 -30890 -58165 -30864
rect -57485 -30236 -57165 -30210
rect -57485 -30864 -57479 -30236
rect -57171 -30864 -57165 -30236
rect -57485 -30890 -57165 -30864
rect -56485 -30236 -56165 -30210
rect -56485 -30864 -56479 -30236
rect -56171 -30864 -56165 -30236
rect -56485 -30890 -56165 -30864
rect -55485 -30236 -55165 -30210
rect -55485 -30864 -55479 -30236
rect -55171 -30864 -55165 -30236
rect -55485 -30890 -55165 -30864
rect -54485 -30236 -54165 -30210
rect -54485 -30864 -54479 -30236
rect -54171 -30864 -54165 -30236
rect -54485 -30890 -54165 -30864
rect -53485 -30236 -53165 -30210
rect -53485 -30864 -53479 -30236
rect -53171 -30864 -53165 -30236
rect -53485 -30890 -53165 -30864
rect -52485 -30236 -52165 -30210
rect -52485 -30864 -52479 -30236
rect -52171 -30864 -52165 -30236
rect -52485 -30890 -52165 -30864
rect -51485 -30236 -51165 -30210
rect -51485 -30864 -51479 -30236
rect -51171 -30864 -51165 -30236
rect -51485 -30890 -51165 -30864
rect -50485 -30236 -50165 -30210
rect -50485 -30864 -50479 -30236
rect -50171 -30864 -50165 -30236
rect -50485 -30890 -50165 -30864
rect -49485 -30236 -49165 -30210
rect -49485 -30864 -49479 -30236
rect -49171 -30864 -49165 -30236
rect -49485 -30890 -49165 -30864
rect 8615 -30236 8935 -30210
rect 8615 -30864 8621 -30236
rect 8929 -30864 8935 -30236
rect 8615 -30890 8935 -30864
rect 9615 -30236 9935 -30210
rect 9615 -30864 9621 -30236
rect 9929 -30864 9935 -30236
rect 9615 -30890 9935 -30864
rect 10615 -30236 10935 -30210
rect 10615 -30864 10621 -30236
rect 10929 -30864 10935 -30236
rect 10615 -30890 10935 -30864
rect 11615 -30236 11935 -30210
rect 11615 -30864 11621 -30236
rect 11929 -30864 11935 -30236
rect 11615 -30890 11935 -30864
rect 12615 -30236 12935 -30210
rect 12615 -30864 12621 -30236
rect 12929 -30864 12935 -30236
rect 12615 -30890 12935 -30864
rect 13615 -30236 13935 -30210
rect 13615 -30864 13621 -30236
rect 13929 -30864 13935 -30236
rect 13615 -30890 13935 -30864
rect 14615 -30236 14935 -30210
rect 14615 -30864 14621 -30236
rect 14929 -30864 14935 -30236
rect 14615 -30890 14935 -30864
rect 15615 -30236 15935 -30210
rect 15615 -30864 15621 -30236
rect 15929 -30864 15935 -30236
rect 15615 -30890 15935 -30864
rect 16615 -30236 16935 -30210
rect 16615 -30864 16621 -30236
rect 16929 -30864 16935 -30236
rect 16615 -30890 16935 -30864
rect 17615 -30236 17935 -30210
rect 17615 -30864 17621 -30236
rect 17929 -30864 17935 -30236
rect 17615 -30890 17935 -30864
rect 18615 -30236 18935 -30210
rect 18615 -30864 18621 -30236
rect 18929 -30864 18935 -30236
rect 18615 -30890 18935 -30864
rect 19615 -30236 19935 -30210
rect 19615 -30864 19621 -30236
rect 19929 -30864 19935 -30236
rect 19615 -30890 19935 -30864
rect 20615 -30236 20935 -30210
rect 20615 -30864 20621 -30236
rect 20929 -30864 20935 -30236
rect 20615 -30890 20935 -30864
rect 21615 -30236 21935 -30210
rect 21615 -30864 21621 -30236
rect 21929 -30864 21935 -30236
rect 21615 -30890 21935 -30864
rect 22615 -30236 22935 -30210
rect 22615 -30864 22621 -30236
rect 22929 -30864 22935 -30236
rect 22615 -30890 22935 -30864
rect 23615 -30236 23935 -30210
rect 23615 -30864 23621 -30236
rect 23929 -30864 23935 -30236
rect 23615 -30890 23935 -30864
rect 24615 -30236 24935 -30210
rect 24615 -30864 24621 -30236
rect 24929 -30864 24935 -30236
rect 24615 -30890 24935 -30864
rect 25615 -30236 25935 -30210
rect 25615 -30864 25621 -30236
rect 25929 -30864 25935 -30236
rect 25615 -30890 25935 -30864
rect 26615 -30236 26935 -30210
rect 26615 -30864 26621 -30236
rect 26929 -30864 26935 -30236
rect 26615 -30890 26935 -30864
rect 27615 -30236 27935 -30210
rect 27615 -30864 27621 -30236
rect 27929 -30864 27935 -30236
rect 27615 -30890 27935 -30864
rect 28615 -30236 28935 -30210
rect 28615 -30864 28621 -30236
rect 28929 -30864 28935 -30236
rect 28615 -30890 28935 -30864
rect 29615 -30236 29935 -30210
rect 29615 -30864 29621 -30236
rect 29929 -30864 29935 -30236
rect 29615 -30890 29935 -30864
rect 30615 -30236 30935 -30210
rect 30615 -30864 30621 -30236
rect 30929 -30864 30935 -30236
rect 30615 -30890 30935 -30864
rect 31615 -30236 31935 -30210
rect 31615 -30864 31621 -30236
rect 31929 -30864 31935 -30236
rect 31615 -30890 31935 -30864
rect 32615 -30236 32935 -30210
rect 32615 -30864 32621 -30236
rect 32929 -30864 32935 -30236
rect 32615 -30890 32935 -30864
rect 33615 -30236 33935 -30210
rect 33615 -30864 33621 -30236
rect 33929 -30864 33935 -30236
rect 33615 -30890 33935 -30864
rect -74825 -30896 -48825 -30890
rect -74825 -31204 -74819 -30896
rect -74511 -30928 -74139 -30896
rect -74511 -31172 -74447 -30928
rect -74203 -31172 -74139 -30928
rect -74511 -31204 -74139 -31172
rect -73511 -30928 -73139 -30896
rect -73511 -31172 -73447 -30928
rect -73203 -31172 -73139 -30928
rect -73511 -31204 -73139 -31172
rect -72511 -30928 -72139 -30896
rect -72511 -31172 -72447 -30928
rect -72203 -31172 -72139 -30928
rect -72511 -31204 -72139 -31172
rect -71511 -30928 -71139 -30896
rect -71511 -31172 -71447 -30928
rect -71203 -31172 -71139 -30928
rect -71511 -31204 -71139 -31172
rect -70511 -30928 -70139 -30896
rect -70511 -31172 -70447 -30928
rect -70203 -31172 -70139 -30928
rect -70511 -31204 -70139 -31172
rect -69511 -30928 -69139 -30896
rect -69511 -31172 -69447 -30928
rect -69203 -31172 -69139 -30928
rect -69511 -31204 -69139 -31172
rect -68511 -30928 -68139 -30896
rect -68511 -31172 -68447 -30928
rect -68203 -31172 -68139 -30928
rect -68511 -31204 -68139 -31172
rect -67511 -30928 -67139 -30896
rect -67511 -31172 -67447 -30928
rect -67203 -31172 -67139 -30928
rect -67511 -31204 -67139 -31172
rect -66511 -30928 -66139 -30896
rect -66511 -31172 -66447 -30928
rect -66203 -31172 -66139 -30928
rect -66511 -31204 -66139 -31172
rect -65511 -30928 -65139 -30896
rect -65511 -31172 -65447 -30928
rect -65203 -31172 -65139 -30928
rect -65511 -31204 -65139 -31172
rect -64511 -30928 -64139 -30896
rect -64511 -31172 -64447 -30928
rect -64203 -31172 -64139 -30928
rect -64511 -31204 -64139 -31172
rect -63511 -30928 -63139 -30896
rect -63511 -31172 -63447 -30928
rect -63203 -31172 -63139 -30928
rect -63511 -31204 -63139 -31172
rect -62511 -30928 -62139 -30896
rect -62511 -31172 -62447 -30928
rect -62203 -31172 -62139 -30928
rect -62511 -31204 -62139 -31172
rect -61511 -30928 -61139 -30896
rect -61511 -31172 -61447 -30928
rect -61203 -31172 -61139 -30928
rect -61511 -31204 -61139 -31172
rect -60511 -30928 -60139 -30896
rect -60511 -31172 -60447 -30928
rect -60203 -31172 -60139 -30928
rect -60511 -31204 -60139 -31172
rect -59511 -30928 -59139 -30896
rect -59511 -31172 -59447 -30928
rect -59203 -31172 -59139 -30928
rect -59511 -31204 -59139 -31172
rect -58511 -30928 -58139 -30896
rect -58511 -31172 -58447 -30928
rect -58203 -31172 -58139 -30928
rect -58511 -31204 -58139 -31172
rect -57511 -30928 -57139 -30896
rect -57511 -31172 -57447 -30928
rect -57203 -31172 -57139 -30928
rect -57511 -31204 -57139 -31172
rect -56511 -30928 -56139 -30896
rect -56511 -31172 -56447 -30928
rect -56203 -31172 -56139 -30928
rect -56511 -31204 -56139 -31172
rect -55511 -30928 -55139 -30896
rect -55511 -31172 -55447 -30928
rect -55203 -31172 -55139 -30928
rect -55511 -31204 -55139 -31172
rect -54511 -30928 -54139 -30896
rect -54511 -31172 -54447 -30928
rect -54203 -31172 -54139 -30928
rect -54511 -31204 -54139 -31172
rect -53511 -30928 -53139 -30896
rect -53511 -31172 -53447 -30928
rect -53203 -31172 -53139 -30928
rect -53511 -31204 -53139 -31172
rect -52511 -30928 -52139 -30896
rect -52511 -31172 -52447 -30928
rect -52203 -31172 -52139 -30928
rect -52511 -31204 -52139 -31172
rect -51511 -30928 -51139 -30896
rect -51511 -31172 -51447 -30928
rect -51203 -31172 -51139 -30928
rect -51511 -31204 -51139 -31172
rect -50511 -30928 -50139 -30896
rect -50511 -31172 -50447 -30928
rect -50203 -31172 -50139 -30928
rect -50511 -31204 -50139 -31172
rect -49511 -30928 -49139 -30896
rect -49511 -31172 -49447 -30928
rect -49203 -31172 -49139 -30928
rect -49511 -31204 -49139 -31172
rect -48831 -31204 -48825 -30896
rect -74825 -31210 -48825 -31204
rect 8275 -30896 34275 -30890
rect 8275 -31204 8281 -30896
rect 8589 -30928 8961 -30896
rect 8589 -31172 8653 -30928
rect 8897 -31172 8961 -30928
rect 8589 -31204 8961 -31172
rect 9589 -30928 9961 -30896
rect 9589 -31172 9653 -30928
rect 9897 -31172 9961 -30928
rect 9589 -31204 9961 -31172
rect 10589 -30928 10961 -30896
rect 10589 -31172 10653 -30928
rect 10897 -31172 10961 -30928
rect 10589 -31204 10961 -31172
rect 11589 -30928 11961 -30896
rect 11589 -31172 11653 -30928
rect 11897 -31172 11961 -30928
rect 11589 -31204 11961 -31172
rect 12589 -30928 12961 -30896
rect 12589 -31172 12653 -30928
rect 12897 -31172 12961 -30928
rect 12589 -31204 12961 -31172
rect 13589 -30928 13961 -30896
rect 13589 -31172 13653 -30928
rect 13897 -31172 13961 -30928
rect 13589 -31204 13961 -31172
rect 14589 -30928 14961 -30896
rect 14589 -31172 14653 -30928
rect 14897 -31172 14961 -30928
rect 14589 -31204 14961 -31172
rect 15589 -30928 15961 -30896
rect 15589 -31172 15653 -30928
rect 15897 -31172 15961 -30928
rect 15589 -31204 15961 -31172
rect 16589 -30928 16961 -30896
rect 16589 -31172 16653 -30928
rect 16897 -31172 16961 -30928
rect 16589 -31204 16961 -31172
rect 17589 -30928 17961 -30896
rect 17589 -31172 17653 -30928
rect 17897 -31172 17961 -30928
rect 17589 -31204 17961 -31172
rect 18589 -30928 18961 -30896
rect 18589 -31172 18653 -30928
rect 18897 -31172 18961 -30928
rect 18589 -31204 18961 -31172
rect 19589 -30928 19961 -30896
rect 19589 -31172 19653 -30928
rect 19897 -31172 19961 -30928
rect 19589 -31204 19961 -31172
rect 20589 -30928 20961 -30896
rect 20589 -31172 20653 -30928
rect 20897 -31172 20961 -30928
rect 20589 -31204 20961 -31172
rect 21589 -30928 21961 -30896
rect 21589 -31172 21653 -30928
rect 21897 -31172 21961 -30928
rect 21589 -31204 21961 -31172
rect 22589 -30928 22961 -30896
rect 22589 -31172 22653 -30928
rect 22897 -31172 22961 -30928
rect 22589 -31204 22961 -31172
rect 23589 -30928 23961 -30896
rect 23589 -31172 23653 -30928
rect 23897 -31172 23961 -30928
rect 23589 -31204 23961 -31172
rect 24589 -30928 24961 -30896
rect 24589 -31172 24653 -30928
rect 24897 -31172 24961 -30928
rect 24589 -31204 24961 -31172
rect 25589 -30928 25961 -30896
rect 25589 -31172 25653 -30928
rect 25897 -31172 25961 -30928
rect 25589 -31204 25961 -31172
rect 26589 -30928 26961 -30896
rect 26589 -31172 26653 -30928
rect 26897 -31172 26961 -30928
rect 26589 -31204 26961 -31172
rect 27589 -30928 27961 -30896
rect 27589 -31172 27653 -30928
rect 27897 -31172 27961 -30928
rect 27589 -31204 27961 -31172
rect 28589 -30928 28961 -30896
rect 28589 -31172 28653 -30928
rect 28897 -31172 28961 -30928
rect 28589 -31204 28961 -31172
rect 29589 -30928 29961 -30896
rect 29589 -31172 29653 -30928
rect 29897 -31172 29961 -30928
rect 29589 -31204 29961 -31172
rect 30589 -30928 30961 -30896
rect 30589 -31172 30653 -30928
rect 30897 -31172 30961 -30928
rect 30589 -31204 30961 -31172
rect 31589 -30928 31961 -30896
rect 31589 -31172 31653 -30928
rect 31897 -31172 31961 -30928
rect 31589 -31204 31961 -31172
rect 32589 -30928 32961 -30896
rect 32589 -31172 32653 -30928
rect 32897 -31172 32961 -30928
rect 32589 -31204 32961 -31172
rect 33589 -30928 33961 -30896
rect 33589 -31172 33653 -30928
rect 33897 -31172 33961 -30928
rect 33589 -31204 33961 -31172
rect 34269 -31204 34275 -30896
rect 8275 -31210 34275 -31204
rect -74485 -31236 -74165 -31210
rect -74485 -31864 -74479 -31236
rect -74171 -31864 -74165 -31236
rect -74485 -31890 -74165 -31864
rect -73485 -31236 -73165 -31210
rect -73485 -31864 -73479 -31236
rect -73171 -31864 -73165 -31236
rect -73485 -31890 -73165 -31864
rect -72485 -31236 -72165 -31210
rect -72485 -31864 -72479 -31236
rect -72171 -31864 -72165 -31236
rect -72485 -31890 -72165 -31864
rect -71485 -31236 -71165 -31210
rect -71485 -31864 -71479 -31236
rect -71171 -31864 -71165 -31236
rect -71485 -31890 -71165 -31864
rect -70485 -31236 -70165 -31210
rect -70485 -31864 -70479 -31236
rect -70171 -31864 -70165 -31236
rect -70485 -31890 -70165 -31864
rect -69485 -31236 -69165 -31210
rect -69485 -31864 -69479 -31236
rect -69171 -31864 -69165 -31236
rect -69485 -31890 -69165 -31864
rect -68485 -31236 -68165 -31210
rect -68485 -31864 -68479 -31236
rect -68171 -31864 -68165 -31236
rect -68485 -31890 -68165 -31864
rect -67485 -31236 -67165 -31210
rect -67485 -31864 -67479 -31236
rect -67171 -31864 -67165 -31236
rect -67485 -31890 -67165 -31864
rect -66485 -31236 -66165 -31210
rect -66485 -31864 -66479 -31236
rect -66171 -31864 -66165 -31236
rect -66485 -31890 -66165 -31864
rect -65485 -31236 -65165 -31210
rect -65485 -31864 -65479 -31236
rect -65171 -31864 -65165 -31236
rect -65485 -31890 -65165 -31864
rect -64485 -31236 -64165 -31210
rect -64485 -31864 -64479 -31236
rect -64171 -31864 -64165 -31236
rect -64485 -31890 -64165 -31864
rect -63485 -31236 -63165 -31210
rect -63485 -31864 -63479 -31236
rect -63171 -31864 -63165 -31236
rect -63485 -31890 -63165 -31864
rect -62485 -31236 -62165 -31210
rect -62485 -31864 -62479 -31236
rect -62171 -31864 -62165 -31236
rect -62485 -31890 -62165 -31864
rect -61485 -31236 -61165 -31210
rect -61485 -31864 -61479 -31236
rect -61171 -31864 -61165 -31236
rect -61485 -31890 -61165 -31864
rect -60485 -31236 -60165 -31210
rect -60485 -31864 -60479 -31236
rect -60171 -31864 -60165 -31236
rect -60485 -31890 -60165 -31864
rect -59485 -31236 -59165 -31210
rect -59485 -31864 -59479 -31236
rect -59171 -31864 -59165 -31236
rect -59485 -31890 -59165 -31864
rect -58485 -31236 -58165 -31210
rect -58485 -31864 -58479 -31236
rect -58171 -31864 -58165 -31236
rect -58485 -31890 -58165 -31864
rect -57485 -31236 -57165 -31210
rect -57485 -31864 -57479 -31236
rect -57171 -31864 -57165 -31236
rect -57485 -31890 -57165 -31864
rect -56485 -31236 -56165 -31210
rect -56485 -31864 -56479 -31236
rect -56171 -31864 -56165 -31236
rect -56485 -31890 -56165 -31864
rect -55485 -31236 -55165 -31210
rect -55485 -31864 -55479 -31236
rect -55171 -31864 -55165 -31236
rect -55485 -31890 -55165 -31864
rect -54485 -31236 -54165 -31210
rect -54485 -31864 -54479 -31236
rect -54171 -31864 -54165 -31236
rect -54485 -31890 -54165 -31864
rect -53485 -31236 -53165 -31210
rect -53485 -31864 -53479 -31236
rect -53171 -31864 -53165 -31236
rect -53485 -31890 -53165 -31864
rect -52485 -31236 -52165 -31210
rect -52485 -31864 -52479 -31236
rect -52171 -31864 -52165 -31236
rect -52485 -31890 -52165 -31864
rect -51485 -31236 -51165 -31210
rect -51485 -31864 -51479 -31236
rect -51171 -31864 -51165 -31236
rect -51485 -31890 -51165 -31864
rect -50485 -31236 -50165 -31210
rect -50485 -31864 -50479 -31236
rect -50171 -31864 -50165 -31236
rect -50485 -31890 -50165 -31864
rect -49485 -31236 -49165 -31210
rect -49485 -31864 -49479 -31236
rect -49171 -31864 -49165 -31236
rect -49485 -31890 -49165 -31864
rect 8615 -31236 8935 -31210
rect 8615 -31864 8621 -31236
rect 8929 -31864 8935 -31236
rect 8615 -31890 8935 -31864
rect 9615 -31236 9935 -31210
rect 9615 -31864 9621 -31236
rect 9929 -31864 9935 -31236
rect 9615 -31890 9935 -31864
rect 10615 -31236 10935 -31210
rect 10615 -31864 10621 -31236
rect 10929 -31864 10935 -31236
rect 10615 -31890 10935 -31864
rect 11615 -31236 11935 -31210
rect 11615 -31864 11621 -31236
rect 11929 -31864 11935 -31236
rect 11615 -31890 11935 -31864
rect 12615 -31236 12935 -31210
rect 12615 -31864 12621 -31236
rect 12929 -31864 12935 -31236
rect 12615 -31890 12935 -31864
rect 13615 -31236 13935 -31210
rect 13615 -31864 13621 -31236
rect 13929 -31864 13935 -31236
rect 13615 -31890 13935 -31864
rect 14615 -31236 14935 -31210
rect 14615 -31864 14621 -31236
rect 14929 -31864 14935 -31236
rect 14615 -31890 14935 -31864
rect 15615 -31236 15935 -31210
rect 15615 -31864 15621 -31236
rect 15929 -31864 15935 -31236
rect 15615 -31890 15935 -31864
rect 16615 -31236 16935 -31210
rect 16615 -31864 16621 -31236
rect 16929 -31864 16935 -31236
rect 16615 -31890 16935 -31864
rect 17615 -31236 17935 -31210
rect 17615 -31864 17621 -31236
rect 17929 -31864 17935 -31236
rect 17615 -31890 17935 -31864
rect 18615 -31236 18935 -31210
rect 18615 -31864 18621 -31236
rect 18929 -31864 18935 -31236
rect 18615 -31890 18935 -31864
rect 19615 -31236 19935 -31210
rect 19615 -31864 19621 -31236
rect 19929 -31864 19935 -31236
rect 19615 -31890 19935 -31864
rect 20615 -31236 20935 -31210
rect 20615 -31864 20621 -31236
rect 20929 -31864 20935 -31236
rect 20615 -31890 20935 -31864
rect 21615 -31236 21935 -31210
rect 21615 -31864 21621 -31236
rect 21929 -31864 21935 -31236
rect 21615 -31890 21935 -31864
rect 22615 -31236 22935 -31210
rect 22615 -31864 22621 -31236
rect 22929 -31864 22935 -31236
rect 22615 -31890 22935 -31864
rect 23615 -31236 23935 -31210
rect 23615 -31864 23621 -31236
rect 23929 -31864 23935 -31236
rect 23615 -31890 23935 -31864
rect 24615 -31236 24935 -31210
rect 24615 -31864 24621 -31236
rect 24929 -31864 24935 -31236
rect 24615 -31890 24935 -31864
rect 25615 -31236 25935 -31210
rect 25615 -31864 25621 -31236
rect 25929 -31864 25935 -31236
rect 25615 -31890 25935 -31864
rect 26615 -31236 26935 -31210
rect 26615 -31864 26621 -31236
rect 26929 -31864 26935 -31236
rect 26615 -31890 26935 -31864
rect 27615 -31236 27935 -31210
rect 27615 -31864 27621 -31236
rect 27929 -31864 27935 -31236
rect 27615 -31890 27935 -31864
rect 28615 -31236 28935 -31210
rect 28615 -31864 28621 -31236
rect 28929 -31864 28935 -31236
rect 28615 -31890 28935 -31864
rect 29615 -31236 29935 -31210
rect 29615 -31864 29621 -31236
rect 29929 -31864 29935 -31236
rect 29615 -31890 29935 -31864
rect 30615 -31236 30935 -31210
rect 30615 -31864 30621 -31236
rect 30929 -31864 30935 -31236
rect 30615 -31890 30935 -31864
rect 31615 -31236 31935 -31210
rect 31615 -31864 31621 -31236
rect 31929 -31864 31935 -31236
rect 31615 -31890 31935 -31864
rect 32615 -31236 32935 -31210
rect 32615 -31864 32621 -31236
rect 32929 -31864 32935 -31236
rect 32615 -31890 32935 -31864
rect 33615 -31236 33935 -31210
rect 33615 -31864 33621 -31236
rect 33929 -31864 33935 -31236
rect 33615 -31890 33935 -31864
rect -74825 -31896 -48825 -31890
rect -74825 -32204 -74819 -31896
rect -74511 -31928 -74139 -31896
rect -74511 -32172 -74447 -31928
rect -74203 -32172 -74139 -31928
rect -74511 -32204 -74139 -32172
rect -73511 -31928 -73139 -31896
rect -73511 -32172 -73447 -31928
rect -73203 -32172 -73139 -31928
rect -73511 -32204 -73139 -32172
rect -72511 -31928 -72139 -31896
rect -72511 -32172 -72447 -31928
rect -72203 -32172 -72139 -31928
rect -72511 -32204 -72139 -32172
rect -71511 -31928 -71139 -31896
rect -71511 -32172 -71447 -31928
rect -71203 -32172 -71139 -31928
rect -71511 -32204 -71139 -32172
rect -70511 -31928 -70139 -31896
rect -70511 -32172 -70447 -31928
rect -70203 -32172 -70139 -31928
rect -70511 -32204 -70139 -32172
rect -69511 -31928 -69139 -31896
rect -69511 -32172 -69447 -31928
rect -69203 -32172 -69139 -31928
rect -69511 -32204 -69139 -32172
rect -68511 -31928 -68139 -31896
rect -68511 -32172 -68447 -31928
rect -68203 -32172 -68139 -31928
rect -68511 -32204 -68139 -32172
rect -67511 -31928 -67139 -31896
rect -67511 -32172 -67447 -31928
rect -67203 -32172 -67139 -31928
rect -67511 -32204 -67139 -32172
rect -66511 -31928 -66139 -31896
rect -66511 -32172 -66447 -31928
rect -66203 -32172 -66139 -31928
rect -66511 -32204 -66139 -32172
rect -65511 -31928 -65139 -31896
rect -65511 -32172 -65447 -31928
rect -65203 -32172 -65139 -31928
rect -65511 -32204 -65139 -32172
rect -64511 -31928 -64139 -31896
rect -64511 -32172 -64447 -31928
rect -64203 -32172 -64139 -31928
rect -64511 -32204 -64139 -32172
rect -63511 -31928 -63139 -31896
rect -63511 -32172 -63447 -31928
rect -63203 -32172 -63139 -31928
rect -63511 -32204 -63139 -32172
rect -62511 -31928 -62139 -31896
rect -62511 -32172 -62447 -31928
rect -62203 -32172 -62139 -31928
rect -62511 -32204 -62139 -32172
rect -61511 -31928 -61139 -31896
rect -61511 -32172 -61447 -31928
rect -61203 -32172 -61139 -31928
rect -61511 -32204 -61139 -32172
rect -60511 -31928 -60139 -31896
rect -60511 -32172 -60447 -31928
rect -60203 -32172 -60139 -31928
rect -60511 -32204 -60139 -32172
rect -59511 -31928 -59139 -31896
rect -59511 -32172 -59447 -31928
rect -59203 -32172 -59139 -31928
rect -59511 -32204 -59139 -32172
rect -58511 -31928 -58139 -31896
rect -58511 -32172 -58447 -31928
rect -58203 -32172 -58139 -31928
rect -58511 -32204 -58139 -32172
rect -57511 -31928 -57139 -31896
rect -57511 -32172 -57447 -31928
rect -57203 -32172 -57139 -31928
rect -57511 -32204 -57139 -32172
rect -56511 -31928 -56139 -31896
rect -56511 -32172 -56447 -31928
rect -56203 -32172 -56139 -31928
rect -56511 -32204 -56139 -32172
rect -55511 -31928 -55139 -31896
rect -55511 -32172 -55447 -31928
rect -55203 -32172 -55139 -31928
rect -55511 -32204 -55139 -32172
rect -54511 -31928 -54139 -31896
rect -54511 -32172 -54447 -31928
rect -54203 -32172 -54139 -31928
rect -54511 -32204 -54139 -32172
rect -53511 -31928 -53139 -31896
rect -53511 -32172 -53447 -31928
rect -53203 -32172 -53139 -31928
rect -53511 -32204 -53139 -32172
rect -52511 -31928 -52139 -31896
rect -52511 -32172 -52447 -31928
rect -52203 -32172 -52139 -31928
rect -52511 -32204 -52139 -32172
rect -51511 -31928 -51139 -31896
rect -51511 -32172 -51447 -31928
rect -51203 -32172 -51139 -31928
rect -51511 -32204 -51139 -32172
rect -50511 -31928 -50139 -31896
rect -50511 -32172 -50447 -31928
rect -50203 -32172 -50139 -31928
rect -50511 -32204 -50139 -32172
rect -49511 -31928 -49139 -31896
rect -49511 -32172 -49447 -31928
rect -49203 -32172 -49139 -31928
rect -49511 -32204 -49139 -32172
rect -48831 -32204 -48825 -31896
rect -74825 -32210 -48825 -32204
rect 8275 -31896 34275 -31890
rect 8275 -32204 8281 -31896
rect 8589 -31928 8961 -31896
rect 8589 -32172 8653 -31928
rect 8897 -32172 8961 -31928
rect 8589 -32204 8961 -32172
rect 9589 -31928 9961 -31896
rect 9589 -32172 9653 -31928
rect 9897 -32172 9961 -31928
rect 9589 -32204 9961 -32172
rect 10589 -31928 10961 -31896
rect 10589 -32172 10653 -31928
rect 10897 -32172 10961 -31928
rect 10589 -32204 10961 -32172
rect 11589 -31928 11961 -31896
rect 11589 -32172 11653 -31928
rect 11897 -32172 11961 -31928
rect 11589 -32204 11961 -32172
rect 12589 -31928 12961 -31896
rect 12589 -32172 12653 -31928
rect 12897 -32172 12961 -31928
rect 12589 -32204 12961 -32172
rect 13589 -31928 13961 -31896
rect 13589 -32172 13653 -31928
rect 13897 -32172 13961 -31928
rect 13589 -32204 13961 -32172
rect 14589 -31928 14961 -31896
rect 14589 -32172 14653 -31928
rect 14897 -32172 14961 -31928
rect 14589 -32204 14961 -32172
rect 15589 -31928 15961 -31896
rect 15589 -32172 15653 -31928
rect 15897 -32172 15961 -31928
rect 15589 -32204 15961 -32172
rect 16589 -31928 16961 -31896
rect 16589 -32172 16653 -31928
rect 16897 -32172 16961 -31928
rect 16589 -32204 16961 -32172
rect 17589 -31928 17961 -31896
rect 17589 -32172 17653 -31928
rect 17897 -32172 17961 -31928
rect 17589 -32204 17961 -32172
rect 18589 -31928 18961 -31896
rect 18589 -32172 18653 -31928
rect 18897 -32172 18961 -31928
rect 18589 -32204 18961 -32172
rect 19589 -31928 19961 -31896
rect 19589 -32172 19653 -31928
rect 19897 -32172 19961 -31928
rect 19589 -32204 19961 -32172
rect 20589 -31928 20961 -31896
rect 20589 -32172 20653 -31928
rect 20897 -32172 20961 -31928
rect 20589 -32204 20961 -32172
rect 21589 -31928 21961 -31896
rect 21589 -32172 21653 -31928
rect 21897 -32172 21961 -31928
rect 21589 -32204 21961 -32172
rect 22589 -31928 22961 -31896
rect 22589 -32172 22653 -31928
rect 22897 -32172 22961 -31928
rect 22589 -32204 22961 -32172
rect 23589 -31928 23961 -31896
rect 23589 -32172 23653 -31928
rect 23897 -32172 23961 -31928
rect 23589 -32204 23961 -32172
rect 24589 -31928 24961 -31896
rect 24589 -32172 24653 -31928
rect 24897 -32172 24961 -31928
rect 24589 -32204 24961 -32172
rect 25589 -31928 25961 -31896
rect 25589 -32172 25653 -31928
rect 25897 -32172 25961 -31928
rect 25589 -32204 25961 -32172
rect 26589 -31928 26961 -31896
rect 26589 -32172 26653 -31928
rect 26897 -32172 26961 -31928
rect 26589 -32204 26961 -32172
rect 27589 -31928 27961 -31896
rect 27589 -32172 27653 -31928
rect 27897 -32172 27961 -31928
rect 27589 -32204 27961 -32172
rect 28589 -31928 28961 -31896
rect 28589 -32172 28653 -31928
rect 28897 -32172 28961 -31928
rect 28589 -32204 28961 -32172
rect 29589 -31928 29961 -31896
rect 29589 -32172 29653 -31928
rect 29897 -32172 29961 -31928
rect 29589 -32204 29961 -32172
rect 30589 -31928 30961 -31896
rect 30589 -32172 30653 -31928
rect 30897 -32172 30961 -31928
rect 30589 -32204 30961 -32172
rect 31589 -31928 31961 -31896
rect 31589 -32172 31653 -31928
rect 31897 -32172 31961 -31928
rect 31589 -32204 31961 -32172
rect 32589 -31928 32961 -31896
rect 32589 -32172 32653 -31928
rect 32897 -32172 32961 -31928
rect 32589 -32204 32961 -32172
rect 33589 -31928 33961 -31896
rect 33589 -32172 33653 -31928
rect 33897 -32172 33961 -31928
rect 33589 -32204 33961 -32172
rect 34269 -32204 34275 -31896
rect 8275 -32210 34275 -32204
rect -74485 -32236 -74165 -32210
rect -74485 -32864 -74479 -32236
rect -74171 -32864 -74165 -32236
rect -74485 -32890 -74165 -32864
rect -73485 -32236 -73165 -32210
rect -73485 -32864 -73479 -32236
rect -73171 -32864 -73165 -32236
rect -73485 -32890 -73165 -32864
rect -72485 -32236 -72165 -32210
rect -72485 -32864 -72479 -32236
rect -72171 -32864 -72165 -32236
rect -72485 -32890 -72165 -32864
rect -71485 -32236 -71165 -32210
rect -71485 -32864 -71479 -32236
rect -71171 -32864 -71165 -32236
rect -71485 -32890 -71165 -32864
rect -70485 -32236 -70165 -32210
rect -70485 -32864 -70479 -32236
rect -70171 -32864 -70165 -32236
rect -70485 -32890 -70165 -32864
rect -69485 -32236 -69165 -32210
rect -69485 -32864 -69479 -32236
rect -69171 -32864 -69165 -32236
rect -69485 -32890 -69165 -32864
rect -68485 -32236 -68165 -32210
rect -68485 -32864 -68479 -32236
rect -68171 -32864 -68165 -32236
rect -68485 -32890 -68165 -32864
rect -67485 -32236 -67165 -32210
rect -67485 -32864 -67479 -32236
rect -67171 -32864 -67165 -32236
rect -67485 -32890 -67165 -32864
rect -66485 -32236 -66165 -32210
rect -66485 -32864 -66479 -32236
rect -66171 -32864 -66165 -32236
rect -66485 -32890 -66165 -32864
rect -65485 -32236 -65165 -32210
rect -65485 -32864 -65479 -32236
rect -65171 -32864 -65165 -32236
rect -65485 -32890 -65165 -32864
rect -64485 -32236 -64165 -32210
rect -64485 -32864 -64479 -32236
rect -64171 -32864 -64165 -32236
rect -64485 -32890 -64165 -32864
rect -63485 -32236 -63165 -32210
rect -63485 -32864 -63479 -32236
rect -63171 -32864 -63165 -32236
rect -63485 -32890 -63165 -32864
rect -62485 -32236 -62165 -32210
rect -62485 -32864 -62479 -32236
rect -62171 -32864 -62165 -32236
rect -62485 -32890 -62165 -32864
rect -61485 -32236 -61165 -32210
rect -61485 -32864 -61479 -32236
rect -61171 -32864 -61165 -32236
rect -61485 -32890 -61165 -32864
rect -60485 -32236 -60165 -32210
rect -60485 -32864 -60479 -32236
rect -60171 -32864 -60165 -32236
rect -60485 -32890 -60165 -32864
rect -59485 -32236 -59165 -32210
rect -59485 -32864 -59479 -32236
rect -59171 -32864 -59165 -32236
rect -59485 -32890 -59165 -32864
rect -58485 -32236 -58165 -32210
rect -58485 -32864 -58479 -32236
rect -58171 -32864 -58165 -32236
rect -58485 -32890 -58165 -32864
rect -57485 -32236 -57165 -32210
rect -57485 -32864 -57479 -32236
rect -57171 -32864 -57165 -32236
rect -57485 -32890 -57165 -32864
rect -56485 -32236 -56165 -32210
rect -56485 -32864 -56479 -32236
rect -56171 -32864 -56165 -32236
rect -56485 -32890 -56165 -32864
rect -55485 -32236 -55165 -32210
rect -55485 -32864 -55479 -32236
rect -55171 -32864 -55165 -32236
rect -55485 -32890 -55165 -32864
rect -54485 -32236 -54165 -32210
rect -54485 -32864 -54479 -32236
rect -54171 -32864 -54165 -32236
rect -54485 -32890 -54165 -32864
rect -53485 -32236 -53165 -32210
rect -53485 -32864 -53479 -32236
rect -53171 -32864 -53165 -32236
rect -53485 -32890 -53165 -32864
rect -52485 -32236 -52165 -32210
rect -52485 -32864 -52479 -32236
rect -52171 -32864 -52165 -32236
rect -52485 -32890 -52165 -32864
rect -51485 -32236 -51165 -32210
rect -51485 -32864 -51479 -32236
rect -51171 -32864 -51165 -32236
rect -51485 -32890 -51165 -32864
rect -50485 -32236 -50165 -32210
rect -50485 -32864 -50479 -32236
rect -50171 -32864 -50165 -32236
rect -50485 -32890 -50165 -32864
rect -49485 -32236 -49165 -32210
rect -49485 -32864 -49479 -32236
rect -49171 -32864 -49165 -32236
rect 8615 -32236 8935 -32210
rect -49485 -32890 -49165 -32864
rect -46275 -32604 -27875 -32550
rect -74825 -32896 -48825 -32890
rect -74825 -33204 -74819 -32896
rect -74511 -32928 -74139 -32896
rect -74511 -33172 -74447 -32928
rect -74203 -33172 -74139 -32928
rect -74511 -33204 -74139 -33172
rect -73511 -32928 -73139 -32896
rect -73511 -33172 -73447 -32928
rect -73203 -33172 -73139 -32928
rect -73511 -33204 -73139 -33172
rect -72511 -32928 -72139 -32896
rect -72511 -33172 -72447 -32928
rect -72203 -33172 -72139 -32928
rect -72511 -33204 -72139 -33172
rect -71511 -32928 -71139 -32896
rect -71511 -33172 -71447 -32928
rect -71203 -33172 -71139 -32928
rect -71511 -33204 -71139 -33172
rect -70511 -32928 -70139 -32896
rect -70511 -33172 -70447 -32928
rect -70203 -33172 -70139 -32928
rect -70511 -33204 -70139 -33172
rect -69511 -32928 -69139 -32896
rect -69511 -33172 -69447 -32928
rect -69203 -33172 -69139 -32928
rect -69511 -33204 -69139 -33172
rect -68511 -32928 -68139 -32896
rect -68511 -33172 -68447 -32928
rect -68203 -33172 -68139 -32928
rect -68511 -33204 -68139 -33172
rect -67511 -32928 -67139 -32896
rect -67511 -33172 -67447 -32928
rect -67203 -33172 -67139 -32928
rect -67511 -33204 -67139 -33172
rect -66511 -32928 -66139 -32896
rect -66511 -33172 -66447 -32928
rect -66203 -33172 -66139 -32928
rect -66511 -33204 -66139 -33172
rect -65511 -32928 -65139 -32896
rect -65511 -33172 -65447 -32928
rect -65203 -33172 -65139 -32928
rect -65511 -33204 -65139 -33172
rect -64511 -32928 -64139 -32896
rect -64511 -33172 -64447 -32928
rect -64203 -33172 -64139 -32928
rect -64511 -33204 -64139 -33172
rect -63511 -32928 -63139 -32896
rect -63511 -33172 -63447 -32928
rect -63203 -33172 -63139 -32928
rect -63511 -33204 -63139 -33172
rect -62511 -32928 -62139 -32896
rect -62511 -33172 -62447 -32928
rect -62203 -33172 -62139 -32928
rect -62511 -33204 -62139 -33172
rect -61511 -32928 -61139 -32896
rect -61511 -33172 -61447 -32928
rect -61203 -33172 -61139 -32928
rect -61511 -33204 -61139 -33172
rect -60511 -32928 -60139 -32896
rect -60511 -33172 -60447 -32928
rect -60203 -33172 -60139 -32928
rect -60511 -33204 -60139 -33172
rect -59511 -32928 -59139 -32896
rect -59511 -33172 -59447 -32928
rect -59203 -33172 -59139 -32928
rect -59511 -33204 -59139 -33172
rect -58511 -32928 -58139 -32896
rect -58511 -33172 -58447 -32928
rect -58203 -33172 -58139 -32928
rect -58511 -33204 -58139 -33172
rect -57511 -32928 -57139 -32896
rect -57511 -33172 -57447 -32928
rect -57203 -33172 -57139 -32928
rect -57511 -33204 -57139 -33172
rect -56511 -32928 -56139 -32896
rect -56511 -33172 -56447 -32928
rect -56203 -33172 -56139 -32928
rect -56511 -33204 -56139 -33172
rect -55511 -32928 -55139 -32896
rect -55511 -33172 -55447 -32928
rect -55203 -33172 -55139 -32928
rect -55511 -33204 -55139 -33172
rect -54511 -32928 -54139 -32896
rect -54511 -33172 -54447 -32928
rect -54203 -33172 -54139 -32928
rect -54511 -33204 -54139 -33172
rect -53511 -32928 -53139 -32896
rect -53511 -33172 -53447 -32928
rect -53203 -33172 -53139 -32928
rect -53511 -33204 -53139 -33172
rect -52511 -32928 -52139 -32896
rect -52511 -33172 -52447 -32928
rect -52203 -33172 -52139 -32928
rect -52511 -33204 -52139 -33172
rect -51511 -32928 -51139 -32896
rect -51511 -33172 -51447 -32928
rect -51203 -33172 -51139 -32928
rect -51511 -33204 -51139 -33172
rect -50511 -32928 -50139 -32896
rect -50511 -33172 -50447 -32928
rect -50203 -33172 -50139 -32928
rect -50511 -33204 -50139 -33172
rect -49511 -32928 -49139 -32896
rect -49511 -33172 -49447 -32928
rect -49203 -33172 -49139 -32928
rect -49511 -33204 -49139 -33172
rect -48831 -33204 -48825 -32896
rect -74825 -33210 -48825 -33204
rect -74485 -33236 -74165 -33210
rect -74485 -33864 -74479 -33236
rect -74171 -33864 -74165 -33236
rect -74485 -33890 -74165 -33864
rect -73485 -33236 -73165 -33210
rect -73485 -33864 -73479 -33236
rect -73171 -33864 -73165 -33236
rect -73485 -33890 -73165 -33864
rect -72485 -33236 -72165 -33210
rect -72485 -33864 -72479 -33236
rect -72171 -33864 -72165 -33236
rect -72485 -33890 -72165 -33864
rect -71485 -33236 -71165 -33210
rect -71485 -33864 -71479 -33236
rect -71171 -33864 -71165 -33236
rect -71485 -33890 -71165 -33864
rect -70485 -33236 -70165 -33210
rect -70485 -33864 -70479 -33236
rect -70171 -33864 -70165 -33236
rect -70485 -33890 -70165 -33864
rect -69485 -33236 -69165 -33210
rect -69485 -33864 -69479 -33236
rect -69171 -33864 -69165 -33236
rect -69485 -33890 -69165 -33864
rect -68485 -33236 -68165 -33210
rect -68485 -33864 -68479 -33236
rect -68171 -33864 -68165 -33236
rect -68485 -33890 -68165 -33864
rect -67485 -33236 -67165 -33210
rect -67485 -33864 -67479 -33236
rect -67171 -33864 -67165 -33236
rect -67485 -33890 -67165 -33864
rect -66485 -33236 -66165 -33210
rect -66485 -33864 -66479 -33236
rect -66171 -33864 -66165 -33236
rect -66485 -33890 -66165 -33864
rect -65485 -33236 -65165 -33210
rect -65485 -33864 -65479 -33236
rect -65171 -33864 -65165 -33236
rect -65485 -33890 -65165 -33864
rect -64485 -33236 -64165 -33210
rect -64485 -33864 -64479 -33236
rect -64171 -33864 -64165 -33236
rect -64485 -33890 -64165 -33864
rect -63485 -33236 -63165 -33210
rect -63485 -33864 -63479 -33236
rect -63171 -33864 -63165 -33236
rect -63485 -33890 -63165 -33864
rect -62485 -33236 -62165 -33210
rect -62485 -33864 -62479 -33236
rect -62171 -33864 -62165 -33236
rect -62485 -33890 -62165 -33864
rect -61485 -33236 -61165 -33210
rect -61485 -33864 -61479 -33236
rect -61171 -33864 -61165 -33236
rect -61485 -33890 -61165 -33864
rect -60485 -33236 -60165 -33210
rect -60485 -33864 -60479 -33236
rect -60171 -33864 -60165 -33236
rect -60485 -33890 -60165 -33864
rect -59485 -33236 -59165 -33210
rect -59485 -33864 -59479 -33236
rect -59171 -33864 -59165 -33236
rect -59485 -33890 -59165 -33864
rect -58485 -33236 -58165 -33210
rect -58485 -33864 -58479 -33236
rect -58171 -33864 -58165 -33236
rect -58485 -33890 -58165 -33864
rect -57485 -33236 -57165 -33210
rect -57485 -33864 -57479 -33236
rect -57171 -33864 -57165 -33236
rect -57485 -33890 -57165 -33864
rect -56485 -33236 -56165 -33210
rect -56485 -33864 -56479 -33236
rect -56171 -33864 -56165 -33236
rect -56485 -33890 -56165 -33864
rect -55485 -33236 -55165 -33210
rect -55485 -33864 -55479 -33236
rect -55171 -33864 -55165 -33236
rect -55485 -33890 -55165 -33864
rect -54485 -33236 -54165 -33210
rect -54485 -33864 -54479 -33236
rect -54171 -33864 -54165 -33236
rect -54485 -33890 -54165 -33864
rect -53485 -33236 -53165 -33210
rect -53485 -33864 -53479 -33236
rect -53171 -33864 -53165 -33236
rect -53485 -33890 -53165 -33864
rect -52485 -33236 -52165 -33210
rect -52485 -33864 -52479 -33236
rect -52171 -33864 -52165 -33236
rect -52485 -33890 -52165 -33864
rect -51485 -33236 -51165 -33210
rect -51485 -33864 -51479 -33236
rect -51171 -33864 -51165 -33236
rect -51485 -33890 -51165 -33864
rect -50485 -33236 -50165 -33210
rect -50485 -33864 -50479 -33236
rect -50171 -33864 -50165 -33236
rect -50485 -33890 -50165 -33864
rect -49485 -33236 -49165 -33210
rect -49485 -33864 -49479 -33236
rect -49171 -33864 -49165 -33236
rect -49485 -33890 -49165 -33864
rect -74825 -33896 -48825 -33890
rect -74825 -34204 -74819 -33896
rect -74511 -33928 -74139 -33896
rect -74511 -34172 -74447 -33928
rect -74203 -34172 -74139 -33928
rect -74511 -34204 -74139 -34172
rect -73511 -33928 -73139 -33896
rect -73511 -34172 -73447 -33928
rect -73203 -34172 -73139 -33928
rect -73511 -34204 -73139 -34172
rect -72511 -33928 -72139 -33896
rect -72511 -34172 -72447 -33928
rect -72203 -34172 -72139 -33928
rect -72511 -34204 -72139 -34172
rect -71511 -33928 -71139 -33896
rect -71511 -34172 -71447 -33928
rect -71203 -34172 -71139 -33928
rect -71511 -34204 -71139 -34172
rect -70511 -33928 -70139 -33896
rect -70511 -34172 -70447 -33928
rect -70203 -34172 -70139 -33928
rect -70511 -34204 -70139 -34172
rect -69511 -33928 -69139 -33896
rect -69511 -34172 -69447 -33928
rect -69203 -34172 -69139 -33928
rect -69511 -34204 -69139 -34172
rect -68511 -33928 -68139 -33896
rect -68511 -34172 -68447 -33928
rect -68203 -34172 -68139 -33928
rect -68511 -34204 -68139 -34172
rect -67511 -33928 -67139 -33896
rect -67511 -34172 -67447 -33928
rect -67203 -34172 -67139 -33928
rect -67511 -34204 -67139 -34172
rect -66511 -33928 -66139 -33896
rect -66511 -34172 -66447 -33928
rect -66203 -34172 -66139 -33928
rect -66511 -34204 -66139 -34172
rect -65511 -33928 -65139 -33896
rect -65511 -34172 -65447 -33928
rect -65203 -34172 -65139 -33928
rect -65511 -34204 -65139 -34172
rect -64511 -33928 -64139 -33896
rect -64511 -34172 -64447 -33928
rect -64203 -34172 -64139 -33928
rect -64511 -34204 -64139 -34172
rect -63511 -33928 -63139 -33896
rect -63511 -34172 -63447 -33928
rect -63203 -34172 -63139 -33928
rect -63511 -34204 -63139 -34172
rect -62511 -33928 -62139 -33896
rect -62511 -34172 -62447 -33928
rect -62203 -34172 -62139 -33928
rect -62511 -34204 -62139 -34172
rect -61511 -33928 -61139 -33896
rect -61511 -34172 -61447 -33928
rect -61203 -34172 -61139 -33928
rect -61511 -34204 -61139 -34172
rect -60511 -33928 -60139 -33896
rect -60511 -34172 -60447 -33928
rect -60203 -34172 -60139 -33928
rect -60511 -34204 -60139 -34172
rect -59511 -33928 -59139 -33896
rect -59511 -34172 -59447 -33928
rect -59203 -34172 -59139 -33928
rect -59511 -34204 -59139 -34172
rect -58511 -33928 -58139 -33896
rect -58511 -34172 -58447 -33928
rect -58203 -34172 -58139 -33928
rect -58511 -34204 -58139 -34172
rect -57511 -33928 -57139 -33896
rect -57511 -34172 -57447 -33928
rect -57203 -34172 -57139 -33928
rect -57511 -34204 -57139 -34172
rect -56511 -33928 -56139 -33896
rect -56511 -34172 -56447 -33928
rect -56203 -34172 -56139 -33928
rect -56511 -34204 -56139 -34172
rect -55511 -33928 -55139 -33896
rect -55511 -34172 -55447 -33928
rect -55203 -34172 -55139 -33928
rect -55511 -34204 -55139 -34172
rect -54511 -33928 -54139 -33896
rect -54511 -34172 -54447 -33928
rect -54203 -34172 -54139 -33928
rect -54511 -34204 -54139 -34172
rect -53511 -33928 -53139 -33896
rect -53511 -34172 -53447 -33928
rect -53203 -34172 -53139 -33928
rect -53511 -34204 -53139 -34172
rect -52511 -33928 -52139 -33896
rect -52511 -34172 -52447 -33928
rect -52203 -34172 -52139 -33928
rect -52511 -34204 -52139 -34172
rect -51511 -33928 -51139 -33896
rect -51511 -34172 -51447 -33928
rect -51203 -34172 -51139 -33928
rect -51511 -34204 -51139 -34172
rect -50511 -33928 -50139 -33896
rect -50511 -34172 -50447 -33928
rect -50203 -34172 -50139 -33928
rect -50511 -34204 -50139 -34172
rect -49511 -33928 -49139 -33896
rect -49511 -34172 -49447 -33928
rect -49203 -34172 -49139 -33928
rect -49511 -34204 -49139 -34172
rect -48831 -34204 -48825 -33896
rect -74825 -34210 -48825 -34204
rect -74485 -34236 -74165 -34210
rect -74485 -34864 -74479 -34236
rect -74171 -34864 -74165 -34236
rect -74485 -34890 -74165 -34864
rect -73485 -34236 -73165 -34210
rect -73485 -34864 -73479 -34236
rect -73171 -34864 -73165 -34236
rect -73485 -34890 -73165 -34864
rect -72485 -34236 -72165 -34210
rect -72485 -34864 -72479 -34236
rect -72171 -34864 -72165 -34236
rect -72485 -34890 -72165 -34864
rect -71485 -34236 -71165 -34210
rect -71485 -34864 -71479 -34236
rect -71171 -34864 -71165 -34236
rect -71485 -34890 -71165 -34864
rect -70485 -34236 -70165 -34210
rect -70485 -34864 -70479 -34236
rect -70171 -34864 -70165 -34236
rect -70485 -34890 -70165 -34864
rect -69485 -34236 -69165 -34210
rect -69485 -34864 -69479 -34236
rect -69171 -34864 -69165 -34236
rect -69485 -34890 -69165 -34864
rect -68485 -34236 -68165 -34210
rect -68485 -34864 -68479 -34236
rect -68171 -34864 -68165 -34236
rect -68485 -34890 -68165 -34864
rect -67485 -34236 -67165 -34210
rect -67485 -34864 -67479 -34236
rect -67171 -34864 -67165 -34236
rect -67485 -34890 -67165 -34864
rect -66485 -34236 -66165 -34210
rect -66485 -34864 -66479 -34236
rect -66171 -34864 -66165 -34236
rect -66485 -34890 -66165 -34864
rect -65485 -34236 -65165 -34210
rect -65485 -34864 -65479 -34236
rect -65171 -34864 -65165 -34236
rect -65485 -34890 -65165 -34864
rect -64485 -34236 -64165 -34210
rect -64485 -34864 -64479 -34236
rect -64171 -34864 -64165 -34236
rect -64485 -34890 -64165 -34864
rect -63485 -34236 -63165 -34210
rect -63485 -34864 -63479 -34236
rect -63171 -34864 -63165 -34236
rect -63485 -34890 -63165 -34864
rect -62485 -34236 -62165 -34210
rect -62485 -34864 -62479 -34236
rect -62171 -34864 -62165 -34236
rect -62485 -34890 -62165 -34864
rect -61485 -34236 -61165 -34210
rect -61485 -34864 -61479 -34236
rect -61171 -34864 -61165 -34236
rect -61485 -34890 -61165 -34864
rect -60485 -34236 -60165 -34210
rect -60485 -34864 -60479 -34236
rect -60171 -34864 -60165 -34236
rect -60485 -34890 -60165 -34864
rect -59485 -34236 -59165 -34210
rect -59485 -34864 -59479 -34236
rect -59171 -34864 -59165 -34236
rect -59485 -34890 -59165 -34864
rect -58485 -34236 -58165 -34210
rect -58485 -34864 -58479 -34236
rect -58171 -34864 -58165 -34236
rect -58485 -34890 -58165 -34864
rect -57485 -34236 -57165 -34210
rect -57485 -34864 -57479 -34236
rect -57171 -34864 -57165 -34236
rect -57485 -34890 -57165 -34864
rect -56485 -34236 -56165 -34210
rect -56485 -34864 -56479 -34236
rect -56171 -34864 -56165 -34236
rect -56485 -34890 -56165 -34864
rect -55485 -34236 -55165 -34210
rect -55485 -34864 -55479 -34236
rect -55171 -34864 -55165 -34236
rect -55485 -34890 -55165 -34864
rect -54485 -34236 -54165 -34210
rect -54485 -34864 -54479 -34236
rect -54171 -34864 -54165 -34236
rect -54485 -34890 -54165 -34864
rect -53485 -34236 -53165 -34210
rect -53485 -34864 -53479 -34236
rect -53171 -34864 -53165 -34236
rect -53485 -34890 -53165 -34864
rect -52485 -34236 -52165 -34210
rect -52485 -34864 -52479 -34236
rect -52171 -34864 -52165 -34236
rect -52485 -34890 -52165 -34864
rect -51485 -34236 -51165 -34210
rect -51485 -34864 -51479 -34236
rect -51171 -34864 -51165 -34236
rect -51485 -34890 -51165 -34864
rect -50485 -34236 -50165 -34210
rect -50485 -34864 -50479 -34236
rect -50171 -34864 -50165 -34236
rect -50485 -34890 -50165 -34864
rect -49485 -34236 -49165 -34210
rect -49485 -34864 -49479 -34236
rect -49171 -34864 -49165 -34236
rect -49485 -34890 -49165 -34864
rect -74825 -34896 -48825 -34890
rect -74825 -35204 -74819 -34896
rect -74511 -34928 -74139 -34896
rect -74511 -35172 -74447 -34928
rect -74203 -35172 -74139 -34928
rect -74511 -35204 -74139 -35172
rect -73511 -34928 -73139 -34896
rect -73511 -35172 -73447 -34928
rect -73203 -35172 -73139 -34928
rect -73511 -35204 -73139 -35172
rect -72511 -34928 -72139 -34896
rect -72511 -35172 -72447 -34928
rect -72203 -35172 -72139 -34928
rect -72511 -35204 -72139 -35172
rect -71511 -34928 -71139 -34896
rect -71511 -35172 -71447 -34928
rect -71203 -35172 -71139 -34928
rect -71511 -35204 -71139 -35172
rect -70511 -34928 -70139 -34896
rect -70511 -35172 -70447 -34928
rect -70203 -35172 -70139 -34928
rect -70511 -35204 -70139 -35172
rect -69511 -34928 -69139 -34896
rect -69511 -35172 -69447 -34928
rect -69203 -35172 -69139 -34928
rect -69511 -35204 -69139 -35172
rect -68511 -34928 -68139 -34896
rect -68511 -35172 -68447 -34928
rect -68203 -35172 -68139 -34928
rect -68511 -35204 -68139 -35172
rect -67511 -34928 -67139 -34896
rect -67511 -35172 -67447 -34928
rect -67203 -35172 -67139 -34928
rect -67511 -35204 -67139 -35172
rect -66511 -34928 -66139 -34896
rect -66511 -35172 -66447 -34928
rect -66203 -35172 -66139 -34928
rect -66511 -35204 -66139 -35172
rect -65511 -34928 -65139 -34896
rect -65511 -35172 -65447 -34928
rect -65203 -35172 -65139 -34928
rect -65511 -35204 -65139 -35172
rect -64511 -34928 -64139 -34896
rect -64511 -35172 -64447 -34928
rect -64203 -35172 -64139 -34928
rect -64511 -35204 -64139 -35172
rect -63511 -34928 -63139 -34896
rect -63511 -35172 -63447 -34928
rect -63203 -35172 -63139 -34928
rect -63511 -35204 -63139 -35172
rect -62511 -34928 -62139 -34896
rect -62511 -35172 -62447 -34928
rect -62203 -35172 -62139 -34928
rect -62511 -35204 -62139 -35172
rect -61511 -34928 -61139 -34896
rect -61511 -35172 -61447 -34928
rect -61203 -35172 -61139 -34928
rect -61511 -35204 -61139 -35172
rect -60511 -34928 -60139 -34896
rect -60511 -35172 -60447 -34928
rect -60203 -35172 -60139 -34928
rect -60511 -35204 -60139 -35172
rect -59511 -34928 -59139 -34896
rect -59511 -35172 -59447 -34928
rect -59203 -35172 -59139 -34928
rect -59511 -35204 -59139 -35172
rect -58511 -34928 -58139 -34896
rect -58511 -35172 -58447 -34928
rect -58203 -35172 -58139 -34928
rect -58511 -35204 -58139 -35172
rect -57511 -34928 -57139 -34896
rect -57511 -35172 -57447 -34928
rect -57203 -35172 -57139 -34928
rect -57511 -35204 -57139 -35172
rect -56511 -34928 -56139 -34896
rect -56511 -35172 -56447 -34928
rect -56203 -35172 -56139 -34928
rect -56511 -35204 -56139 -35172
rect -55511 -34928 -55139 -34896
rect -55511 -35172 -55447 -34928
rect -55203 -35172 -55139 -34928
rect -55511 -35204 -55139 -35172
rect -54511 -34928 -54139 -34896
rect -54511 -35172 -54447 -34928
rect -54203 -35172 -54139 -34928
rect -54511 -35204 -54139 -35172
rect -53511 -34928 -53139 -34896
rect -53511 -35172 -53447 -34928
rect -53203 -35172 -53139 -34928
rect -53511 -35204 -53139 -35172
rect -52511 -34928 -52139 -34896
rect -52511 -35172 -52447 -34928
rect -52203 -35172 -52139 -34928
rect -52511 -35204 -52139 -35172
rect -51511 -34928 -51139 -34896
rect -51511 -35172 -51447 -34928
rect -51203 -35172 -51139 -34928
rect -51511 -35204 -51139 -35172
rect -50511 -34928 -50139 -34896
rect -50511 -35172 -50447 -34928
rect -50203 -35172 -50139 -34928
rect -50511 -35204 -50139 -35172
rect -49511 -34928 -49139 -34896
rect -49511 -35172 -49447 -34928
rect -49203 -35172 -49139 -34928
rect -49511 -35204 -49139 -35172
rect -48831 -35204 -48825 -34896
rect -74825 -35210 -48825 -35204
rect -74485 -35236 -74165 -35210
rect -74485 -35864 -74479 -35236
rect -74171 -35864 -74165 -35236
rect -74485 -35890 -74165 -35864
rect -73485 -35236 -73165 -35210
rect -73485 -35864 -73479 -35236
rect -73171 -35864 -73165 -35236
rect -73485 -35890 -73165 -35864
rect -72485 -35236 -72165 -35210
rect -72485 -35864 -72479 -35236
rect -72171 -35864 -72165 -35236
rect -72485 -35890 -72165 -35864
rect -71485 -35236 -71165 -35210
rect -71485 -35864 -71479 -35236
rect -71171 -35864 -71165 -35236
rect -71485 -35890 -71165 -35864
rect -70485 -35236 -70165 -35210
rect -70485 -35864 -70479 -35236
rect -70171 -35864 -70165 -35236
rect -70485 -35890 -70165 -35864
rect -69485 -35236 -69165 -35210
rect -69485 -35864 -69479 -35236
rect -69171 -35864 -69165 -35236
rect -69485 -35890 -69165 -35864
rect -68485 -35236 -68165 -35210
rect -68485 -35864 -68479 -35236
rect -68171 -35864 -68165 -35236
rect -68485 -35890 -68165 -35864
rect -67485 -35236 -67165 -35210
rect -67485 -35864 -67479 -35236
rect -67171 -35864 -67165 -35236
rect -67485 -35890 -67165 -35864
rect -66485 -35236 -66165 -35210
rect -66485 -35864 -66479 -35236
rect -66171 -35864 -66165 -35236
rect -66485 -35890 -66165 -35864
rect -65485 -35236 -65165 -35210
rect -65485 -35864 -65479 -35236
rect -65171 -35864 -65165 -35236
rect -65485 -35890 -65165 -35864
rect -64485 -35236 -64165 -35210
rect -64485 -35864 -64479 -35236
rect -64171 -35864 -64165 -35236
rect -64485 -35890 -64165 -35864
rect -63485 -35236 -63165 -35210
rect -63485 -35864 -63479 -35236
rect -63171 -35864 -63165 -35236
rect -63485 -35890 -63165 -35864
rect -62485 -35236 -62165 -35210
rect -62485 -35864 -62479 -35236
rect -62171 -35864 -62165 -35236
rect -62485 -35890 -62165 -35864
rect -61485 -35236 -61165 -35210
rect -61485 -35864 -61479 -35236
rect -61171 -35864 -61165 -35236
rect -61485 -35890 -61165 -35864
rect -60485 -35236 -60165 -35210
rect -60485 -35864 -60479 -35236
rect -60171 -35864 -60165 -35236
rect -60485 -35890 -60165 -35864
rect -59485 -35236 -59165 -35210
rect -59485 -35864 -59479 -35236
rect -59171 -35864 -59165 -35236
rect -59485 -35890 -59165 -35864
rect -58485 -35236 -58165 -35210
rect -58485 -35864 -58479 -35236
rect -58171 -35864 -58165 -35236
rect -58485 -35890 -58165 -35864
rect -57485 -35236 -57165 -35210
rect -57485 -35864 -57479 -35236
rect -57171 -35864 -57165 -35236
rect -57485 -35890 -57165 -35864
rect -56485 -35236 -56165 -35210
rect -56485 -35864 -56479 -35236
rect -56171 -35864 -56165 -35236
rect -56485 -35890 -56165 -35864
rect -55485 -35236 -55165 -35210
rect -55485 -35864 -55479 -35236
rect -55171 -35864 -55165 -35236
rect -55485 -35890 -55165 -35864
rect -54485 -35236 -54165 -35210
rect -54485 -35864 -54479 -35236
rect -54171 -35864 -54165 -35236
rect -54485 -35890 -54165 -35864
rect -53485 -35236 -53165 -35210
rect -53485 -35864 -53479 -35236
rect -53171 -35864 -53165 -35236
rect -53485 -35890 -53165 -35864
rect -52485 -35236 -52165 -35210
rect -52485 -35864 -52479 -35236
rect -52171 -35864 -52165 -35236
rect -52485 -35890 -52165 -35864
rect -51485 -35236 -51165 -35210
rect -51485 -35864 -51479 -35236
rect -51171 -35864 -51165 -35236
rect -51485 -35890 -51165 -35864
rect -50485 -35236 -50165 -35210
rect -50485 -35864 -50479 -35236
rect -50171 -35864 -50165 -35236
rect -50485 -35890 -50165 -35864
rect -49485 -35236 -49165 -35210
rect -49485 -35864 -49479 -35236
rect -49171 -35864 -49165 -35236
rect -49485 -35890 -49165 -35864
rect -74825 -35896 -48825 -35890
rect -74825 -36204 -74819 -35896
rect -74511 -35928 -74139 -35896
rect -74511 -36172 -74447 -35928
rect -74203 -36172 -74139 -35928
rect -74511 -36204 -74139 -36172
rect -73511 -35928 -73139 -35896
rect -73511 -36172 -73447 -35928
rect -73203 -36172 -73139 -35928
rect -73511 -36204 -73139 -36172
rect -72511 -35928 -72139 -35896
rect -72511 -36172 -72447 -35928
rect -72203 -36172 -72139 -35928
rect -72511 -36204 -72139 -36172
rect -71511 -35928 -71139 -35896
rect -71511 -36172 -71447 -35928
rect -71203 -36172 -71139 -35928
rect -71511 -36204 -71139 -36172
rect -70511 -35928 -70139 -35896
rect -70511 -36172 -70447 -35928
rect -70203 -36172 -70139 -35928
rect -70511 -36204 -70139 -36172
rect -69511 -35928 -69139 -35896
rect -69511 -36172 -69447 -35928
rect -69203 -36172 -69139 -35928
rect -69511 -36204 -69139 -36172
rect -68511 -35928 -68139 -35896
rect -68511 -36172 -68447 -35928
rect -68203 -36172 -68139 -35928
rect -68511 -36204 -68139 -36172
rect -67511 -35928 -67139 -35896
rect -67511 -36172 -67447 -35928
rect -67203 -36172 -67139 -35928
rect -67511 -36204 -67139 -36172
rect -66511 -35928 -66139 -35896
rect -66511 -36172 -66447 -35928
rect -66203 -36172 -66139 -35928
rect -66511 -36204 -66139 -36172
rect -65511 -35928 -65139 -35896
rect -65511 -36172 -65447 -35928
rect -65203 -36172 -65139 -35928
rect -65511 -36204 -65139 -36172
rect -64511 -35928 -64139 -35896
rect -64511 -36172 -64447 -35928
rect -64203 -36172 -64139 -35928
rect -64511 -36204 -64139 -36172
rect -63511 -35928 -63139 -35896
rect -63511 -36172 -63447 -35928
rect -63203 -36172 -63139 -35928
rect -63511 -36204 -63139 -36172
rect -62511 -35928 -62139 -35896
rect -62511 -36172 -62447 -35928
rect -62203 -36172 -62139 -35928
rect -62511 -36204 -62139 -36172
rect -61511 -35928 -61139 -35896
rect -61511 -36172 -61447 -35928
rect -61203 -36172 -61139 -35928
rect -61511 -36204 -61139 -36172
rect -60511 -35928 -60139 -35896
rect -60511 -36172 -60447 -35928
rect -60203 -36172 -60139 -35928
rect -60511 -36204 -60139 -36172
rect -59511 -35928 -59139 -35896
rect -59511 -36172 -59447 -35928
rect -59203 -36172 -59139 -35928
rect -59511 -36204 -59139 -36172
rect -58511 -35928 -58139 -35896
rect -58511 -36172 -58447 -35928
rect -58203 -36172 -58139 -35928
rect -58511 -36204 -58139 -36172
rect -57511 -35928 -57139 -35896
rect -57511 -36172 -57447 -35928
rect -57203 -36172 -57139 -35928
rect -57511 -36204 -57139 -36172
rect -56511 -35928 -56139 -35896
rect -56511 -36172 -56447 -35928
rect -56203 -36172 -56139 -35928
rect -56511 -36204 -56139 -36172
rect -55511 -35928 -55139 -35896
rect -55511 -36172 -55447 -35928
rect -55203 -36172 -55139 -35928
rect -55511 -36204 -55139 -36172
rect -54511 -35928 -54139 -35896
rect -54511 -36172 -54447 -35928
rect -54203 -36172 -54139 -35928
rect -54511 -36204 -54139 -36172
rect -53511 -35928 -53139 -35896
rect -53511 -36172 -53447 -35928
rect -53203 -36172 -53139 -35928
rect -53511 -36204 -53139 -36172
rect -52511 -35928 -52139 -35896
rect -52511 -36172 -52447 -35928
rect -52203 -36172 -52139 -35928
rect -52511 -36204 -52139 -36172
rect -51511 -35928 -51139 -35896
rect -51511 -36172 -51447 -35928
rect -51203 -36172 -51139 -35928
rect -51511 -36204 -51139 -36172
rect -50511 -35928 -50139 -35896
rect -50511 -36172 -50447 -35928
rect -50203 -36172 -50139 -35928
rect -50511 -36204 -50139 -36172
rect -49511 -35928 -49139 -35896
rect -49511 -36172 -49447 -35928
rect -49203 -36172 -49139 -35928
rect -49511 -36204 -49139 -36172
rect -48831 -36204 -48825 -35896
rect -74825 -36210 -48825 -36204
rect -74485 -36236 -74165 -36210
rect -74485 -36864 -74479 -36236
rect -74171 -36864 -74165 -36236
rect -74485 -36890 -74165 -36864
rect -73485 -36236 -73165 -36210
rect -73485 -36864 -73479 -36236
rect -73171 -36864 -73165 -36236
rect -73485 -36890 -73165 -36864
rect -72485 -36236 -72165 -36210
rect -72485 -36864 -72479 -36236
rect -72171 -36864 -72165 -36236
rect -72485 -36890 -72165 -36864
rect -71485 -36236 -71165 -36210
rect -71485 -36864 -71479 -36236
rect -71171 -36864 -71165 -36236
rect -71485 -36890 -71165 -36864
rect -70485 -36236 -70165 -36210
rect -70485 -36864 -70479 -36236
rect -70171 -36864 -70165 -36236
rect -70485 -36890 -70165 -36864
rect -69485 -36236 -69165 -36210
rect -69485 -36864 -69479 -36236
rect -69171 -36864 -69165 -36236
rect -69485 -36890 -69165 -36864
rect -68485 -36236 -68165 -36210
rect -68485 -36864 -68479 -36236
rect -68171 -36864 -68165 -36236
rect -68485 -36890 -68165 -36864
rect -67485 -36236 -67165 -36210
rect -67485 -36864 -67479 -36236
rect -67171 -36864 -67165 -36236
rect -67485 -36890 -67165 -36864
rect -66485 -36236 -66165 -36210
rect -66485 -36864 -66479 -36236
rect -66171 -36864 -66165 -36236
rect -66485 -36890 -66165 -36864
rect -65485 -36236 -65165 -36210
rect -65485 -36864 -65479 -36236
rect -65171 -36864 -65165 -36236
rect -65485 -36890 -65165 -36864
rect -64485 -36236 -64165 -36210
rect -64485 -36864 -64479 -36236
rect -64171 -36864 -64165 -36236
rect -64485 -36890 -64165 -36864
rect -63485 -36236 -63165 -36210
rect -63485 -36864 -63479 -36236
rect -63171 -36864 -63165 -36236
rect -63485 -36890 -63165 -36864
rect -62485 -36236 -62165 -36210
rect -62485 -36864 -62479 -36236
rect -62171 -36864 -62165 -36236
rect -62485 -36890 -62165 -36864
rect -61485 -36236 -61165 -36210
rect -61485 -36864 -61479 -36236
rect -61171 -36864 -61165 -36236
rect -61485 -36890 -61165 -36864
rect -60485 -36236 -60165 -36210
rect -60485 -36864 -60479 -36236
rect -60171 -36864 -60165 -36236
rect -60485 -36890 -60165 -36864
rect -59485 -36236 -59165 -36210
rect -59485 -36864 -59479 -36236
rect -59171 -36864 -59165 -36236
rect -59485 -36890 -59165 -36864
rect -58485 -36236 -58165 -36210
rect -58485 -36864 -58479 -36236
rect -58171 -36864 -58165 -36236
rect -58485 -36890 -58165 -36864
rect -57485 -36236 -57165 -36210
rect -57485 -36864 -57479 -36236
rect -57171 -36864 -57165 -36236
rect -57485 -36890 -57165 -36864
rect -56485 -36236 -56165 -36210
rect -56485 -36864 -56479 -36236
rect -56171 -36864 -56165 -36236
rect -56485 -36890 -56165 -36864
rect -55485 -36236 -55165 -36210
rect -55485 -36864 -55479 -36236
rect -55171 -36864 -55165 -36236
rect -55485 -36890 -55165 -36864
rect -54485 -36236 -54165 -36210
rect -54485 -36864 -54479 -36236
rect -54171 -36864 -54165 -36236
rect -54485 -36890 -54165 -36864
rect -53485 -36236 -53165 -36210
rect -53485 -36864 -53479 -36236
rect -53171 -36864 -53165 -36236
rect -53485 -36890 -53165 -36864
rect -52485 -36236 -52165 -36210
rect -52485 -36864 -52479 -36236
rect -52171 -36864 -52165 -36236
rect -52485 -36890 -52165 -36864
rect -51485 -36236 -51165 -36210
rect -51485 -36864 -51479 -36236
rect -51171 -36864 -51165 -36236
rect -51485 -36890 -51165 -36864
rect -50485 -36236 -50165 -36210
rect -50485 -36864 -50479 -36236
rect -50171 -36864 -50165 -36236
rect -50485 -36890 -50165 -36864
rect -49485 -36236 -49165 -36210
rect -49485 -36864 -49479 -36236
rect -49171 -36864 -49165 -36236
rect -49485 -36890 -49165 -36864
rect -74825 -36896 -48825 -36890
rect -74825 -37204 -74819 -36896
rect -74511 -36928 -74139 -36896
rect -74511 -37172 -74447 -36928
rect -74203 -37172 -74139 -36928
rect -74511 -37204 -74139 -37172
rect -73511 -36928 -73139 -36896
rect -73511 -37172 -73447 -36928
rect -73203 -37172 -73139 -36928
rect -73511 -37204 -73139 -37172
rect -72511 -36928 -72139 -36896
rect -72511 -37172 -72447 -36928
rect -72203 -37172 -72139 -36928
rect -72511 -37204 -72139 -37172
rect -71511 -36928 -71139 -36896
rect -71511 -37172 -71447 -36928
rect -71203 -37172 -71139 -36928
rect -71511 -37204 -71139 -37172
rect -70511 -36928 -70139 -36896
rect -70511 -37172 -70447 -36928
rect -70203 -37172 -70139 -36928
rect -70511 -37204 -70139 -37172
rect -69511 -36928 -69139 -36896
rect -69511 -37172 -69447 -36928
rect -69203 -37172 -69139 -36928
rect -69511 -37204 -69139 -37172
rect -68511 -36928 -68139 -36896
rect -68511 -37172 -68447 -36928
rect -68203 -37172 -68139 -36928
rect -68511 -37204 -68139 -37172
rect -67511 -36928 -67139 -36896
rect -67511 -37172 -67447 -36928
rect -67203 -37172 -67139 -36928
rect -67511 -37204 -67139 -37172
rect -66511 -36928 -66139 -36896
rect -66511 -37172 -66447 -36928
rect -66203 -37172 -66139 -36928
rect -66511 -37204 -66139 -37172
rect -65511 -36928 -65139 -36896
rect -65511 -37172 -65447 -36928
rect -65203 -37172 -65139 -36928
rect -65511 -37204 -65139 -37172
rect -64511 -36928 -64139 -36896
rect -64511 -37172 -64447 -36928
rect -64203 -37172 -64139 -36928
rect -64511 -37204 -64139 -37172
rect -63511 -36928 -63139 -36896
rect -63511 -37172 -63447 -36928
rect -63203 -37172 -63139 -36928
rect -63511 -37204 -63139 -37172
rect -62511 -36928 -62139 -36896
rect -62511 -37172 -62447 -36928
rect -62203 -37172 -62139 -36928
rect -62511 -37204 -62139 -37172
rect -61511 -36928 -61139 -36896
rect -61511 -37172 -61447 -36928
rect -61203 -37172 -61139 -36928
rect -61511 -37204 -61139 -37172
rect -60511 -36928 -60139 -36896
rect -60511 -37172 -60447 -36928
rect -60203 -37172 -60139 -36928
rect -60511 -37204 -60139 -37172
rect -59511 -36928 -59139 -36896
rect -59511 -37172 -59447 -36928
rect -59203 -37172 -59139 -36928
rect -59511 -37204 -59139 -37172
rect -58511 -36928 -58139 -36896
rect -58511 -37172 -58447 -36928
rect -58203 -37172 -58139 -36928
rect -58511 -37204 -58139 -37172
rect -57511 -36928 -57139 -36896
rect -57511 -37172 -57447 -36928
rect -57203 -37172 -57139 -36928
rect -57511 -37204 -57139 -37172
rect -56511 -36928 -56139 -36896
rect -56511 -37172 -56447 -36928
rect -56203 -37172 -56139 -36928
rect -56511 -37204 -56139 -37172
rect -55511 -36928 -55139 -36896
rect -55511 -37172 -55447 -36928
rect -55203 -37172 -55139 -36928
rect -55511 -37204 -55139 -37172
rect -54511 -36928 -54139 -36896
rect -54511 -37172 -54447 -36928
rect -54203 -37172 -54139 -36928
rect -54511 -37204 -54139 -37172
rect -53511 -36928 -53139 -36896
rect -53511 -37172 -53447 -36928
rect -53203 -37172 -53139 -36928
rect -53511 -37204 -53139 -37172
rect -52511 -36928 -52139 -36896
rect -52511 -37172 -52447 -36928
rect -52203 -37172 -52139 -36928
rect -52511 -37204 -52139 -37172
rect -51511 -36928 -51139 -36896
rect -51511 -37172 -51447 -36928
rect -51203 -37172 -51139 -36928
rect -51511 -37204 -51139 -37172
rect -50511 -36928 -50139 -36896
rect -50511 -37172 -50447 -36928
rect -50203 -37172 -50139 -36928
rect -50511 -37204 -50139 -37172
rect -49511 -36928 -49139 -36896
rect -49511 -37172 -49447 -36928
rect -49203 -37172 -49139 -36928
rect -49511 -37204 -49139 -37172
rect -48831 -37204 -48825 -36896
rect -74825 -37210 -48825 -37204
rect -74485 -37236 -74165 -37210
rect -74485 -37864 -74479 -37236
rect -74171 -37864 -74165 -37236
rect -74485 -37890 -74165 -37864
rect -73485 -37236 -73165 -37210
rect -73485 -37864 -73479 -37236
rect -73171 -37864 -73165 -37236
rect -73485 -37890 -73165 -37864
rect -72485 -37236 -72165 -37210
rect -72485 -37864 -72479 -37236
rect -72171 -37864 -72165 -37236
rect -72485 -37890 -72165 -37864
rect -71485 -37236 -71165 -37210
rect -71485 -37864 -71479 -37236
rect -71171 -37864 -71165 -37236
rect -71485 -37890 -71165 -37864
rect -70485 -37236 -70165 -37210
rect -70485 -37864 -70479 -37236
rect -70171 -37864 -70165 -37236
rect -70485 -37890 -70165 -37864
rect -69485 -37236 -69165 -37210
rect -69485 -37864 -69479 -37236
rect -69171 -37864 -69165 -37236
rect -69485 -37890 -69165 -37864
rect -68485 -37236 -68165 -37210
rect -68485 -37864 -68479 -37236
rect -68171 -37864 -68165 -37236
rect -68485 -37890 -68165 -37864
rect -67485 -37236 -67165 -37210
rect -67485 -37864 -67479 -37236
rect -67171 -37864 -67165 -37236
rect -67485 -37890 -67165 -37864
rect -66485 -37236 -66165 -37210
rect -66485 -37864 -66479 -37236
rect -66171 -37864 -66165 -37236
rect -66485 -37890 -66165 -37864
rect -65485 -37236 -65165 -37210
rect -65485 -37864 -65479 -37236
rect -65171 -37864 -65165 -37236
rect -65485 -37890 -65165 -37864
rect -64485 -37236 -64165 -37210
rect -64485 -37864 -64479 -37236
rect -64171 -37864 -64165 -37236
rect -64485 -37890 -64165 -37864
rect -63485 -37236 -63165 -37210
rect -63485 -37864 -63479 -37236
rect -63171 -37864 -63165 -37236
rect -63485 -37890 -63165 -37864
rect -62485 -37236 -62165 -37210
rect -62485 -37864 -62479 -37236
rect -62171 -37864 -62165 -37236
rect -62485 -37890 -62165 -37864
rect -61485 -37236 -61165 -37210
rect -61485 -37864 -61479 -37236
rect -61171 -37864 -61165 -37236
rect -61485 -37890 -61165 -37864
rect -60485 -37236 -60165 -37210
rect -60485 -37864 -60479 -37236
rect -60171 -37864 -60165 -37236
rect -60485 -37890 -60165 -37864
rect -59485 -37236 -59165 -37210
rect -59485 -37864 -59479 -37236
rect -59171 -37864 -59165 -37236
rect -59485 -37890 -59165 -37864
rect -58485 -37236 -58165 -37210
rect -58485 -37864 -58479 -37236
rect -58171 -37864 -58165 -37236
rect -58485 -37890 -58165 -37864
rect -57485 -37236 -57165 -37210
rect -57485 -37864 -57479 -37236
rect -57171 -37864 -57165 -37236
rect -57485 -37890 -57165 -37864
rect -56485 -37236 -56165 -37210
rect -56485 -37864 -56479 -37236
rect -56171 -37864 -56165 -37236
rect -56485 -37890 -56165 -37864
rect -55485 -37236 -55165 -37210
rect -55485 -37864 -55479 -37236
rect -55171 -37864 -55165 -37236
rect -55485 -37890 -55165 -37864
rect -54485 -37236 -54165 -37210
rect -54485 -37864 -54479 -37236
rect -54171 -37864 -54165 -37236
rect -54485 -37890 -54165 -37864
rect -53485 -37236 -53165 -37210
rect -53485 -37864 -53479 -37236
rect -53171 -37864 -53165 -37236
rect -53485 -37890 -53165 -37864
rect -52485 -37236 -52165 -37210
rect -52485 -37864 -52479 -37236
rect -52171 -37864 -52165 -37236
rect -52485 -37890 -52165 -37864
rect -51485 -37236 -51165 -37210
rect -51485 -37864 -51479 -37236
rect -51171 -37864 -51165 -37236
rect -51485 -37890 -51165 -37864
rect -50485 -37236 -50165 -37210
rect -50485 -37864 -50479 -37236
rect -50171 -37864 -50165 -37236
rect -50485 -37890 -50165 -37864
rect -49485 -37236 -49165 -37210
rect -49485 -37864 -49479 -37236
rect -49171 -37864 -49165 -37236
rect -49485 -37890 -49165 -37864
rect -74825 -37896 -48825 -37890
rect -74825 -38204 -74819 -37896
rect -74511 -37928 -74139 -37896
rect -74511 -38172 -74447 -37928
rect -74203 -38172 -74139 -37928
rect -74511 -38204 -74139 -38172
rect -73511 -37928 -73139 -37896
rect -73511 -38172 -73447 -37928
rect -73203 -38172 -73139 -37928
rect -73511 -38204 -73139 -38172
rect -72511 -37928 -72139 -37896
rect -72511 -38172 -72447 -37928
rect -72203 -38172 -72139 -37928
rect -72511 -38204 -72139 -38172
rect -71511 -37928 -71139 -37896
rect -71511 -38172 -71447 -37928
rect -71203 -38172 -71139 -37928
rect -71511 -38204 -71139 -38172
rect -70511 -37928 -70139 -37896
rect -70511 -38172 -70447 -37928
rect -70203 -38172 -70139 -37928
rect -70511 -38204 -70139 -38172
rect -69511 -37928 -69139 -37896
rect -69511 -38172 -69447 -37928
rect -69203 -38172 -69139 -37928
rect -69511 -38204 -69139 -38172
rect -68511 -37928 -68139 -37896
rect -68511 -38172 -68447 -37928
rect -68203 -38172 -68139 -37928
rect -68511 -38204 -68139 -38172
rect -67511 -37928 -67139 -37896
rect -67511 -38172 -67447 -37928
rect -67203 -38172 -67139 -37928
rect -67511 -38204 -67139 -38172
rect -66511 -37928 -66139 -37896
rect -66511 -38172 -66447 -37928
rect -66203 -38172 -66139 -37928
rect -66511 -38204 -66139 -38172
rect -65511 -37928 -65139 -37896
rect -65511 -38172 -65447 -37928
rect -65203 -38172 -65139 -37928
rect -65511 -38204 -65139 -38172
rect -64511 -37928 -64139 -37896
rect -64511 -38172 -64447 -37928
rect -64203 -38172 -64139 -37928
rect -64511 -38204 -64139 -38172
rect -63511 -37928 -63139 -37896
rect -63511 -38172 -63447 -37928
rect -63203 -38172 -63139 -37928
rect -63511 -38204 -63139 -38172
rect -62511 -37928 -62139 -37896
rect -62511 -38172 -62447 -37928
rect -62203 -38172 -62139 -37928
rect -62511 -38204 -62139 -38172
rect -61511 -37928 -61139 -37896
rect -61511 -38172 -61447 -37928
rect -61203 -38172 -61139 -37928
rect -61511 -38204 -61139 -38172
rect -60511 -37928 -60139 -37896
rect -60511 -38172 -60447 -37928
rect -60203 -38172 -60139 -37928
rect -60511 -38204 -60139 -38172
rect -59511 -37928 -59139 -37896
rect -59511 -38172 -59447 -37928
rect -59203 -38172 -59139 -37928
rect -59511 -38204 -59139 -38172
rect -58511 -37928 -58139 -37896
rect -58511 -38172 -58447 -37928
rect -58203 -38172 -58139 -37928
rect -58511 -38204 -58139 -38172
rect -57511 -37928 -57139 -37896
rect -57511 -38172 -57447 -37928
rect -57203 -38172 -57139 -37928
rect -57511 -38204 -57139 -38172
rect -56511 -37928 -56139 -37896
rect -56511 -38172 -56447 -37928
rect -56203 -38172 -56139 -37928
rect -56511 -38204 -56139 -38172
rect -55511 -37928 -55139 -37896
rect -55511 -38172 -55447 -37928
rect -55203 -38172 -55139 -37928
rect -55511 -38204 -55139 -38172
rect -54511 -37928 -54139 -37896
rect -54511 -38172 -54447 -37928
rect -54203 -38172 -54139 -37928
rect -54511 -38204 -54139 -38172
rect -53511 -37928 -53139 -37896
rect -53511 -38172 -53447 -37928
rect -53203 -38172 -53139 -37928
rect -53511 -38204 -53139 -38172
rect -52511 -37928 -52139 -37896
rect -52511 -38172 -52447 -37928
rect -52203 -38172 -52139 -37928
rect -52511 -38204 -52139 -38172
rect -51511 -37928 -51139 -37896
rect -51511 -38172 -51447 -37928
rect -51203 -38172 -51139 -37928
rect -51511 -38204 -51139 -38172
rect -50511 -37928 -50139 -37896
rect -50511 -38172 -50447 -37928
rect -50203 -38172 -50139 -37928
rect -50511 -38204 -50139 -38172
rect -49511 -37928 -49139 -37896
rect -49511 -38172 -49447 -37928
rect -49203 -38172 -49139 -37928
rect -49511 -38204 -49139 -38172
rect -48831 -38204 -48825 -37896
rect -74825 -38210 -48825 -38204
rect -74485 -38236 -74165 -38210
rect -74485 -38864 -74479 -38236
rect -74171 -38864 -74165 -38236
rect -74485 -38890 -74165 -38864
rect -73485 -38236 -73165 -38210
rect -73485 -38864 -73479 -38236
rect -73171 -38864 -73165 -38236
rect -73485 -38890 -73165 -38864
rect -72485 -38236 -72165 -38210
rect -72485 -38864 -72479 -38236
rect -72171 -38864 -72165 -38236
rect -72485 -38890 -72165 -38864
rect -71485 -38236 -71165 -38210
rect -71485 -38864 -71479 -38236
rect -71171 -38864 -71165 -38236
rect -71485 -38890 -71165 -38864
rect -70485 -38236 -70165 -38210
rect -70485 -38864 -70479 -38236
rect -70171 -38864 -70165 -38236
rect -70485 -38890 -70165 -38864
rect -69485 -38236 -69165 -38210
rect -69485 -38864 -69479 -38236
rect -69171 -38864 -69165 -38236
rect -69485 -38890 -69165 -38864
rect -68485 -38236 -68165 -38210
rect -68485 -38864 -68479 -38236
rect -68171 -38864 -68165 -38236
rect -68485 -38890 -68165 -38864
rect -67485 -38236 -67165 -38210
rect -67485 -38864 -67479 -38236
rect -67171 -38864 -67165 -38236
rect -67485 -38890 -67165 -38864
rect -66485 -38236 -66165 -38210
rect -66485 -38864 -66479 -38236
rect -66171 -38864 -66165 -38236
rect -66485 -38890 -66165 -38864
rect -65485 -38236 -65165 -38210
rect -65485 -38864 -65479 -38236
rect -65171 -38864 -65165 -38236
rect -65485 -38890 -65165 -38864
rect -64485 -38236 -64165 -38210
rect -64485 -38864 -64479 -38236
rect -64171 -38864 -64165 -38236
rect -64485 -38890 -64165 -38864
rect -63485 -38236 -63165 -38210
rect -63485 -38864 -63479 -38236
rect -63171 -38864 -63165 -38236
rect -63485 -38890 -63165 -38864
rect -62485 -38236 -62165 -38210
rect -62485 -38864 -62479 -38236
rect -62171 -38864 -62165 -38236
rect -62485 -38890 -62165 -38864
rect -61485 -38236 -61165 -38210
rect -61485 -38864 -61479 -38236
rect -61171 -38864 -61165 -38236
rect -61485 -38890 -61165 -38864
rect -60485 -38236 -60165 -38210
rect -60485 -38864 -60479 -38236
rect -60171 -38864 -60165 -38236
rect -60485 -38890 -60165 -38864
rect -59485 -38236 -59165 -38210
rect -59485 -38864 -59479 -38236
rect -59171 -38864 -59165 -38236
rect -59485 -38890 -59165 -38864
rect -58485 -38236 -58165 -38210
rect -58485 -38864 -58479 -38236
rect -58171 -38864 -58165 -38236
rect -58485 -38890 -58165 -38864
rect -57485 -38236 -57165 -38210
rect -57485 -38864 -57479 -38236
rect -57171 -38864 -57165 -38236
rect -57485 -38890 -57165 -38864
rect -56485 -38236 -56165 -38210
rect -56485 -38864 -56479 -38236
rect -56171 -38864 -56165 -38236
rect -56485 -38890 -56165 -38864
rect -55485 -38236 -55165 -38210
rect -55485 -38864 -55479 -38236
rect -55171 -38864 -55165 -38236
rect -55485 -38890 -55165 -38864
rect -54485 -38236 -54165 -38210
rect -54485 -38864 -54479 -38236
rect -54171 -38864 -54165 -38236
rect -54485 -38890 -54165 -38864
rect -53485 -38236 -53165 -38210
rect -53485 -38864 -53479 -38236
rect -53171 -38864 -53165 -38236
rect -53485 -38890 -53165 -38864
rect -52485 -38236 -52165 -38210
rect -52485 -38864 -52479 -38236
rect -52171 -38864 -52165 -38236
rect -52485 -38890 -52165 -38864
rect -51485 -38236 -51165 -38210
rect -51485 -38864 -51479 -38236
rect -51171 -38864 -51165 -38236
rect -51485 -38890 -51165 -38864
rect -50485 -38236 -50165 -38210
rect -50485 -38864 -50479 -38236
rect -50171 -38864 -50165 -38236
rect -50485 -38890 -50165 -38864
rect -49485 -38236 -49165 -38210
rect -49485 -38864 -49479 -38236
rect -49171 -38864 -49165 -38236
rect -49485 -38890 -49165 -38864
rect -74825 -38896 -48825 -38890
rect -74825 -39204 -74819 -38896
rect -74511 -38928 -74139 -38896
rect -74511 -39172 -74447 -38928
rect -74203 -39172 -74139 -38928
rect -74511 -39204 -74139 -39172
rect -73511 -38928 -73139 -38896
rect -73511 -39172 -73447 -38928
rect -73203 -39172 -73139 -38928
rect -73511 -39204 -73139 -39172
rect -72511 -38928 -72139 -38896
rect -72511 -39172 -72447 -38928
rect -72203 -39172 -72139 -38928
rect -72511 -39204 -72139 -39172
rect -71511 -38928 -71139 -38896
rect -71511 -39172 -71447 -38928
rect -71203 -39172 -71139 -38928
rect -71511 -39204 -71139 -39172
rect -70511 -38928 -70139 -38896
rect -70511 -39172 -70447 -38928
rect -70203 -39172 -70139 -38928
rect -70511 -39204 -70139 -39172
rect -69511 -38928 -69139 -38896
rect -69511 -39172 -69447 -38928
rect -69203 -39172 -69139 -38928
rect -69511 -39204 -69139 -39172
rect -68511 -38928 -68139 -38896
rect -68511 -39172 -68447 -38928
rect -68203 -39172 -68139 -38928
rect -68511 -39204 -68139 -39172
rect -67511 -38928 -67139 -38896
rect -67511 -39172 -67447 -38928
rect -67203 -39172 -67139 -38928
rect -67511 -39204 -67139 -39172
rect -66511 -38928 -66139 -38896
rect -66511 -39172 -66447 -38928
rect -66203 -39172 -66139 -38928
rect -66511 -39204 -66139 -39172
rect -65511 -38928 -65139 -38896
rect -65511 -39172 -65447 -38928
rect -65203 -39172 -65139 -38928
rect -65511 -39204 -65139 -39172
rect -64511 -38928 -64139 -38896
rect -64511 -39172 -64447 -38928
rect -64203 -39172 -64139 -38928
rect -64511 -39204 -64139 -39172
rect -63511 -38928 -63139 -38896
rect -63511 -39172 -63447 -38928
rect -63203 -39172 -63139 -38928
rect -63511 -39204 -63139 -39172
rect -62511 -38928 -62139 -38896
rect -62511 -39172 -62447 -38928
rect -62203 -39172 -62139 -38928
rect -62511 -39204 -62139 -39172
rect -61511 -38928 -61139 -38896
rect -61511 -39172 -61447 -38928
rect -61203 -39172 -61139 -38928
rect -61511 -39204 -61139 -39172
rect -60511 -38928 -60139 -38896
rect -60511 -39172 -60447 -38928
rect -60203 -39172 -60139 -38928
rect -60511 -39204 -60139 -39172
rect -59511 -38928 -59139 -38896
rect -59511 -39172 -59447 -38928
rect -59203 -39172 -59139 -38928
rect -59511 -39204 -59139 -39172
rect -58511 -38928 -58139 -38896
rect -58511 -39172 -58447 -38928
rect -58203 -39172 -58139 -38928
rect -58511 -39204 -58139 -39172
rect -57511 -38928 -57139 -38896
rect -57511 -39172 -57447 -38928
rect -57203 -39172 -57139 -38928
rect -57511 -39204 -57139 -39172
rect -56511 -38928 -56139 -38896
rect -56511 -39172 -56447 -38928
rect -56203 -39172 -56139 -38928
rect -56511 -39204 -56139 -39172
rect -55511 -38928 -55139 -38896
rect -55511 -39172 -55447 -38928
rect -55203 -39172 -55139 -38928
rect -55511 -39204 -55139 -39172
rect -54511 -38928 -54139 -38896
rect -54511 -39172 -54447 -38928
rect -54203 -39172 -54139 -38928
rect -54511 -39204 -54139 -39172
rect -53511 -38928 -53139 -38896
rect -53511 -39172 -53447 -38928
rect -53203 -39172 -53139 -38928
rect -53511 -39204 -53139 -39172
rect -52511 -38928 -52139 -38896
rect -52511 -39172 -52447 -38928
rect -52203 -39172 -52139 -38928
rect -52511 -39204 -52139 -39172
rect -51511 -38928 -51139 -38896
rect -51511 -39172 -51447 -38928
rect -51203 -39172 -51139 -38928
rect -51511 -39204 -51139 -39172
rect -50511 -38928 -50139 -38896
rect -50511 -39172 -50447 -38928
rect -50203 -39172 -50139 -38928
rect -50511 -39204 -50139 -39172
rect -49511 -38928 -49139 -38896
rect -49511 -39172 -49447 -38928
rect -49203 -39172 -49139 -38928
rect -49511 -39204 -49139 -39172
rect -48831 -39204 -48825 -38896
rect -74825 -39210 -48825 -39204
rect -74485 -39236 -74165 -39210
rect -74485 -39864 -74479 -39236
rect -74171 -39864 -74165 -39236
rect -74485 -39890 -74165 -39864
rect -73485 -39236 -73165 -39210
rect -73485 -39864 -73479 -39236
rect -73171 -39864 -73165 -39236
rect -73485 -39890 -73165 -39864
rect -72485 -39236 -72165 -39210
rect -72485 -39864 -72479 -39236
rect -72171 -39864 -72165 -39236
rect -72485 -39890 -72165 -39864
rect -71485 -39236 -71165 -39210
rect -71485 -39864 -71479 -39236
rect -71171 -39864 -71165 -39236
rect -71485 -39890 -71165 -39864
rect -70485 -39236 -70165 -39210
rect -70485 -39864 -70479 -39236
rect -70171 -39864 -70165 -39236
rect -70485 -39890 -70165 -39864
rect -69485 -39236 -69165 -39210
rect -69485 -39864 -69479 -39236
rect -69171 -39864 -69165 -39236
rect -69485 -39890 -69165 -39864
rect -68485 -39236 -68165 -39210
rect -68485 -39864 -68479 -39236
rect -68171 -39864 -68165 -39236
rect -68485 -39890 -68165 -39864
rect -67485 -39236 -67165 -39210
rect -67485 -39864 -67479 -39236
rect -67171 -39864 -67165 -39236
rect -67485 -39890 -67165 -39864
rect -66485 -39236 -66165 -39210
rect -66485 -39864 -66479 -39236
rect -66171 -39864 -66165 -39236
rect -66485 -39890 -66165 -39864
rect -65485 -39236 -65165 -39210
rect -65485 -39864 -65479 -39236
rect -65171 -39864 -65165 -39236
rect -65485 -39890 -65165 -39864
rect -64485 -39236 -64165 -39210
rect -64485 -39864 -64479 -39236
rect -64171 -39864 -64165 -39236
rect -64485 -39890 -64165 -39864
rect -63485 -39236 -63165 -39210
rect -63485 -39864 -63479 -39236
rect -63171 -39864 -63165 -39236
rect -63485 -39890 -63165 -39864
rect -62485 -39236 -62165 -39210
rect -62485 -39864 -62479 -39236
rect -62171 -39864 -62165 -39236
rect -62485 -39890 -62165 -39864
rect -61485 -39236 -61165 -39210
rect -61485 -39864 -61479 -39236
rect -61171 -39864 -61165 -39236
rect -61485 -39890 -61165 -39864
rect -60485 -39236 -60165 -39210
rect -60485 -39864 -60479 -39236
rect -60171 -39864 -60165 -39236
rect -60485 -39890 -60165 -39864
rect -59485 -39236 -59165 -39210
rect -59485 -39864 -59479 -39236
rect -59171 -39864 -59165 -39236
rect -59485 -39890 -59165 -39864
rect -58485 -39236 -58165 -39210
rect -58485 -39864 -58479 -39236
rect -58171 -39864 -58165 -39236
rect -58485 -39890 -58165 -39864
rect -57485 -39236 -57165 -39210
rect -57485 -39864 -57479 -39236
rect -57171 -39864 -57165 -39236
rect -57485 -39890 -57165 -39864
rect -56485 -39236 -56165 -39210
rect -56485 -39864 -56479 -39236
rect -56171 -39864 -56165 -39236
rect -56485 -39890 -56165 -39864
rect -55485 -39236 -55165 -39210
rect -55485 -39864 -55479 -39236
rect -55171 -39864 -55165 -39236
rect -55485 -39890 -55165 -39864
rect -54485 -39236 -54165 -39210
rect -54485 -39864 -54479 -39236
rect -54171 -39864 -54165 -39236
rect -54485 -39890 -54165 -39864
rect -53485 -39236 -53165 -39210
rect -53485 -39864 -53479 -39236
rect -53171 -39864 -53165 -39236
rect -53485 -39890 -53165 -39864
rect -52485 -39236 -52165 -39210
rect -52485 -39864 -52479 -39236
rect -52171 -39864 -52165 -39236
rect -52485 -39890 -52165 -39864
rect -51485 -39236 -51165 -39210
rect -51485 -39864 -51479 -39236
rect -51171 -39864 -51165 -39236
rect -51485 -39890 -51165 -39864
rect -50485 -39236 -50165 -39210
rect -50485 -39864 -50479 -39236
rect -50171 -39864 -50165 -39236
rect -50485 -39890 -50165 -39864
rect -49485 -39236 -49165 -39210
rect -49485 -39864 -49479 -39236
rect -49171 -39864 -49165 -39236
rect -49485 -39890 -49165 -39864
rect -74825 -39896 -48825 -39890
rect -74825 -40204 -74819 -39896
rect -74511 -39928 -74139 -39896
rect -74511 -40172 -74447 -39928
rect -74203 -40172 -74139 -39928
rect -74511 -40204 -74139 -40172
rect -73511 -39928 -73139 -39896
rect -73511 -40172 -73447 -39928
rect -73203 -40172 -73139 -39928
rect -73511 -40204 -73139 -40172
rect -72511 -39928 -72139 -39896
rect -72511 -40172 -72447 -39928
rect -72203 -40172 -72139 -39928
rect -72511 -40204 -72139 -40172
rect -71511 -39928 -71139 -39896
rect -71511 -40172 -71447 -39928
rect -71203 -40172 -71139 -39928
rect -71511 -40204 -71139 -40172
rect -70511 -39928 -70139 -39896
rect -70511 -40172 -70447 -39928
rect -70203 -40172 -70139 -39928
rect -70511 -40204 -70139 -40172
rect -69511 -39928 -69139 -39896
rect -69511 -40172 -69447 -39928
rect -69203 -40172 -69139 -39928
rect -69511 -40204 -69139 -40172
rect -68511 -39928 -68139 -39896
rect -68511 -40172 -68447 -39928
rect -68203 -40172 -68139 -39928
rect -68511 -40204 -68139 -40172
rect -67511 -39928 -67139 -39896
rect -67511 -40172 -67447 -39928
rect -67203 -40172 -67139 -39928
rect -67511 -40204 -67139 -40172
rect -66511 -39928 -66139 -39896
rect -66511 -40172 -66447 -39928
rect -66203 -40172 -66139 -39928
rect -66511 -40204 -66139 -40172
rect -65511 -39928 -65139 -39896
rect -65511 -40172 -65447 -39928
rect -65203 -40172 -65139 -39928
rect -65511 -40204 -65139 -40172
rect -64511 -39928 -64139 -39896
rect -64511 -40172 -64447 -39928
rect -64203 -40172 -64139 -39928
rect -64511 -40204 -64139 -40172
rect -63511 -39928 -63139 -39896
rect -63511 -40172 -63447 -39928
rect -63203 -40172 -63139 -39928
rect -63511 -40204 -63139 -40172
rect -62511 -39928 -62139 -39896
rect -62511 -40172 -62447 -39928
rect -62203 -40172 -62139 -39928
rect -62511 -40204 -62139 -40172
rect -61511 -39928 -61139 -39896
rect -61511 -40172 -61447 -39928
rect -61203 -40172 -61139 -39928
rect -61511 -40204 -61139 -40172
rect -60511 -39928 -60139 -39896
rect -60511 -40172 -60447 -39928
rect -60203 -40172 -60139 -39928
rect -60511 -40204 -60139 -40172
rect -59511 -39928 -59139 -39896
rect -59511 -40172 -59447 -39928
rect -59203 -40172 -59139 -39928
rect -59511 -40204 -59139 -40172
rect -58511 -39928 -58139 -39896
rect -58511 -40172 -58447 -39928
rect -58203 -40172 -58139 -39928
rect -58511 -40204 -58139 -40172
rect -57511 -39928 -57139 -39896
rect -57511 -40172 -57447 -39928
rect -57203 -40172 -57139 -39928
rect -57511 -40204 -57139 -40172
rect -56511 -39928 -56139 -39896
rect -56511 -40172 -56447 -39928
rect -56203 -40172 -56139 -39928
rect -56511 -40204 -56139 -40172
rect -55511 -39928 -55139 -39896
rect -55511 -40172 -55447 -39928
rect -55203 -40172 -55139 -39928
rect -55511 -40204 -55139 -40172
rect -54511 -39928 -54139 -39896
rect -54511 -40172 -54447 -39928
rect -54203 -40172 -54139 -39928
rect -54511 -40204 -54139 -40172
rect -53511 -39928 -53139 -39896
rect -53511 -40172 -53447 -39928
rect -53203 -40172 -53139 -39928
rect -53511 -40204 -53139 -40172
rect -52511 -39928 -52139 -39896
rect -52511 -40172 -52447 -39928
rect -52203 -40172 -52139 -39928
rect -52511 -40204 -52139 -40172
rect -51511 -39928 -51139 -39896
rect -51511 -40172 -51447 -39928
rect -51203 -40172 -51139 -39928
rect -51511 -40204 -51139 -40172
rect -50511 -39928 -50139 -39896
rect -50511 -40172 -50447 -39928
rect -50203 -40172 -50139 -39928
rect -50511 -40204 -50139 -40172
rect -49511 -39928 -49139 -39896
rect -49511 -40172 -49447 -39928
rect -49203 -40172 -49139 -39928
rect -49511 -40204 -49139 -40172
rect -48831 -40204 -48825 -39896
rect -74825 -40210 -48825 -40204
rect -74485 -40236 -74165 -40210
rect -74485 -40864 -74479 -40236
rect -74171 -40864 -74165 -40236
rect -74485 -40890 -74165 -40864
rect -73485 -40236 -73165 -40210
rect -73485 -40864 -73479 -40236
rect -73171 -40864 -73165 -40236
rect -73485 -40890 -73165 -40864
rect -72485 -40236 -72165 -40210
rect -72485 -40864 -72479 -40236
rect -72171 -40864 -72165 -40236
rect -72485 -40890 -72165 -40864
rect -71485 -40236 -71165 -40210
rect -71485 -40864 -71479 -40236
rect -71171 -40864 -71165 -40236
rect -71485 -40890 -71165 -40864
rect -70485 -40236 -70165 -40210
rect -70485 -40864 -70479 -40236
rect -70171 -40864 -70165 -40236
rect -70485 -40890 -70165 -40864
rect -69485 -40236 -69165 -40210
rect -69485 -40864 -69479 -40236
rect -69171 -40864 -69165 -40236
rect -69485 -40890 -69165 -40864
rect -68485 -40236 -68165 -40210
rect -68485 -40864 -68479 -40236
rect -68171 -40864 -68165 -40236
rect -68485 -40890 -68165 -40864
rect -67485 -40236 -67165 -40210
rect -67485 -40864 -67479 -40236
rect -67171 -40864 -67165 -40236
rect -67485 -40890 -67165 -40864
rect -66485 -40236 -66165 -40210
rect -66485 -40864 -66479 -40236
rect -66171 -40864 -66165 -40236
rect -66485 -40890 -66165 -40864
rect -65485 -40236 -65165 -40210
rect -65485 -40864 -65479 -40236
rect -65171 -40864 -65165 -40236
rect -65485 -40890 -65165 -40864
rect -64485 -40236 -64165 -40210
rect -64485 -40864 -64479 -40236
rect -64171 -40864 -64165 -40236
rect -64485 -40890 -64165 -40864
rect -63485 -40236 -63165 -40210
rect -63485 -40864 -63479 -40236
rect -63171 -40864 -63165 -40236
rect -63485 -40890 -63165 -40864
rect -62485 -40236 -62165 -40210
rect -62485 -40864 -62479 -40236
rect -62171 -40864 -62165 -40236
rect -62485 -40890 -62165 -40864
rect -61485 -40236 -61165 -40210
rect -61485 -40864 -61479 -40236
rect -61171 -40864 -61165 -40236
rect -61485 -40890 -61165 -40864
rect -60485 -40236 -60165 -40210
rect -60485 -40864 -60479 -40236
rect -60171 -40864 -60165 -40236
rect -60485 -40890 -60165 -40864
rect -59485 -40236 -59165 -40210
rect -59485 -40864 -59479 -40236
rect -59171 -40864 -59165 -40236
rect -59485 -40890 -59165 -40864
rect -58485 -40236 -58165 -40210
rect -58485 -40864 -58479 -40236
rect -58171 -40864 -58165 -40236
rect -58485 -40890 -58165 -40864
rect -57485 -40236 -57165 -40210
rect -57485 -40864 -57479 -40236
rect -57171 -40864 -57165 -40236
rect -57485 -40890 -57165 -40864
rect -56485 -40236 -56165 -40210
rect -56485 -40864 -56479 -40236
rect -56171 -40864 -56165 -40236
rect -56485 -40890 -56165 -40864
rect -55485 -40236 -55165 -40210
rect -55485 -40864 -55479 -40236
rect -55171 -40864 -55165 -40236
rect -55485 -40890 -55165 -40864
rect -54485 -40236 -54165 -40210
rect -54485 -40864 -54479 -40236
rect -54171 -40864 -54165 -40236
rect -54485 -40890 -54165 -40864
rect -53485 -40236 -53165 -40210
rect -53485 -40864 -53479 -40236
rect -53171 -40864 -53165 -40236
rect -53485 -40890 -53165 -40864
rect -52485 -40236 -52165 -40210
rect -52485 -40864 -52479 -40236
rect -52171 -40864 -52165 -40236
rect -52485 -40890 -52165 -40864
rect -51485 -40236 -51165 -40210
rect -51485 -40864 -51479 -40236
rect -51171 -40864 -51165 -40236
rect -51485 -40890 -51165 -40864
rect -50485 -40236 -50165 -40210
rect -50485 -40864 -50479 -40236
rect -50171 -40864 -50165 -40236
rect -50485 -40890 -50165 -40864
rect -49485 -40236 -49165 -40210
rect -49485 -40864 -49479 -40236
rect -49171 -40864 -49165 -40236
rect -49485 -40890 -49165 -40864
rect -74825 -40896 -48825 -40890
rect -74825 -41204 -74819 -40896
rect -74511 -40928 -74139 -40896
rect -74511 -41172 -74447 -40928
rect -74203 -41172 -74139 -40928
rect -74511 -41204 -74139 -41172
rect -73511 -40928 -73139 -40896
rect -73511 -41172 -73447 -40928
rect -73203 -41172 -73139 -40928
rect -73511 -41204 -73139 -41172
rect -72511 -40928 -72139 -40896
rect -72511 -41172 -72447 -40928
rect -72203 -41172 -72139 -40928
rect -72511 -41204 -72139 -41172
rect -71511 -40928 -71139 -40896
rect -71511 -41172 -71447 -40928
rect -71203 -41172 -71139 -40928
rect -71511 -41204 -71139 -41172
rect -70511 -40928 -70139 -40896
rect -70511 -41172 -70447 -40928
rect -70203 -41172 -70139 -40928
rect -70511 -41204 -70139 -41172
rect -69511 -40928 -69139 -40896
rect -69511 -41172 -69447 -40928
rect -69203 -41172 -69139 -40928
rect -69511 -41204 -69139 -41172
rect -68511 -40928 -68139 -40896
rect -68511 -41172 -68447 -40928
rect -68203 -41172 -68139 -40928
rect -68511 -41204 -68139 -41172
rect -67511 -40928 -67139 -40896
rect -67511 -41172 -67447 -40928
rect -67203 -41172 -67139 -40928
rect -67511 -41204 -67139 -41172
rect -66511 -40928 -66139 -40896
rect -66511 -41172 -66447 -40928
rect -66203 -41172 -66139 -40928
rect -66511 -41204 -66139 -41172
rect -65511 -40928 -65139 -40896
rect -65511 -41172 -65447 -40928
rect -65203 -41172 -65139 -40928
rect -65511 -41204 -65139 -41172
rect -64511 -40928 -64139 -40896
rect -64511 -41172 -64447 -40928
rect -64203 -41172 -64139 -40928
rect -64511 -41204 -64139 -41172
rect -63511 -40928 -63139 -40896
rect -63511 -41172 -63447 -40928
rect -63203 -41172 -63139 -40928
rect -63511 -41204 -63139 -41172
rect -62511 -40928 -62139 -40896
rect -62511 -41172 -62447 -40928
rect -62203 -41172 -62139 -40928
rect -62511 -41204 -62139 -41172
rect -61511 -40928 -61139 -40896
rect -61511 -41172 -61447 -40928
rect -61203 -41172 -61139 -40928
rect -61511 -41204 -61139 -41172
rect -60511 -40928 -60139 -40896
rect -60511 -41172 -60447 -40928
rect -60203 -41172 -60139 -40928
rect -60511 -41204 -60139 -41172
rect -59511 -40928 -59139 -40896
rect -59511 -41172 -59447 -40928
rect -59203 -41172 -59139 -40928
rect -59511 -41204 -59139 -41172
rect -58511 -40928 -58139 -40896
rect -58511 -41172 -58447 -40928
rect -58203 -41172 -58139 -40928
rect -58511 -41204 -58139 -41172
rect -57511 -40928 -57139 -40896
rect -57511 -41172 -57447 -40928
rect -57203 -41172 -57139 -40928
rect -57511 -41204 -57139 -41172
rect -56511 -40928 -56139 -40896
rect -56511 -41172 -56447 -40928
rect -56203 -41172 -56139 -40928
rect -56511 -41204 -56139 -41172
rect -55511 -40928 -55139 -40896
rect -55511 -41172 -55447 -40928
rect -55203 -41172 -55139 -40928
rect -55511 -41204 -55139 -41172
rect -54511 -40928 -54139 -40896
rect -54511 -41172 -54447 -40928
rect -54203 -41172 -54139 -40928
rect -54511 -41204 -54139 -41172
rect -53511 -40928 -53139 -40896
rect -53511 -41172 -53447 -40928
rect -53203 -41172 -53139 -40928
rect -53511 -41204 -53139 -41172
rect -52511 -40928 -52139 -40896
rect -52511 -41172 -52447 -40928
rect -52203 -41172 -52139 -40928
rect -52511 -41204 -52139 -41172
rect -51511 -40928 -51139 -40896
rect -51511 -41172 -51447 -40928
rect -51203 -41172 -51139 -40928
rect -51511 -41204 -51139 -41172
rect -50511 -40928 -50139 -40896
rect -50511 -41172 -50447 -40928
rect -50203 -41172 -50139 -40928
rect -50511 -41204 -50139 -41172
rect -49511 -40928 -49139 -40896
rect -49511 -41172 -49447 -40928
rect -49203 -41172 -49139 -40928
rect -49511 -41204 -49139 -41172
rect -48831 -41204 -48825 -40896
rect -74825 -41210 -48825 -41204
rect -74485 -41236 -74165 -41210
rect -74485 -41864 -74479 -41236
rect -74171 -41864 -74165 -41236
rect -74485 -41890 -74165 -41864
rect -73485 -41236 -73165 -41210
rect -73485 -41864 -73479 -41236
rect -73171 -41864 -73165 -41236
rect -73485 -41890 -73165 -41864
rect -72485 -41236 -72165 -41210
rect -72485 -41864 -72479 -41236
rect -72171 -41864 -72165 -41236
rect -72485 -41890 -72165 -41864
rect -71485 -41236 -71165 -41210
rect -71485 -41864 -71479 -41236
rect -71171 -41864 -71165 -41236
rect -71485 -41890 -71165 -41864
rect -70485 -41236 -70165 -41210
rect -70485 -41864 -70479 -41236
rect -70171 -41864 -70165 -41236
rect -70485 -41890 -70165 -41864
rect -69485 -41236 -69165 -41210
rect -69485 -41864 -69479 -41236
rect -69171 -41864 -69165 -41236
rect -69485 -41890 -69165 -41864
rect -68485 -41236 -68165 -41210
rect -68485 -41864 -68479 -41236
rect -68171 -41864 -68165 -41236
rect -68485 -41890 -68165 -41864
rect -67485 -41236 -67165 -41210
rect -67485 -41864 -67479 -41236
rect -67171 -41864 -67165 -41236
rect -67485 -41890 -67165 -41864
rect -66485 -41236 -66165 -41210
rect -66485 -41864 -66479 -41236
rect -66171 -41864 -66165 -41236
rect -66485 -41890 -66165 -41864
rect -65485 -41236 -65165 -41210
rect -65485 -41864 -65479 -41236
rect -65171 -41864 -65165 -41236
rect -65485 -41890 -65165 -41864
rect -64485 -41236 -64165 -41210
rect -64485 -41864 -64479 -41236
rect -64171 -41864 -64165 -41236
rect -64485 -41890 -64165 -41864
rect -63485 -41236 -63165 -41210
rect -63485 -41864 -63479 -41236
rect -63171 -41864 -63165 -41236
rect -63485 -41890 -63165 -41864
rect -62485 -41236 -62165 -41210
rect -62485 -41864 -62479 -41236
rect -62171 -41864 -62165 -41236
rect -62485 -41890 -62165 -41864
rect -61485 -41236 -61165 -41210
rect -61485 -41864 -61479 -41236
rect -61171 -41864 -61165 -41236
rect -61485 -41890 -61165 -41864
rect -60485 -41236 -60165 -41210
rect -60485 -41864 -60479 -41236
rect -60171 -41864 -60165 -41236
rect -60485 -41890 -60165 -41864
rect -59485 -41236 -59165 -41210
rect -59485 -41864 -59479 -41236
rect -59171 -41864 -59165 -41236
rect -59485 -41890 -59165 -41864
rect -58485 -41236 -58165 -41210
rect -58485 -41864 -58479 -41236
rect -58171 -41864 -58165 -41236
rect -58485 -41890 -58165 -41864
rect -57485 -41236 -57165 -41210
rect -57485 -41864 -57479 -41236
rect -57171 -41864 -57165 -41236
rect -57485 -41890 -57165 -41864
rect -56485 -41236 -56165 -41210
rect -56485 -41864 -56479 -41236
rect -56171 -41864 -56165 -41236
rect -56485 -41890 -56165 -41864
rect -55485 -41236 -55165 -41210
rect -55485 -41864 -55479 -41236
rect -55171 -41864 -55165 -41236
rect -55485 -41890 -55165 -41864
rect -54485 -41236 -54165 -41210
rect -54485 -41864 -54479 -41236
rect -54171 -41864 -54165 -41236
rect -54485 -41890 -54165 -41864
rect -53485 -41236 -53165 -41210
rect -53485 -41864 -53479 -41236
rect -53171 -41864 -53165 -41236
rect -53485 -41890 -53165 -41864
rect -52485 -41236 -52165 -41210
rect -52485 -41864 -52479 -41236
rect -52171 -41864 -52165 -41236
rect -52485 -41890 -52165 -41864
rect -51485 -41236 -51165 -41210
rect -51485 -41864 -51479 -41236
rect -51171 -41864 -51165 -41236
rect -51485 -41890 -51165 -41864
rect -50485 -41236 -50165 -41210
rect -50485 -41864 -50479 -41236
rect -50171 -41864 -50165 -41236
rect -50485 -41890 -50165 -41864
rect -49485 -41236 -49165 -41210
rect -49485 -41864 -49479 -41236
rect -49171 -41864 -49165 -41236
rect -49485 -41890 -49165 -41864
rect -74825 -41896 -48825 -41890
rect -74825 -42204 -74819 -41896
rect -74511 -41928 -74139 -41896
rect -74511 -42172 -74447 -41928
rect -74203 -42172 -74139 -41928
rect -74511 -42204 -74139 -42172
rect -73511 -41928 -73139 -41896
rect -73511 -42172 -73447 -41928
rect -73203 -42172 -73139 -41928
rect -73511 -42204 -73139 -42172
rect -72511 -41928 -72139 -41896
rect -72511 -42172 -72447 -41928
rect -72203 -42172 -72139 -41928
rect -72511 -42204 -72139 -42172
rect -71511 -41928 -71139 -41896
rect -71511 -42172 -71447 -41928
rect -71203 -42172 -71139 -41928
rect -71511 -42204 -71139 -42172
rect -70511 -41928 -70139 -41896
rect -70511 -42172 -70447 -41928
rect -70203 -42172 -70139 -41928
rect -70511 -42204 -70139 -42172
rect -69511 -41928 -69139 -41896
rect -69511 -42172 -69447 -41928
rect -69203 -42172 -69139 -41928
rect -69511 -42204 -69139 -42172
rect -68511 -41928 -68139 -41896
rect -68511 -42172 -68447 -41928
rect -68203 -42172 -68139 -41928
rect -68511 -42204 -68139 -42172
rect -67511 -41928 -67139 -41896
rect -67511 -42172 -67447 -41928
rect -67203 -42172 -67139 -41928
rect -67511 -42204 -67139 -42172
rect -66511 -41928 -66139 -41896
rect -66511 -42172 -66447 -41928
rect -66203 -42172 -66139 -41928
rect -66511 -42204 -66139 -42172
rect -65511 -41928 -65139 -41896
rect -65511 -42172 -65447 -41928
rect -65203 -42172 -65139 -41928
rect -65511 -42204 -65139 -42172
rect -64511 -41928 -64139 -41896
rect -64511 -42172 -64447 -41928
rect -64203 -42172 -64139 -41928
rect -64511 -42204 -64139 -42172
rect -63511 -41928 -63139 -41896
rect -63511 -42172 -63447 -41928
rect -63203 -42172 -63139 -41928
rect -63511 -42204 -63139 -42172
rect -62511 -41928 -62139 -41896
rect -62511 -42172 -62447 -41928
rect -62203 -42172 -62139 -41928
rect -62511 -42204 -62139 -42172
rect -61511 -41928 -61139 -41896
rect -61511 -42172 -61447 -41928
rect -61203 -42172 -61139 -41928
rect -61511 -42204 -61139 -42172
rect -60511 -41928 -60139 -41896
rect -60511 -42172 -60447 -41928
rect -60203 -42172 -60139 -41928
rect -60511 -42204 -60139 -42172
rect -59511 -41928 -59139 -41896
rect -59511 -42172 -59447 -41928
rect -59203 -42172 -59139 -41928
rect -59511 -42204 -59139 -42172
rect -58511 -41928 -58139 -41896
rect -58511 -42172 -58447 -41928
rect -58203 -42172 -58139 -41928
rect -58511 -42204 -58139 -42172
rect -57511 -41928 -57139 -41896
rect -57511 -42172 -57447 -41928
rect -57203 -42172 -57139 -41928
rect -57511 -42204 -57139 -42172
rect -56511 -41928 -56139 -41896
rect -56511 -42172 -56447 -41928
rect -56203 -42172 -56139 -41928
rect -56511 -42204 -56139 -42172
rect -55511 -41928 -55139 -41896
rect -55511 -42172 -55447 -41928
rect -55203 -42172 -55139 -41928
rect -55511 -42204 -55139 -42172
rect -54511 -41928 -54139 -41896
rect -54511 -42172 -54447 -41928
rect -54203 -42172 -54139 -41928
rect -54511 -42204 -54139 -42172
rect -53511 -41928 -53139 -41896
rect -53511 -42172 -53447 -41928
rect -53203 -42172 -53139 -41928
rect -53511 -42204 -53139 -42172
rect -52511 -41928 -52139 -41896
rect -52511 -42172 -52447 -41928
rect -52203 -42172 -52139 -41928
rect -52511 -42204 -52139 -42172
rect -51511 -41928 -51139 -41896
rect -51511 -42172 -51447 -41928
rect -51203 -42172 -51139 -41928
rect -51511 -42204 -51139 -42172
rect -50511 -41928 -50139 -41896
rect -50511 -42172 -50447 -41928
rect -50203 -42172 -50139 -41928
rect -50511 -42204 -50139 -42172
rect -49511 -41928 -49139 -41896
rect -49511 -42172 -49447 -41928
rect -49203 -42172 -49139 -41928
rect -49511 -42204 -49139 -42172
rect -48831 -42204 -48825 -41896
rect -74825 -42210 -48825 -42204
rect -74485 -42236 -74165 -42210
rect -74485 -42864 -74479 -42236
rect -74171 -42864 -74165 -42236
rect -74485 -42890 -74165 -42864
rect -73485 -42236 -73165 -42210
rect -73485 -42864 -73479 -42236
rect -73171 -42864 -73165 -42236
rect -73485 -42890 -73165 -42864
rect -72485 -42236 -72165 -42210
rect -72485 -42864 -72479 -42236
rect -72171 -42864 -72165 -42236
rect -72485 -42890 -72165 -42864
rect -71485 -42236 -71165 -42210
rect -71485 -42864 -71479 -42236
rect -71171 -42864 -71165 -42236
rect -71485 -42890 -71165 -42864
rect -70485 -42236 -70165 -42210
rect -70485 -42864 -70479 -42236
rect -70171 -42864 -70165 -42236
rect -70485 -42890 -70165 -42864
rect -69485 -42236 -69165 -42210
rect -69485 -42864 -69479 -42236
rect -69171 -42864 -69165 -42236
rect -69485 -42890 -69165 -42864
rect -68485 -42236 -68165 -42210
rect -68485 -42864 -68479 -42236
rect -68171 -42864 -68165 -42236
rect -68485 -42890 -68165 -42864
rect -67485 -42236 -67165 -42210
rect -67485 -42864 -67479 -42236
rect -67171 -42864 -67165 -42236
rect -67485 -42890 -67165 -42864
rect -66485 -42236 -66165 -42210
rect -66485 -42864 -66479 -42236
rect -66171 -42864 -66165 -42236
rect -66485 -42890 -66165 -42864
rect -65485 -42236 -65165 -42210
rect -65485 -42864 -65479 -42236
rect -65171 -42864 -65165 -42236
rect -65485 -42890 -65165 -42864
rect -64485 -42236 -64165 -42210
rect -64485 -42864 -64479 -42236
rect -64171 -42864 -64165 -42236
rect -64485 -42890 -64165 -42864
rect -63485 -42236 -63165 -42210
rect -63485 -42864 -63479 -42236
rect -63171 -42864 -63165 -42236
rect -63485 -42890 -63165 -42864
rect -62485 -42236 -62165 -42210
rect -62485 -42864 -62479 -42236
rect -62171 -42864 -62165 -42236
rect -62485 -42890 -62165 -42864
rect -61485 -42236 -61165 -42210
rect -61485 -42864 -61479 -42236
rect -61171 -42864 -61165 -42236
rect -61485 -42890 -61165 -42864
rect -60485 -42236 -60165 -42210
rect -60485 -42864 -60479 -42236
rect -60171 -42864 -60165 -42236
rect -60485 -42890 -60165 -42864
rect -59485 -42236 -59165 -42210
rect -59485 -42864 -59479 -42236
rect -59171 -42864 -59165 -42236
rect -59485 -42890 -59165 -42864
rect -58485 -42236 -58165 -42210
rect -58485 -42864 -58479 -42236
rect -58171 -42864 -58165 -42236
rect -58485 -42890 -58165 -42864
rect -57485 -42236 -57165 -42210
rect -57485 -42864 -57479 -42236
rect -57171 -42864 -57165 -42236
rect -57485 -42890 -57165 -42864
rect -56485 -42236 -56165 -42210
rect -56485 -42864 -56479 -42236
rect -56171 -42864 -56165 -42236
rect -56485 -42890 -56165 -42864
rect -55485 -42236 -55165 -42210
rect -55485 -42864 -55479 -42236
rect -55171 -42864 -55165 -42236
rect -55485 -42890 -55165 -42864
rect -54485 -42236 -54165 -42210
rect -54485 -42864 -54479 -42236
rect -54171 -42864 -54165 -42236
rect -54485 -42890 -54165 -42864
rect -53485 -42236 -53165 -42210
rect -53485 -42864 -53479 -42236
rect -53171 -42864 -53165 -42236
rect -53485 -42890 -53165 -42864
rect -52485 -42236 -52165 -42210
rect -52485 -42864 -52479 -42236
rect -52171 -42864 -52165 -42236
rect -52485 -42890 -52165 -42864
rect -51485 -42236 -51165 -42210
rect -51485 -42864 -51479 -42236
rect -51171 -42864 -51165 -42236
rect -51485 -42890 -51165 -42864
rect -50485 -42236 -50165 -42210
rect -50485 -42864 -50479 -42236
rect -50171 -42864 -50165 -42236
rect -50485 -42890 -50165 -42864
rect -49485 -42236 -49165 -42210
rect -49485 -42864 -49479 -42236
rect -49171 -42864 -49165 -42236
rect -49485 -42890 -49165 -42864
rect -74825 -42896 -48825 -42890
rect -74825 -43204 -74819 -42896
rect -74511 -42928 -74139 -42896
rect -74511 -43172 -74447 -42928
rect -74203 -43172 -74139 -42928
rect -74511 -43204 -74139 -43172
rect -73511 -42928 -73139 -42896
rect -73511 -43172 -73447 -42928
rect -73203 -43172 -73139 -42928
rect -73511 -43204 -73139 -43172
rect -72511 -42928 -72139 -42896
rect -72511 -43172 -72447 -42928
rect -72203 -43172 -72139 -42928
rect -72511 -43204 -72139 -43172
rect -71511 -42928 -71139 -42896
rect -71511 -43172 -71447 -42928
rect -71203 -43172 -71139 -42928
rect -71511 -43204 -71139 -43172
rect -70511 -42928 -70139 -42896
rect -70511 -43172 -70447 -42928
rect -70203 -43172 -70139 -42928
rect -70511 -43204 -70139 -43172
rect -69511 -42928 -69139 -42896
rect -69511 -43172 -69447 -42928
rect -69203 -43172 -69139 -42928
rect -69511 -43204 -69139 -43172
rect -68511 -42928 -68139 -42896
rect -68511 -43172 -68447 -42928
rect -68203 -43172 -68139 -42928
rect -68511 -43204 -68139 -43172
rect -67511 -42928 -67139 -42896
rect -67511 -43172 -67447 -42928
rect -67203 -43172 -67139 -42928
rect -67511 -43204 -67139 -43172
rect -66511 -42928 -66139 -42896
rect -66511 -43172 -66447 -42928
rect -66203 -43172 -66139 -42928
rect -66511 -43204 -66139 -43172
rect -65511 -42928 -65139 -42896
rect -65511 -43172 -65447 -42928
rect -65203 -43172 -65139 -42928
rect -65511 -43204 -65139 -43172
rect -64511 -42928 -64139 -42896
rect -64511 -43172 -64447 -42928
rect -64203 -43172 -64139 -42928
rect -64511 -43204 -64139 -43172
rect -63511 -42928 -63139 -42896
rect -63511 -43172 -63447 -42928
rect -63203 -43172 -63139 -42928
rect -63511 -43204 -63139 -43172
rect -62511 -42928 -62139 -42896
rect -62511 -43172 -62447 -42928
rect -62203 -43172 -62139 -42928
rect -62511 -43204 -62139 -43172
rect -61511 -42928 -61139 -42896
rect -61511 -43172 -61447 -42928
rect -61203 -43172 -61139 -42928
rect -61511 -43204 -61139 -43172
rect -60511 -42928 -60139 -42896
rect -60511 -43172 -60447 -42928
rect -60203 -43172 -60139 -42928
rect -60511 -43204 -60139 -43172
rect -59511 -42928 -59139 -42896
rect -59511 -43172 -59447 -42928
rect -59203 -43172 -59139 -42928
rect -59511 -43204 -59139 -43172
rect -58511 -42928 -58139 -42896
rect -58511 -43172 -58447 -42928
rect -58203 -43172 -58139 -42928
rect -58511 -43204 -58139 -43172
rect -57511 -42928 -57139 -42896
rect -57511 -43172 -57447 -42928
rect -57203 -43172 -57139 -42928
rect -57511 -43204 -57139 -43172
rect -56511 -42928 -56139 -42896
rect -56511 -43172 -56447 -42928
rect -56203 -43172 -56139 -42928
rect -56511 -43204 -56139 -43172
rect -55511 -42928 -55139 -42896
rect -55511 -43172 -55447 -42928
rect -55203 -43172 -55139 -42928
rect -55511 -43204 -55139 -43172
rect -54511 -42928 -54139 -42896
rect -54511 -43172 -54447 -42928
rect -54203 -43172 -54139 -42928
rect -54511 -43204 -54139 -43172
rect -53511 -42928 -53139 -42896
rect -53511 -43172 -53447 -42928
rect -53203 -43172 -53139 -42928
rect -53511 -43204 -53139 -43172
rect -52511 -42928 -52139 -42896
rect -52511 -43172 -52447 -42928
rect -52203 -43172 -52139 -42928
rect -52511 -43204 -52139 -43172
rect -51511 -42928 -51139 -42896
rect -51511 -43172 -51447 -42928
rect -51203 -43172 -51139 -42928
rect -51511 -43204 -51139 -43172
rect -50511 -42928 -50139 -42896
rect -50511 -43172 -50447 -42928
rect -50203 -43172 -50139 -42928
rect -50511 -43204 -50139 -43172
rect -49511 -42928 -49139 -42896
rect -49511 -43172 -49447 -42928
rect -49203 -43172 -49139 -42928
rect -49511 -43204 -49139 -43172
rect -48831 -43204 -48825 -42896
rect -74825 -43210 -48825 -43204
rect -74485 -43236 -74165 -43210
rect -74485 -43864 -74479 -43236
rect -74171 -43864 -74165 -43236
rect -74485 -43890 -74165 -43864
rect -73485 -43236 -73165 -43210
rect -73485 -43864 -73479 -43236
rect -73171 -43864 -73165 -43236
rect -73485 -43890 -73165 -43864
rect -72485 -43236 -72165 -43210
rect -72485 -43864 -72479 -43236
rect -72171 -43864 -72165 -43236
rect -72485 -43890 -72165 -43864
rect -71485 -43236 -71165 -43210
rect -71485 -43864 -71479 -43236
rect -71171 -43864 -71165 -43236
rect -71485 -43890 -71165 -43864
rect -70485 -43236 -70165 -43210
rect -70485 -43864 -70479 -43236
rect -70171 -43864 -70165 -43236
rect -70485 -43890 -70165 -43864
rect -69485 -43236 -69165 -43210
rect -69485 -43864 -69479 -43236
rect -69171 -43864 -69165 -43236
rect -69485 -43890 -69165 -43864
rect -68485 -43236 -68165 -43210
rect -68485 -43864 -68479 -43236
rect -68171 -43864 -68165 -43236
rect -68485 -43890 -68165 -43864
rect -67485 -43236 -67165 -43210
rect -67485 -43864 -67479 -43236
rect -67171 -43864 -67165 -43236
rect -67485 -43890 -67165 -43864
rect -66485 -43236 -66165 -43210
rect -66485 -43864 -66479 -43236
rect -66171 -43864 -66165 -43236
rect -66485 -43890 -66165 -43864
rect -65485 -43236 -65165 -43210
rect -65485 -43864 -65479 -43236
rect -65171 -43864 -65165 -43236
rect -65485 -43890 -65165 -43864
rect -64485 -43236 -64165 -43210
rect -64485 -43864 -64479 -43236
rect -64171 -43864 -64165 -43236
rect -64485 -43890 -64165 -43864
rect -63485 -43236 -63165 -43210
rect -63485 -43864 -63479 -43236
rect -63171 -43864 -63165 -43236
rect -63485 -43890 -63165 -43864
rect -62485 -43236 -62165 -43210
rect -62485 -43864 -62479 -43236
rect -62171 -43864 -62165 -43236
rect -62485 -43890 -62165 -43864
rect -61485 -43236 -61165 -43210
rect -61485 -43864 -61479 -43236
rect -61171 -43864 -61165 -43236
rect -61485 -43890 -61165 -43864
rect -60485 -43236 -60165 -43210
rect -60485 -43864 -60479 -43236
rect -60171 -43864 -60165 -43236
rect -60485 -43890 -60165 -43864
rect -59485 -43236 -59165 -43210
rect -59485 -43864 -59479 -43236
rect -59171 -43864 -59165 -43236
rect -59485 -43890 -59165 -43864
rect -58485 -43236 -58165 -43210
rect -58485 -43864 -58479 -43236
rect -58171 -43864 -58165 -43236
rect -58485 -43890 -58165 -43864
rect -57485 -43236 -57165 -43210
rect -57485 -43864 -57479 -43236
rect -57171 -43864 -57165 -43236
rect -57485 -43890 -57165 -43864
rect -56485 -43236 -56165 -43210
rect -56485 -43864 -56479 -43236
rect -56171 -43864 -56165 -43236
rect -56485 -43890 -56165 -43864
rect -55485 -43236 -55165 -43210
rect -55485 -43864 -55479 -43236
rect -55171 -43864 -55165 -43236
rect -55485 -43890 -55165 -43864
rect -54485 -43236 -54165 -43210
rect -54485 -43864 -54479 -43236
rect -54171 -43864 -54165 -43236
rect -54485 -43890 -54165 -43864
rect -53485 -43236 -53165 -43210
rect -53485 -43864 -53479 -43236
rect -53171 -43864 -53165 -43236
rect -53485 -43890 -53165 -43864
rect -52485 -43236 -52165 -43210
rect -52485 -43864 -52479 -43236
rect -52171 -43864 -52165 -43236
rect -52485 -43890 -52165 -43864
rect -51485 -43236 -51165 -43210
rect -51485 -43864 -51479 -43236
rect -51171 -43864 -51165 -43236
rect -51485 -43890 -51165 -43864
rect -50485 -43236 -50165 -43210
rect -50485 -43864 -50479 -43236
rect -50171 -43864 -50165 -43236
rect -50485 -43890 -50165 -43864
rect -49485 -43236 -49165 -43210
rect -49485 -43864 -49479 -43236
rect -49171 -43864 -49165 -43236
rect -49485 -43890 -49165 -43864
rect -74825 -43896 -48825 -43890
rect -74825 -44204 -74819 -43896
rect -74511 -43928 -74139 -43896
rect -74511 -44172 -74447 -43928
rect -74203 -44172 -74139 -43928
rect -74511 -44204 -74139 -44172
rect -73511 -43928 -73139 -43896
rect -73511 -44172 -73447 -43928
rect -73203 -44172 -73139 -43928
rect -73511 -44204 -73139 -44172
rect -72511 -43928 -72139 -43896
rect -72511 -44172 -72447 -43928
rect -72203 -44172 -72139 -43928
rect -72511 -44204 -72139 -44172
rect -71511 -43928 -71139 -43896
rect -71511 -44172 -71447 -43928
rect -71203 -44172 -71139 -43928
rect -71511 -44204 -71139 -44172
rect -70511 -43928 -70139 -43896
rect -70511 -44172 -70447 -43928
rect -70203 -44172 -70139 -43928
rect -70511 -44204 -70139 -44172
rect -69511 -43928 -69139 -43896
rect -69511 -44172 -69447 -43928
rect -69203 -44172 -69139 -43928
rect -69511 -44204 -69139 -44172
rect -68511 -43928 -68139 -43896
rect -68511 -44172 -68447 -43928
rect -68203 -44172 -68139 -43928
rect -68511 -44204 -68139 -44172
rect -67511 -43928 -67139 -43896
rect -67511 -44172 -67447 -43928
rect -67203 -44172 -67139 -43928
rect -67511 -44204 -67139 -44172
rect -66511 -43928 -66139 -43896
rect -66511 -44172 -66447 -43928
rect -66203 -44172 -66139 -43928
rect -66511 -44204 -66139 -44172
rect -65511 -43928 -65139 -43896
rect -65511 -44172 -65447 -43928
rect -65203 -44172 -65139 -43928
rect -65511 -44204 -65139 -44172
rect -64511 -43928 -64139 -43896
rect -64511 -44172 -64447 -43928
rect -64203 -44172 -64139 -43928
rect -64511 -44204 -64139 -44172
rect -63511 -43928 -63139 -43896
rect -63511 -44172 -63447 -43928
rect -63203 -44172 -63139 -43928
rect -63511 -44204 -63139 -44172
rect -62511 -43928 -62139 -43896
rect -62511 -44172 -62447 -43928
rect -62203 -44172 -62139 -43928
rect -62511 -44204 -62139 -44172
rect -61511 -43928 -61139 -43896
rect -61511 -44172 -61447 -43928
rect -61203 -44172 -61139 -43928
rect -61511 -44204 -61139 -44172
rect -60511 -43928 -60139 -43896
rect -60511 -44172 -60447 -43928
rect -60203 -44172 -60139 -43928
rect -60511 -44204 -60139 -44172
rect -59511 -43928 -59139 -43896
rect -59511 -44172 -59447 -43928
rect -59203 -44172 -59139 -43928
rect -59511 -44204 -59139 -44172
rect -58511 -43928 -58139 -43896
rect -58511 -44172 -58447 -43928
rect -58203 -44172 -58139 -43928
rect -58511 -44204 -58139 -44172
rect -57511 -43928 -57139 -43896
rect -57511 -44172 -57447 -43928
rect -57203 -44172 -57139 -43928
rect -57511 -44204 -57139 -44172
rect -56511 -43928 -56139 -43896
rect -56511 -44172 -56447 -43928
rect -56203 -44172 -56139 -43928
rect -56511 -44204 -56139 -44172
rect -55511 -43928 -55139 -43896
rect -55511 -44172 -55447 -43928
rect -55203 -44172 -55139 -43928
rect -55511 -44204 -55139 -44172
rect -54511 -43928 -54139 -43896
rect -54511 -44172 -54447 -43928
rect -54203 -44172 -54139 -43928
rect -54511 -44204 -54139 -44172
rect -53511 -43928 -53139 -43896
rect -53511 -44172 -53447 -43928
rect -53203 -44172 -53139 -43928
rect -53511 -44204 -53139 -44172
rect -52511 -43928 -52139 -43896
rect -52511 -44172 -52447 -43928
rect -52203 -44172 -52139 -43928
rect -52511 -44204 -52139 -44172
rect -51511 -43928 -51139 -43896
rect -51511 -44172 -51447 -43928
rect -51203 -44172 -51139 -43928
rect -51511 -44204 -51139 -44172
rect -50511 -43928 -50139 -43896
rect -50511 -44172 -50447 -43928
rect -50203 -44172 -50139 -43928
rect -50511 -44204 -50139 -44172
rect -49511 -43928 -49139 -43896
rect -49511 -44172 -49447 -43928
rect -49203 -44172 -49139 -43928
rect -49511 -44204 -49139 -44172
rect -48831 -44204 -48825 -43896
rect -74825 -44210 -48825 -44204
rect -74485 -44236 -74165 -44210
rect -74485 -44864 -74479 -44236
rect -74171 -44864 -74165 -44236
rect -74485 -44890 -74165 -44864
rect -73485 -44236 -73165 -44210
rect -73485 -44864 -73479 -44236
rect -73171 -44864 -73165 -44236
rect -73485 -44890 -73165 -44864
rect -72485 -44236 -72165 -44210
rect -72485 -44864 -72479 -44236
rect -72171 -44864 -72165 -44236
rect -72485 -44890 -72165 -44864
rect -71485 -44236 -71165 -44210
rect -71485 -44864 -71479 -44236
rect -71171 -44864 -71165 -44236
rect -71485 -44890 -71165 -44864
rect -70485 -44236 -70165 -44210
rect -70485 -44864 -70479 -44236
rect -70171 -44864 -70165 -44236
rect -70485 -44890 -70165 -44864
rect -69485 -44236 -69165 -44210
rect -69485 -44864 -69479 -44236
rect -69171 -44864 -69165 -44236
rect -69485 -44890 -69165 -44864
rect -68485 -44236 -68165 -44210
rect -68485 -44864 -68479 -44236
rect -68171 -44864 -68165 -44236
rect -68485 -44890 -68165 -44864
rect -67485 -44236 -67165 -44210
rect -67485 -44864 -67479 -44236
rect -67171 -44864 -67165 -44236
rect -67485 -44890 -67165 -44864
rect -66485 -44236 -66165 -44210
rect -66485 -44864 -66479 -44236
rect -66171 -44864 -66165 -44236
rect -66485 -44890 -66165 -44864
rect -65485 -44236 -65165 -44210
rect -65485 -44864 -65479 -44236
rect -65171 -44864 -65165 -44236
rect -65485 -44890 -65165 -44864
rect -64485 -44236 -64165 -44210
rect -64485 -44864 -64479 -44236
rect -64171 -44864 -64165 -44236
rect -64485 -44890 -64165 -44864
rect -63485 -44236 -63165 -44210
rect -63485 -44864 -63479 -44236
rect -63171 -44864 -63165 -44236
rect -63485 -44890 -63165 -44864
rect -62485 -44236 -62165 -44210
rect -62485 -44864 -62479 -44236
rect -62171 -44864 -62165 -44236
rect -62485 -44890 -62165 -44864
rect -61485 -44236 -61165 -44210
rect -61485 -44864 -61479 -44236
rect -61171 -44864 -61165 -44236
rect -61485 -44890 -61165 -44864
rect -60485 -44236 -60165 -44210
rect -60485 -44864 -60479 -44236
rect -60171 -44864 -60165 -44236
rect -60485 -44890 -60165 -44864
rect -59485 -44236 -59165 -44210
rect -59485 -44864 -59479 -44236
rect -59171 -44864 -59165 -44236
rect -59485 -44890 -59165 -44864
rect -58485 -44236 -58165 -44210
rect -58485 -44864 -58479 -44236
rect -58171 -44864 -58165 -44236
rect -58485 -44890 -58165 -44864
rect -57485 -44236 -57165 -44210
rect -57485 -44864 -57479 -44236
rect -57171 -44864 -57165 -44236
rect -57485 -44890 -57165 -44864
rect -56485 -44236 -56165 -44210
rect -56485 -44864 -56479 -44236
rect -56171 -44864 -56165 -44236
rect -56485 -44890 -56165 -44864
rect -55485 -44236 -55165 -44210
rect -55485 -44864 -55479 -44236
rect -55171 -44864 -55165 -44236
rect -55485 -44890 -55165 -44864
rect -54485 -44236 -54165 -44210
rect -54485 -44864 -54479 -44236
rect -54171 -44864 -54165 -44236
rect -54485 -44890 -54165 -44864
rect -53485 -44236 -53165 -44210
rect -53485 -44864 -53479 -44236
rect -53171 -44864 -53165 -44236
rect -53485 -44890 -53165 -44864
rect -52485 -44236 -52165 -44210
rect -52485 -44864 -52479 -44236
rect -52171 -44864 -52165 -44236
rect -52485 -44890 -52165 -44864
rect -51485 -44236 -51165 -44210
rect -51485 -44864 -51479 -44236
rect -51171 -44864 -51165 -44236
rect -51485 -44890 -51165 -44864
rect -50485 -44236 -50165 -44210
rect -50485 -44864 -50479 -44236
rect -50171 -44864 -50165 -44236
rect -50485 -44890 -50165 -44864
rect -49485 -44236 -49165 -44210
rect -49485 -44864 -49479 -44236
rect -49171 -44864 -49165 -44236
rect -46275 -44496 -46234 -32604
rect -36326 -33850 -27875 -32604
rect -12675 -32604 5725 -32550
rect -12675 -33850 -4234 -32604
rect -36326 -35350 -4234 -33850
rect -36326 -36150 -27875 -35350
rect -12675 -36150 -4234 -35350
rect -36326 -37650 -4234 -36150
rect -36326 -38450 -27875 -37650
rect -12675 -38450 -4234 -37650
rect -36326 -39950 -4234 -38450
rect -36326 -40750 -27875 -39950
rect -12675 -40750 -4234 -39950
rect -36326 -42250 -4234 -40750
rect -36326 -43050 -27875 -42250
rect -12675 -43050 -4234 -42250
rect -36326 -44496 -4234 -43050
rect 5674 -44496 5725 -32604
rect 8615 -32864 8621 -32236
rect 8929 -32864 8935 -32236
rect 8615 -32890 8935 -32864
rect 9615 -32236 9935 -32210
rect 9615 -32864 9621 -32236
rect 9929 -32864 9935 -32236
rect 9615 -32890 9935 -32864
rect 10615 -32236 10935 -32210
rect 10615 -32864 10621 -32236
rect 10929 -32864 10935 -32236
rect 10615 -32890 10935 -32864
rect 11615 -32236 11935 -32210
rect 11615 -32864 11621 -32236
rect 11929 -32864 11935 -32236
rect 11615 -32890 11935 -32864
rect 12615 -32236 12935 -32210
rect 12615 -32864 12621 -32236
rect 12929 -32864 12935 -32236
rect 12615 -32890 12935 -32864
rect 13615 -32236 13935 -32210
rect 13615 -32864 13621 -32236
rect 13929 -32864 13935 -32236
rect 13615 -32890 13935 -32864
rect 14615 -32236 14935 -32210
rect 14615 -32864 14621 -32236
rect 14929 -32864 14935 -32236
rect 14615 -32890 14935 -32864
rect 15615 -32236 15935 -32210
rect 15615 -32864 15621 -32236
rect 15929 -32864 15935 -32236
rect 15615 -32890 15935 -32864
rect 16615 -32236 16935 -32210
rect 16615 -32864 16621 -32236
rect 16929 -32864 16935 -32236
rect 16615 -32890 16935 -32864
rect 17615 -32236 17935 -32210
rect 17615 -32864 17621 -32236
rect 17929 -32864 17935 -32236
rect 17615 -32890 17935 -32864
rect 18615 -32236 18935 -32210
rect 18615 -32864 18621 -32236
rect 18929 -32864 18935 -32236
rect 18615 -32890 18935 -32864
rect 19615 -32236 19935 -32210
rect 19615 -32864 19621 -32236
rect 19929 -32864 19935 -32236
rect 19615 -32890 19935 -32864
rect 20615 -32236 20935 -32210
rect 20615 -32864 20621 -32236
rect 20929 -32864 20935 -32236
rect 20615 -32890 20935 -32864
rect 21615 -32236 21935 -32210
rect 21615 -32864 21621 -32236
rect 21929 -32864 21935 -32236
rect 21615 -32890 21935 -32864
rect 22615 -32236 22935 -32210
rect 22615 -32864 22621 -32236
rect 22929 -32864 22935 -32236
rect 22615 -32890 22935 -32864
rect 23615 -32236 23935 -32210
rect 23615 -32864 23621 -32236
rect 23929 -32864 23935 -32236
rect 23615 -32890 23935 -32864
rect 24615 -32236 24935 -32210
rect 24615 -32864 24621 -32236
rect 24929 -32864 24935 -32236
rect 24615 -32890 24935 -32864
rect 25615 -32236 25935 -32210
rect 25615 -32864 25621 -32236
rect 25929 -32864 25935 -32236
rect 25615 -32890 25935 -32864
rect 26615 -32236 26935 -32210
rect 26615 -32864 26621 -32236
rect 26929 -32864 26935 -32236
rect 26615 -32890 26935 -32864
rect 27615 -32236 27935 -32210
rect 27615 -32864 27621 -32236
rect 27929 -32864 27935 -32236
rect 27615 -32890 27935 -32864
rect 28615 -32236 28935 -32210
rect 28615 -32864 28621 -32236
rect 28929 -32864 28935 -32236
rect 28615 -32890 28935 -32864
rect 29615 -32236 29935 -32210
rect 29615 -32864 29621 -32236
rect 29929 -32864 29935 -32236
rect 29615 -32890 29935 -32864
rect 30615 -32236 30935 -32210
rect 30615 -32864 30621 -32236
rect 30929 -32864 30935 -32236
rect 30615 -32890 30935 -32864
rect 31615 -32236 31935 -32210
rect 31615 -32864 31621 -32236
rect 31929 -32864 31935 -32236
rect 31615 -32890 31935 -32864
rect 32615 -32236 32935 -32210
rect 32615 -32864 32621 -32236
rect 32929 -32864 32935 -32236
rect 32615 -32890 32935 -32864
rect 33615 -32236 33935 -32210
rect 33615 -32864 33621 -32236
rect 33929 -32864 33935 -32236
rect 33615 -32890 33935 -32864
rect 8275 -32896 34275 -32890
rect 8275 -33204 8281 -32896
rect 8589 -32928 8961 -32896
rect 8589 -33172 8653 -32928
rect 8897 -33172 8961 -32928
rect 8589 -33204 8961 -33172
rect 9589 -32928 9961 -32896
rect 9589 -33172 9653 -32928
rect 9897 -33172 9961 -32928
rect 9589 -33204 9961 -33172
rect 10589 -32928 10961 -32896
rect 10589 -33172 10653 -32928
rect 10897 -33172 10961 -32928
rect 10589 -33204 10961 -33172
rect 11589 -32928 11961 -32896
rect 11589 -33172 11653 -32928
rect 11897 -33172 11961 -32928
rect 11589 -33204 11961 -33172
rect 12589 -32928 12961 -32896
rect 12589 -33172 12653 -32928
rect 12897 -33172 12961 -32928
rect 12589 -33204 12961 -33172
rect 13589 -32928 13961 -32896
rect 13589 -33172 13653 -32928
rect 13897 -33172 13961 -32928
rect 13589 -33204 13961 -33172
rect 14589 -32928 14961 -32896
rect 14589 -33172 14653 -32928
rect 14897 -33172 14961 -32928
rect 14589 -33204 14961 -33172
rect 15589 -32928 15961 -32896
rect 15589 -33172 15653 -32928
rect 15897 -33172 15961 -32928
rect 15589 -33204 15961 -33172
rect 16589 -32928 16961 -32896
rect 16589 -33172 16653 -32928
rect 16897 -33172 16961 -32928
rect 16589 -33204 16961 -33172
rect 17589 -32928 17961 -32896
rect 17589 -33172 17653 -32928
rect 17897 -33172 17961 -32928
rect 17589 -33204 17961 -33172
rect 18589 -32928 18961 -32896
rect 18589 -33172 18653 -32928
rect 18897 -33172 18961 -32928
rect 18589 -33204 18961 -33172
rect 19589 -32928 19961 -32896
rect 19589 -33172 19653 -32928
rect 19897 -33172 19961 -32928
rect 19589 -33204 19961 -33172
rect 20589 -32928 20961 -32896
rect 20589 -33172 20653 -32928
rect 20897 -33172 20961 -32928
rect 20589 -33204 20961 -33172
rect 21589 -32928 21961 -32896
rect 21589 -33172 21653 -32928
rect 21897 -33172 21961 -32928
rect 21589 -33204 21961 -33172
rect 22589 -32928 22961 -32896
rect 22589 -33172 22653 -32928
rect 22897 -33172 22961 -32928
rect 22589 -33204 22961 -33172
rect 23589 -32928 23961 -32896
rect 23589 -33172 23653 -32928
rect 23897 -33172 23961 -32928
rect 23589 -33204 23961 -33172
rect 24589 -32928 24961 -32896
rect 24589 -33172 24653 -32928
rect 24897 -33172 24961 -32928
rect 24589 -33204 24961 -33172
rect 25589 -32928 25961 -32896
rect 25589 -33172 25653 -32928
rect 25897 -33172 25961 -32928
rect 25589 -33204 25961 -33172
rect 26589 -32928 26961 -32896
rect 26589 -33172 26653 -32928
rect 26897 -33172 26961 -32928
rect 26589 -33204 26961 -33172
rect 27589 -32928 27961 -32896
rect 27589 -33172 27653 -32928
rect 27897 -33172 27961 -32928
rect 27589 -33204 27961 -33172
rect 28589 -32928 28961 -32896
rect 28589 -33172 28653 -32928
rect 28897 -33172 28961 -32928
rect 28589 -33204 28961 -33172
rect 29589 -32928 29961 -32896
rect 29589 -33172 29653 -32928
rect 29897 -33172 29961 -32928
rect 29589 -33204 29961 -33172
rect 30589 -32928 30961 -32896
rect 30589 -33172 30653 -32928
rect 30897 -33172 30961 -32928
rect 30589 -33204 30961 -33172
rect 31589 -32928 31961 -32896
rect 31589 -33172 31653 -32928
rect 31897 -33172 31961 -32928
rect 31589 -33204 31961 -33172
rect 32589 -32928 32961 -32896
rect 32589 -33172 32653 -32928
rect 32897 -33172 32961 -32928
rect 32589 -33204 32961 -33172
rect 33589 -32928 33961 -32896
rect 33589 -33172 33653 -32928
rect 33897 -33172 33961 -32928
rect 33589 -33204 33961 -33172
rect 34269 -33204 34275 -32896
rect 8275 -33210 34275 -33204
rect 8615 -33236 8935 -33210
rect 8615 -33864 8621 -33236
rect 8929 -33864 8935 -33236
rect 8615 -33890 8935 -33864
rect 9615 -33236 9935 -33210
rect 9615 -33864 9621 -33236
rect 9929 -33864 9935 -33236
rect 9615 -33890 9935 -33864
rect 10615 -33236 10935 -33210
rect 10615 -33864 10621 -33236
rect 10929 -33864 10935 -33236
rect 10615 -33890 10935 -33864
rect 11615 -33236 11935 -33210
rect 11615 -33864 11621 -33236
rect 11929 -33864 11935 -33236
rect 11615 -33890 11935 -33864
rect 12615 -33236 12935 -33210
rect 12615 -33864 12621 -33236
rect 12929 -33864 12935 -33236
rect 12615 -33890 12935 -33864
rect 13615 -33236 13935 -33210
rect 13615 -33864 13621 -33236
rect 13929 -33864 13935 -33236
rect 13615 -33890 13935 -33864
rect 14615 -33236 14935 -33210
rect 14615 -33864 14621 -33236
rect 14929 -33864 14935 -33236
rect 14615 -33890 14935 -33864
rect 15615 -33236 15935 -33210
rect 15615 -33864 15621 -33236
rect 15929 -33864 15935 -33236
rect 15615 -33890 15935 -33864
rect 16615 -33236 16935 -33210
rect 16615 -33864 16621 -33236
rect 16929 -33864 16935 -33236
rect 16615 -33890 16935 -33864
rect 17615 -33236 17935 -33210
rect 17615 -33864 17621 -33236
rect 17929 -33864 17935 -33236
rect 17615 -33890 17935 -33864
rect 18615 -33236 18935 -33210
rect 18615 -33864 18621 -33236
rect 18929 -33864 18935 -33236
rect 18615 -33890 18935 -33864
rect 19615 -33236 19935 -33210
rect 19615 -33864 19621 -33236
rect 19929 -33864 19935 -33236
rect 19615 -33890 19935 -33864
rect 20615 -33236 20935 -33210
rect 20615 -33864 20621 -33236
rect 20929 -33864 20935 -33236
rect 20615 -33890 20935 -33864
rect 21615 -33236 21935 -33210
rect 21615 -33864 21621 -33236
rect 21929 -33864 21935 -33236
rect 21615 -33890 21935 -33864
rect 22615 -33236 22935 -33210
rect 22615 -33864 22621 -33236
rect 22929 -33864 22935 -33236
rect 22615 -33890 22935 -33864
rect 23615 -33236 23935 -33210
rect 23615 -33864 23621 -33236
rect 23929 -33864 23935 -33236
rect 23615 -33890 23935 -33864
rect 24615 -33236 24935 -33210
rect 24615 -33864 24621 -33236
rect 24929 -33864 24935 -33236
rect 24615 -33890 24935 -33864
rect 25615 -33236 25935 -33210
rect 25615 -33864 25621 -33236
rect 25929 -33864 25935 -33236
rect 25615 -33890 25935 -33864
rect 26615 -33236 26935 -33210
rect 26615 -33864 26621 -33236
rect 26929 -33864 26935 -33236
rect 26615 -33890 26935 -33864
rect 27615 -33236 27935 -33210
rect 27615 -33864 27621 -33236
rect 27929 -33864 27935 -33236
rect 27615 -33890 27935 -33864
rect 28615 -33236 28935 -33210
rect 28615 -33864 28621 -33236
rect 28929 -33864 28935 -33236
rect 28615 -33890 28935 -33864
rect 29615 -33236 29935 -33210
rect 29615 -33864 29621 -33236
rect 29929 -33864 29935 -33236
rect 29615 -33890 29935 -33864
rect 30615 -33236 30935 -33210
rect 30615 -33864 30621 -33236
rect 30929 -33864 30935 -33236
rect 30615 -33890 30935 -33864
rect 31615 -33236 31935 -33210
rect 31615 -33864 31621 -33236
rect 31929 -33864 31935 -33236
rect 31615 -33890 31935 -33864
rect 32615 -33236 32935 -33210
rect 32615 -33864 32621 -33236
rect 32929 -33864 32935 -33236
rect 32615 -33890 32935 -33864
rect 33615 -33236 33935 -33210
rect 33615 -33864 33621 -33236
rect 33929 -33864 33935 -33236
rect 33615 -33890 33935 -33864
rect 8275 -33896 34275 -33890
rect 8275 -34204 8281 -33896
rect 8589 -33928 8961 -33896
rect 8589 -34172 8653 -33928
rect 8897 -34172 8961 -33928
rect 8589 -34204 8961 -34172
rect 9589 -33928 9961 -33896
rect 9589 -34172 9653 -33928
rect 9897 -34172 9961 -33928
rect 9589 -34204 9961 -34172
rect 10589 -33928 10961 -33896
rect 10589 -34172 10653 -33928
rect 10897 -34172 10961 -33928
rect 10589 -34204 10961 -34172
rect 11589 -33928 11961 -33896
rect 11589 -34172 11653 -33928
rect 11897 -34172 11961 -33928
rect 11589 -34204 11961 -34172
rect 12589 -33928 12961 -33896
rect 12589 -34172 12653 -33928
rect 12897 -34172 12961 -33928
rect 12589 -34204 12961 -34172
rect 13589 -33928 13961 -33896
rect 13589 -34172 13653 -33928
rect 13897 -34172 13961 -33928
rect 13589 -34204 13961 -34172
rect 14589 -33928 14961 -33896
rect 14589 -34172 14653 -33928
rect 14897 -34172 14961 -33928
rect 14589 -34204 14961 -34172
rect 15589 -33928 15961 -33896
rect 15589 -34172 15653 -33928
rect 15897 -34172 15961 -33928
rect 15589 -34204 15961 -34172
rect 16589 -33928 16961 -33896
rect 16589 -34172 16653 -33928
rect 16897 -34172 16961 -33928
rect 16589 -34204 16961 -34172
rect 17589 -33928 17961 -33896
rect 17589 -34172 17653 -33928
rect 17897 -34172 17961 -33928
rect 17589 -34204 17961 -34172
rect 18589 -33928 18961 -33896
rect 18589 -34172 18653 -33928
rect 18897 -34172 18961 -33928
rect 18589 -34204 18961 -34172
rect 19589 -33928 19961 -33896
rect 19589 -34172 19653 -33928
rect 19897 -34172 19961 -33928
rect 19589 -34204 19961 -34172
rect 20589 -33928 20961 -33896
rect 20589 -34172 20653 -33928
rect 20897 -34172 20961 -33928
rect 20589 -34204 20961 -34172
rect 21589 -33928 21961 -33896
rect 21589 -34172 21653 -33928
rect 21897 -34172 21961 -33928
rect 21589 -34204 21961 -34172
rect 22589 -33928 22961 -33896
rect 22589 -34172 22653 -33928
rect 22897 -34172 22961 -33928
rect 22589 -34204 22961 -34172
rect 23589 -33928 23961 -33896
rect 23589 -34172 23653 -33928
rect 23897 -34172 23961 -33928
rect 23589 -34204 23961 -34172
rect 24589 -33928 24961 -33896
rect 24589 -34172 24653 -33928
rect 24897 -34172 24961 -33928
rect 24589 -34204 24961 -34172
rect 25589 -33928 25961 -33896
rect 25589 -34172 25653 -33928
rect 25897 -34172 25961 -33928
rect 25589 -34204 25961 -34172
rect 26589 -33928 26961 -33896
rect 26589 -34172 26653 -33928
rect 26897 -34172 26961 -33928
rect 26589 -34204 26961 -34172
rect 27589 -33928 27961 -33896
rect 27589 -34172 27653 -33928
rect 27897 -34172 27961 -33928
rect 27589 -34204 27961 -34172
rect 28589 -33928 28961 -33896
rect 28589 -34172 28653 -33928
rect 28897 -34172 28961 -33928
rect 28589 -34204 28961 -34172
rect 29589 -33928 29961 -33896
rect 29589 -34172 29653 -33928
rect 29897 -34172 29961 -33928
rect 29589 -34204 29961 -34172
rect 30589 -33928 30961 -33896
rect 30589 -34172 30653 -33928
rect 30897 -34172 30961 -33928
rect 30589 -34204 30961 -34172
rect 31589 -33928 31961 -33896
rect 31589 -34172 31653 -33928
rect 31897 -34172 31961 -33928
rect 31589 -34204 31961 -34172
rect 32589 -33928 32961 -33896
rect 32589 -34172 32653 -33928
rect 32897 -34172 32961 -33928
rect 32589 -34204 32961 -34172
rect 33589 -33928 33961 -33896
rect 33589 -34172 33653 -33928
rect 33897 -34172 33961 -33928
rect 33589 -34204 33961 -34172
rect 34269 -34204 34275 -33896
rect 8275 -34210 34275 -34204
rect 8615 -34236 8935 -34210
rect 8615 -34864 8621 -34236
rect 8929 -34864 8935 -34236
rect 8615 -34890 8935 -34864
rect 9615 -34236 9935 -34210
rect 9615 -34864 9621 -34236
rect 9929 -34864 9935 -34236
rect 9615 -34890 9935 -34864
rect 10615 -34236 10935 -34210
rect 10615 -34864 10621 -34236
rect 10929 -34864 10935 -34236
rect 10615 -34890 10935 -34864
rect 11615 -34236 11935 -34210
rect 11615 -34864 11621 -34236
rect 11929 -34864 11935 -34236
rect 11615 -34890 11935 -34864
rect 12615 -34236 12935 -34210
rect 12615 -34864 12621 -34236
rect 12929 -34864 12935 -34236
rect 12615 -34890 12935 -34864
rect 13615 -34236 13935 -34210
rect 13615 -34864 13621 -34236
rect 13929 -34864 13935 -34236
rect 13615 -34890 13935 -34864
rect 14615 -34236 14935 -34210
rect 14615 -34864 14621 -34236
rect 14929 -34864 14935 -34236
rect 14615 -34890 14935 -34864
rect 15615 -34236 15935 -34210
rect 15615 -34864 15621 -34236
rect 15929 -34864 15935 -34236
rect 15615 -34890 15935 -34864
rect 16615 -34236 16935 -34210
rect 16615 -34864 16621 -34236
rect 16929 -34864 16935 -34236
rect 16615 -34890 16935 -34864
rect 17615 -34236 17935 -34210
rect 17615 -34864 17621 -34236
rect 17929 -34864 17935 -34236
rect 17615 -34890 17935 -34864
rect 18615 -34236 18935 -34210
rect 18615 -34864 18621 -34236
rect 18929 -34864 18935 -34236
rect 18615 -34890 18935 -34864
rect 19615 -34236 19935 -34210
rect 19615 -34864 19621 -34236
rect 19929 -34864 19935 -34236
rect 19615 -34890 19935 -34864
rect 20615 -34236 20935 -34210
rect 20615 -34864 20621 -34236
rect 20929 -34864 20935 -34236
rect 20615 -34890 20935 -34864
rect 21615 -34236 21935 -34210
rect 21615 -34864 21621 -34236
rect 21929 -34864 21935 -34236
rect 21615 -34890 21935 -34864
rect 22615 -34236 22935 -34210
rect 22615 -34864 22621 -34236
rect 22929 -34864 22935 -34236
rect 22615 -34890 22935 -34864
rect 23615 -34236 23935 -34210
rect 23615 -34864 23621 -34236
rect 23929 -34864 23935 -34236
rect 23615 -34890 23935 -34864
rect 24615 -34236 24935 -34210
rect 24615 -34864 24621 -34236
rect 24929 -34864 24935 -34236
rect 24615 -34890 24935 -34864
rect 25615 -34236 25935 -34210
rect 25615 -34864 25621 -34236
rect 25929 -34864 25935 -34236
rect 25615 -34890 25935 -34864
rect 26615 -34236 26935 -34210
rect 26615 -34864 26621 -34236
rect 26929 -34864 26935 -34236
rect 26615 -34890 26935 -34864
rect 27615 -34236 27935 -34210
rect 27615 -34864 27621 -34236
rect 27929 -34864 27935 -34236
rect 27615 -34890 27935 -34864
rect 28615 -34236 28935 -34210
rect 28615 -34864 28621 -34236
rect 28929 -34864 28935 -34236
rect 28615 -34890 28935 -34864
rect 29615 -34236 29935 -34210
rect 29615 -34864 29621 -34236
rect 29929 -34864 29935 -34236
rect 29615 -34890 29935 -34864
rect 30615 -34236 30935 -34210
rect 30615 -34864 30621 -34236
rect 30929 -34864 30935 -34236
rect 30615 -34890 30935 -34864
rect 31615 -34236 31935 -34210
rect 31615 -34864 31621 -34236
rect 31929 -34864 31935 -34236
rect 31615 -34890 31935 -34864
rect 32615 -34236 32935 -34210
rect 32615 -34864 32621 -34236
rect 32929 -34864 32935 -34236
rect 32615 -34890 32935 -34864
rect 33615 -34236 33935 -34210
rect 33615 -34864 33621 -34236
rect 33929 -34864 33935 -34236
rect 33615 -34890 33935 -34864
rect 8275 -34896 34275 -34890
rect 8275 -35204 8281 -34896
rect 8589 -34928 8961 -34896
rect 8589 -35172 8653 -34928
rect 8897 -35172 8961 -34928
rect 8589 -35204 8961 -35172
rect 9589 -34928 9961 -34896
rect 9589 -35172 9653 -34928
rect 9897 -35172 9961 -34928
rect 9589 -35204 9961 -35172
rect 10589 -34928 10961 -34896
rect 10589 -35172 10653 -34928
rect 10897 -35172 10961 -34928
rect 10589 -35204 10961 -35172
rect 11589 -34928 11961 -34896
rect 11589 -35172 11653 -34928
rect 11897 -35172 11961 -34928
rect 11589 -35204 11961 -35172
rect 12589 -34928 12961 -34896
rect 12589 -35172 12653 -34928
rect 12897 -35172 12961 -34928
rect 12589 -35204 12961 -35172
rect 13589 -34928 13961 -34896
rect 13589 -35172 13653 -34928
rect 13897 -35172 13961 -34928
rect 13589 -35204 13961 -35172
rect 14589 -34928 14961 -34896
rect 14589 -35172 14653 -34928
rect 14897 -35172 14961 -34928
rect 14589 -35204 14961 -35172
rect 15589 -34928 15961 -34896
rect 15589 -35172 15653 -34928
rect 15897 -35172 15961 -34928
rect 15589 -35204 15961 -35172
rect 16589 -34928 16961 -34896
rect 16589 -35172 16653 -34928
rect 16897 -35172 16961 -34928
rect 16589 -35204 16961 -35172
rect 17589 -34928 17961 -34896
rect 17589 -35172 17653 -34928
rect 17897 -35172 17961 -34928
rect 17589 -35204 17961 -35172
rect 18589 -34928 18961 -34896
rect 18589 -35172 18653 -34928
rect 18897 -35172 18961 -34928
rect 18589 -35204 18961 -35172
rect 19589 -34928 19961 -34896
rect 19589 -35172 19653 -34928
rect 19897 -35172 19961 -34928
rect 19589 -35204 19961 -35172
rect 20589 -34928 20961 -34896
rect 20589 -35172 20653 -34928
rect 20897 -35172 20961 -34928
rect 20589 -35204 20961 -35172
rect 21589 -34928 21961 -34896
rect 21589 -35172 21653 -34928
rect 21897 -35172 21961 -34928
rect 21589 -35204 21961 -35172
rect 22589 -34928 22961 -34896
rect 22589 -35172 22653 -34928
rect 22897 -35172 22961 -34928
rect 22589 -35204 22961 -35172
rect 23589 -34928 23961 -34896
rect 23589 -35172 23653 -34928
rect 23897 -35172 23961 -34928
rect 23589 -35204 23961 -35172
rect 24589 -34928 24961 -34896
rect 24589 -35172 24653 -34928
rect 24897 -35172 24961 -34928
rect 24589 -35204 24961 -35172
rect 25589 -34928 25961 -34896
rect 25589 -35172 25653 -34928
rect 25897 -35172 25961 -34928
rect 25589 -35204 25961 -35172
rect 26589 -34928 26961 -34896
rect 26589 -35172 26653 -34928
rect 26897 -35172 26961 -34928
rect 26589 -35204 26961 -35172
rect 27589 -34928 27961 -34896
rect 27589 -35172 27653 -34928
rect 27897 -35172 27961 -34928
rect 27589 -35204 27961 -35172
rect 28589 -34928 28961 -34896
rect 28589 -35172 28653 -34928
rect 28897 -35172 28961 -34928
rect 28589 -35204 28961 -35172
rect 29589 -34928 29961 -34896
rect 29589 -35172 29653 -34928
rect 29897 -35172 29961 -34928
rect 29589 -35204 29961 -35172
rect 30589 -34928 30961 -34896
rect 30589 -35172 30653 -34928
rect 30897 -35172 30961 -34928
rect 30589 -35204 30961 -35172
rect 31589 -34928 31961 -34896
rect 31589 -35172 31653 -34928
rect 31897 -35172 31961 -34928
rect 31589 -35204 31961 -35172
rect 32589 -34928 32961 -34896
rect 32589 -35172 32653 -34928
rect 32897 -35172 32961 -34928
rect 32589 -35204 32961 -35172
rect 33589 -34928 33961 -34896
rect 33589 -35172 33653 -34928
rect 33897 -35172 33961 -34928
rect 33589 -35204 33961 -35172
rect 34269 -35204 34275 -34896
rect 8275 -35210 34275 -35204
rect 8615 -35236 8935 -35210
rect 8615 -35864 8621 -35236
rect 8929 -35864 8935 -35236
rect 8615 -35890 8935 -35864
rect 9615 -35236 9935 -35210
rect 9615 -35864 9621 -35236
rect 9929 -35864 9935 -35236
rect 9615 -35890 9935 -35864
rect 10615 -35236 10935 -35210
rect 10615 -35864 10621 -35236
rect 10929 -35864 10935 -35236
rect 10615 -35890 10935 -35864
rect 11615 -35236 11935 -35210
rect 11615 -35864 11621 -35236
rect 11929 -35864 11935 -35236
rect 11615 -35890 11935 -35864
rect 12615 -35236 12935 -35210
rect 12615 -35864 12621 -35236
rect 12929 -35864 12935 -35236
rect 12615 -35890 12935 -35864
rect 13615 -35236 13935 -35210
rect 13615 -35864 13621 -35236
rect 13929 -35864 13935 -35236
rect 13615 -35890 13935 -35864
rect 14615 -35236 14935 -35210
rect 14615 -35864 14621 -35236
rect 14929 -35864 14935 -35236
rect 14615 -35890 14935 -35864
rect 15615 -35236 15935 -35210
rect 15615 -35864 15621 -35236
rect 15929 -35864 15935 -35236
rect 15615 -35890 15935 -35864
rect 16615 -35236 16935 -35210
rect 16615 -35864 16621 -35236
rect 16929 -35864 16935 -35236
rect 16615 -35890 16935 -35864
rect 17615 -35236 17935 -35210
rect 17615 -35864 17621 -35236
rect 17929 -35864 17935 -35236
rect 17615 -35890 17935 -35864
rect 18615 -35236 18935 -35210
rect 18615 -35864 18621 -35236
rect 18929 -35864 18935 -35236
rect 18615 -35890 18935 -35864
rect 19615 -35236 19935 -35210
rect 19615 -35864 19621 -35236
rect 19929 -35864 19935 -35236
rect 19615 -35890 19935 -35864
rect 20615 -35236 20935 -35210
rect 20615 -35864 20621 -35236
rect 20929 -35864 20935 -35236
rect 20615 -35890 20935 -35864
rect 21615 -35236 21935 -35210
rect 21615 -35864 21621 -35236
rect 21929 -35864 21935 -35236
rect 21615 -35890 21935 -35864
rect 22615 -35236 22935 -35210
rect 22615 -35864 22621 -35236
rect 22929 -35864 22935 -35236
rect 22615 -35890 22935 -35864
rect 23615 -35236 23935 -35210
rect 23615 -35864 23621 -35236
rect 23929 -35864 23935 -35236
rect 23615 -35890 23935 -35864
rect 24615 -35236 24935 -35210
rect 24615 -35864 24621 -35236
rect 24929 -35864 24935 -35236
rect 24615 -35890 24935 -35864
rect 25615 -35236 25935 -35210
rect 25615 -35864 25621 -35236
rect 25929 -35864 25935 -35236
rect 25615 -35890 25935 -35864
rect 26615 -35236 26935 -35210
rect 26615 -35864 26621 -35236
rect 26929 -35864 26935 -35236
rect 26615 -35890 26935 -35864
rect 27615 -35236 27935 -35210
rect 27615 -35864 27621 -35236
rect 27929 -35864 27935 -35236
rect 27615 -35890 27935 -35864
rect 28615 -35236 28935 -35210
rect 28615 -35864 28621 -35236
rect 28929 -35864 28935 -35236
rect 28615 -35890 28935 -35864
rect 29615 -35236 29935 -35210
rect 29615 -35864 29621 -35236
rect 29929 -35864 29935 -35236
rect 29615 -35890 29935 -35864
rect 30615 -35236 30935 -35210
rect 30615 -35864 30621 -35236
rect 30929 -35864 30935 -35236
rect 30615 -35890 30935 -35864
rect 31615 -35236 31935 -35210
rect 31615 -35864 31621 -35236
rect 31929 -35864 31935 -35236
rect 31615 -35890 31935 -35864
rect 32615 -35236 32935 -35210
rect 32615 -35864 32621 -35236
rect 32929 -35864 32935 -35236
rect 32615 -35890 32935 -35864
rect 33615 -35236 33935 -35210
rect 33615 -35864 33621 -35236
rect 33929 -35864 33935 -35236
rect 33615 -35890 33935 -35864
rect 8275 -35896 34275 -35890
rect 8275 -36204 8281 -35896
rect 8589 -35928 8961 -35896
rect 8589 -36172 8653 -35928
rect 8897 -36172 8961 -35928
rect 8589 -36204 8961 -36172
rect 9589 -35928 9961 -35896
rect 9589 -36172 9653 -35928
rect 9897 -36172 9961 -35928
rect 9589 -36204 9961 -36172
rect 10589 -35928 10961 -35896
rect 10589 -36172 10653 -35928
rect 10897 -36172 10961 -35928
rect 10589 -36204 10961 -36172
rect 11589 -35928 11961 -35896
rect 11589 -36172 11653 -35928
rect 11897 -36172 11961 -35928
rect 11589 -36204 11961 -36172
rect 12589 -35928 12961 -35896
rect 12589 -36172 12653 -35928
rect 12897 -36172 12961 -35928
rect 12589 -36204 12961 -36172
rect 13589 -35928 13961 -35896
rect 13589 -36172 13653 -35928
rect 13897 -36172 13961 -35928
rect 13589 -36204 13961 -36172
rect 14589 -35928 14961 -35896
rect 14589 -36172 14653 -35928
rect 14897 -36172 14961 -35928
rect 14589 -36204 14961 -36172
rect 15589 -35928 15961 -35896
rect 15589 -36172 15653 -35928
rect 15897 -36172 15961 -35928
rect 15589 -36204 15961 -36172
rect 16589 -35928 16961 -35896
rect 16589 -36172 16653 -35928
rect 16897 -36172 16961 -35928
rect 16589 -36204 16961 -36172
rect 17589 -35928 17961 -35896
rect 17589 -36172 17653 -35928
rect 17897 -36172 17961 -35928
rect 17589 -36204 17961 -36172
rect 18589 -35928 18961 -35896
rect 18589 -36172 18653 -35928
rect 18897 -36172 18961 -35928
rect 18589 -36204 18961 -36172
rect 19589 -35928 19961 -35896
rect 19589 -36172 19653 -35928
rect 19897 -36172 19961 -35928
rect 19589 -36204 19961 -36172
rect 20589 -35928 20961 -35896
rect 20589 -36172 20653 -35928
rect 20897 -36172 20961 -35928
rect 20589 -36204 20961 -36172
rect 21589 -35928 21961 -35896
rect 21589 -36172 21653 -35928
rect 21897 -36172 21961 -35928
rect 21589 -36204 21961 -36172
rect 22589 -35928 22961 -35896
rect 22589 -36172 22653 -35928
rect 22897 -36172 22961 -35928
rect 22589 -36204 22961 -36172
rect 23589 -35928 23961 -35896
rect 23589 -36172 23653 -35928
rect 23897 -36172 23961 -35928
rect 23589 -36204 23961 -36172
rect 24589 -35928 24961 -35896
rect 24589 -36172 24653 -35928
rect 24897 -36172 24961 -35928
rect 24589 -36204 24961 -36172
rect 25589 -35928 25961 -35896
rect 25589 -36172 25653 -35928
rect 25897 -36172 25961 -35928
rect 25589 -36204 25961 -36172
rect 26589 -35928 26961 -35896
rect 26589 -36172 26653 -35928
rect 26897 -36172 26961 -35928
rect 26589 -36204 26961 -36172
rect 27589 -35928 27961 -35896
rect 27589 -36172 27653 -35928
rect 27897 -36172 27961 -35928
rect 27589 -36204 27961 -36172
rect 28589 -35928 28961 -35896
rect 28589 -36172 28653 -35928
rect 28897 -36172 28961 -35928
rect 28589 -36204 28961 -36172
rect 29589 -35928 29961 -35896
rect 29589 -36172 29653 -35928
rect 29897 -36172 29961 -35928
rect 29589 -36204 29961 -36172
rect 30589 -35928 30961 -35896
rect 30589 -36172 30653 -35928
rect 30897 -36172 30961 -35928
rect 30589 -36204 30961 -36172
rect 31589 -35928 31961 -35896
rect 31589 -36172 31653 -35928
rect 31897 -36172 31961 -35928
rect 31589 -36204 31961 -36172
rect 32589 -35928 32961 -35896
rect 32589 -36172 32653 -35928
rect 32897 -36172 32961 -35928
rect 32589 -36204 32961 -36172
rect 33589 -35928 33961 -35896
rect 33589 -36172 33653 -35928
rect 33897 -36172 33961 -35928
rect 33589 -36204 33961 -36172
rect 34269 -36204 34275 -35896
rect 8275 -36210 34275 -36204
rect 8615 -36236 8935 -36210
rect 8615 -36864 8621 -36236
rect 8929 -36864 8935 -36236
rect 8615 -36890 8935 -36864
rect 9615 -36236 9935 -36210
rect 9615 -36864 9621 -36236
rect 9929 -36864 9935 -36236
rect 9615 -36890 9935 -36864
rect 10615 -36236 10935 -36210
rect 10615 -36864 10621 -36236
rect 10929 -36864 10935 -36236
rect 10615 -36890 10935 -36864
rect 11615 -36236 11935 -36210
rect 11615 -36864 11621 -36236
rect 11929 -36864 11935 -36236
rect 11615 -36890 11935 -36864
rect 12615 -36236 12935 -36210
rect 12615 -36864 12621 -36236
rect 12929 -36864 12935 -36236
rect 12615 -36890 12935 -36864
rect 13615 -36236 13935 -36210
rect 13615 -36864 13621 -36236
rect 13929 -36864 13935 -36236
rect 13615 -36890 13935 -36864
rect 14615 -36236 14935 -36210
rect 14615 -36864 14621 -36236
rect 14929 -36864 14935 -36236
rect 14615 -36890 14935 -36864
rect 15615 -36236 15935 -36210
rect 15615 -36864 15621 -36236
rect 15929 -36864 15935 -36236
rect 15615 -36890 15935 -36864
rect 16615 -36236 16935 -36210
rect 16615 -36864 16621 -36236
rect 16929 -36864 16935 -36236
rect 16615 -36890 16935 -36864
rect 17615 -36236 17935 -36210
rect 17615 -36864 17621 -36236
rect 17929 -36864 17935 -36236
rect 17615 -36890 17935 -36864
rect 18615 -36236 18935 -36210
rect 18615 -36864 18621 -36236
rect 18929 -36864 18935 -36236
rect 18615 -36890 18935 -36864
rect 19615 -36236 19935 -36210
rect 19615 -36864 19621 -36236
rect 19929 -36864 19935 -36236
rect 19615 -36890 19935 -36864
rect 20615 -36236 20935 -36210
rect 20615 -36864 20621 -36236
rect 20929 -36864 20935 -36236
rect 20615 -36890 20935 -36864
rect 21615 -36236 21935 -36210
rect 21615 -36864 21621 -36236
rect 21929 -36864 21935 -36236
rect 21615 -36890 21935 -36864
rect 22615 -36236 22935 -36210
rect 22615 -36864 22621 -36236
rect 22929 -36864 22935 -36236
rect 22615 -36890 22935 -36864
rect 23615 -36236 23935 -36210
rect 23615 -36864 23621 -36236
rect 23929 -36864 23935 -36236
rect 23615 -36890 23935 -36864
rect 24615 -36236 24935 -36210
rect 24615 -36864 24621 -36236
rect 24929 -36864 24935 -36236
rect 24615 -36890 24935 -36864
rect 25615 -36236 25935 -36210
rect 25615 -36864 25621 -36236
rect 25929 -36864 25935 -36236
rect 25615 -36890 25935 -36864
rect 26615 -36236 26935 -36210
rect 26615 -36864 26621 -36236
rect 26929 -36864 26935 -36236
rect 26615 -36890 26935 -36864
rect 27615 -36236 27935 -36210
rect 27615 -36864 27621 -36236
rect 27929 -36864 27935 -36236
rect 27615 -36890 27935 -36864
rect 28615 -36236 28935 -36210
rect 28615 -36864 28621 -36236
rect 28929 -36864 28935 -36236
rect 28615 -36890 28935 -36864
rect 29615 -36236 29935 -36210
rect 29615 -36864 29621 -36236
rect 29929 -36864 29935 -36236
rect 29615 -36890 29935 -36864
rect 30615 -36236 30935 -36210
rect 30615 -36864 30621 -36236
rect 30929 -36864 30935 -36236
rect 30615 -36890 30935 -36864
rect 31615 -36236 31935 -36210
rect 31615 -36864 31621 -36236
rect 31929 -36864 31935 -36236
rect 31615 -36890 31935 -36864
rect 32615 -36236 32935 -36210
rect 32615 -36864 32621 -36236
rect 32929 -36864 32935 -36236
rect 32615 -36890 32935 -36864
rect 33615 -36236 33935 -36210
rect 33615 -36864 33621 -36236
rect 33929 -36864 33935 -36236
rect 33615 -36890 33935 -36864
rect 8275 -36896 34275 -36890
rect 8275 -37204 8281 -36896
rect 8589 -36928 8961 -36896
rect 8589 -37172 8653 -36928
rect 8897 -37172 8961 -36928
rect 8589 -37204 8961 -37172
rect 9589 -36928 9961 -36896
rect 9589 -37172 9653 -36928
rect 9897 -37172 9961 -36928
rect 9589 -37204 9961 -37172
rect 10589 -36928 10961 -36896
rect 10589 -37172 10653 -36928
rect 10897 -37172 10961 -36928
rect 10589 -37204 10961 -37172
rect 11589 -36928 11961 -36896
rect 11589 -37172 11653 -36928
rect 11897 -37172 11961 -36928
rect 11589 -37204 11961 -37172
rect 12589 -36928 12961 -36896
rect 12589 -37172 12653 -36928
rect 12897 -37172 12961 -36928
rect 12589 -37204 12961 -37172
rect 13589 -36928 13961 -36896
rect 13589 -37172 13653 -36928
rect 13897 -37172 13961 -36928
rect 13589 -37204 13961 -37172
rect 14589 -36928 14961 -36896
rect 14589 -37172 14653 -36928
rect 14897 -37172 14961 -36928
rect 14589 -37204 14961 -37172
rect 15589 -36928 15961 -36896
rect 15589 -37172 15653 -36928
rect 15897 -37172 15961 -36928
rect 15589 -37204 15961 -37172
rect 16589 -36928 16961 -36896
rect 16589 -37172 16653 -36928
rect 16897 -37172 16961 -36928
rect 16589 -37204 16961 -37172
rect 17589 -36928 17961 -36896
rect 17589 -37172 17653 -36928
rect 17897 -37172 17961 -36928
rect 17589 -37204 17961 -37172
rect 18589 -36928 18961 -36896
rect 18589 -37172 18653 -36928
rect 18897 -37172 18961 -36928
rect 18589 -37204 18961 -37172
rect 19589 -36928 19961 -36896
rect 19589 -37172 19653 -36928
rect 19897 -37172 19961 -36928
rect 19589 -37204 19961 -37172
rect 20589 -36928 20961 -36896
rect 20589 -37172 20653 -36928
rect 20897 -37172 20961 -36928
rect 20589 -37204 20961 -37172
rect 21589 -36928 21961 -36896
rect 21589 -37172 21653 -36928
rect 21897 -37172 21961 -36928
rect 21589 -37204 21961 -37172
rect 22589 -36928 22961 -36896
rect 22589 -37172 22653 -36928
rect 22897 -37172 22961 -36928
rect 22589 -37204 22961 -37172
rect 23589 -36928 23961 -36896
rect 23589 -37172 23653 -36928
rect 23897 -37172 23961 -36928
rect 23589 -37204 23961 -37172
rect 24589 -36928 24961 -36896
rect 24589 -37172 24653 -36928
rect 24897 -37172 24961 -36928
rect 24589 -37204 24961 -37172
rect 25589 -36928 25961 -36896
rect 25589 -37172 25653 -36928
rect 25897 -37172 25961 -36928
rect 25589 -37204 25961 -37172
rect 26589 -36928 26961 -36896
rect 26589 -37172 26653 -36928
rect 26897 -37172 26961 -36928
rect 26589 -37204 26961 -37172
rect 27589 -36928 27961 -36896
rect 27589 -37172 27653 -36928
rect 27897 -37172 27961 -36928
rect 27589 -37204 27961 -37172
rect 28589 -36928 28961 -36896
rect 28589 -37172 28653 -36928
rect 28897 -37172 28961 -36928
rect 28589 -37204 28961 -37172
rect 29589 -36928 29961 -36896
rect 29589 -37172 29653 -36928
rect 29897 -37172 29961 -36928
rect 29589 -37204 29961 -37172
rect 30589 -36928 30961 -36896
rect 30589 -37172 30653 -36928
rect 30897 -37172 30961 -36928
rect 30589 -37204 30961 -37172
rect 31589 -36928 31961 -36896
rect 31589 -37172 31653 -36928
rect 31897 -37172 31961 -36928
rect 31589 -37204 31961 -37172
rect 32589 -36928 32961 -36896
rect 32589 -37172 32653 -36928
rect 32897 -37172 32961 -36928
rect 32589 -37204 32961 -37172
rect 33589 -36928 33961 -36896
rect 33589 -37172 33653 -36928
rect 33897 -37172 33961 -36928
rect 33589 -37204 33961 -37172
rect 34269 -37204 34275 -36896
rect 8275 -37210 34275 -37204
rect 8615 -37236 8935 -37210
rect 8615 -37864 8621 -37236
rect 8929 -37864 8935 -37236
rect 8615 -37890 8935 -37864
rect 9615 -37236 9935 -37210
rect 9615 -37864 9621 -37236
rect 9929 -37864 9935 -37236
rect 9615 -37890 9935 -37864
rect 10615 -37236 10935 -37210
rect 10615 -37864 10621 -37236
rect 10929 -37864 10935 -37236
rect 10615 -37890 10935 -37864
rect 11615 -37236 11935 -37210
rect 11615 -37864 11621 -37236
rect 11929 -37864 11935 -37236
rect 11615 -37890 11935 -37864
rect 12615 -37236 12935 -37210
rect 12615 -37864 12621 -37236
rect 12929 -37864 12935 -37236
rect 12615 -37890 12935 -37864
rect 13615 -37236 13935 -37210
rect 13615 -37864 13621 -37236
rect 13929 -37864 13935 -37236
rect 13615 -37890 13935 -37864
rect 14615 -37236 14935 -37210
rect 14615 -37864 14621 -37236
rect 14929 -37864 14935 -37236
rect 14615 -37890 14935 -37864
rect 15615 -37236 15935 -37210
rect 15615 -37864 15621 -37236
rect 15929 -37864 15935 -37236
rect 15615 -37890 15935 -37864
rect 16615 -37236 16935 -37210
rect 16615 -37864 16621 -37236
rect 16929 -37864 16935 -37236
rect 16615 -37890 16935 -37864
rect 17615 -37236 17935 -37210
rect 17615 -37864 17621 -37236
rect 17929 -37864 17935 -37236
rect 17615 -37890 17935 -37864
rect 18615 -37236 18935 -37210
rect 18615 -37864 18621 -37236
rect 18929 -37864 18935 -37236
rect 18615 -37890 18935 -37864
rect 19615 -37236 19935 -37210
rect 19615 -37864 19621 -37236
rect 19929 -37864 19935 -37236
rect 19615 -37890 19935 -37864
rect 20615 -37236 20935 -37210
rect 20615 -37864 20621 -37236
rect 20929 -37864 20935 -37236
rect 20615 -37890 20935 -37864
rect 21615 -37236 21935 -37210
rect 21615 -37864 21621 -37236
rect 21929 -37864 21935 -37236
rect 21615 -37890 21935 -37864
rect 22615 -37236 22935 -37210
rect 22615 -37864 22621 -37236
rect 22929 -37864 22935 -37236
rect 22615 -37890 22935 -37864
rect 23615 -37236 23935 -37210
rect 23615 -37864 23621 -37236
rect 23929 -37864 23935 -37236
rect 23615 -37890 23935 -37864
rect 24615 -37236 24935 -37210
rect 24615 -37864 24621 -37236
rect 24929 -37864 24935 -37236
rect 24615 -37890 24935 -37864
rect 25615 -37236 25935 -37210
rect 25615 -37864 25621 -37236
rect 25929 -37864 25935 -37236
rect 25615 -37890 25935 -37864
rect 26615 -37236 26935 -37210
rect 26615 -37864 26621 -37236
rect 26929 -37864 26935 -37236
rect 26615 -37890 26935 -37864
rect 27615 -37236 27935 -37210
rect 27615 -37864 27621 -37236
rect 27929 -37864 27935 -37236
rect 27615 -37890 27935 -37864
rect 28615 -37236 28935 -37210
rect 28615 -37864 28621 -37236
rect 28929 -37864 28935 -37236
rect 28615 -37890 28935 -37864
rect 29615 -37236 29935 -37210
rect 29615 -37864 29621 -37236
rect 29929 -37864 29935 -37236
rect 29615 -37890 29935 -37864
rect 30615 -37236 30935 -37210
rect 30615 -37864 30621 -37236
rect 30929 -37864 30935 -37236
rect 30615 -37890 30935 -37864
rect 31615 -37236 31935 -37210
rect 31615 -37864 31621 -37236
rect 31929 -37864 31935 -37236
rect 31615 -37890 31935 -37864
rect 32615 -37236 32935 -37210
rect 32615 -37864 32621 -37236
rect 32929 -37864 32935 -37236
rect 32615 -37890 32935 -37864
rect 33615 -37236 33935 -37210
rect 33615 -37864 33621 -37236
rect 33929 -37864 33935 -37236
rect 33615 -37890 33935 -37864
rect 8275 -37896 34275 -37890
rect 8275 -38204 8281 -37896
rect 8589 -37928 8961 -37896
rect 8589 -38172 8653 -37928
rect 8897 -38172 8961 -37928
rect 8589 -38204 8961 -38172
rect 9589 -37928 9961 -37896
rect 9589 -38172 9653 -37928
rect 9897 -38172 9961 -37928
rect 9589 -38204 9961 -38172
rect 10589 -37928 10961 -37896
rect 10589 -38172 10653 -37928
rect 10897 -38172 10961 -37928
rect 10589 -38204 10961 -38172
rect 11589 -37928 11961 -37896
rect 11589 -38172 11653 -37928
rect 11897 -38172 11961 -37928
rect 11589 -38204 11961 -38172
rect 12589 -37928 12961 -37896
rect 12589 -38172 12653 -37928
rect 12897 -38172 12961 -37928
rect 12589 -38204 12961 -38172
rect 13589 -37928 13961 -37896
rect 13589 -38172 13653 -37928
rect 13897 -38172 13961 -37928
rect 13589 -38204 13961 -38172
rect 14589 -37928 14961 -37896
rect 14589 -38172 14653 -37928
rect 14897 -38172 14961 -37928
rect 14589 -38204 14961 -38172
rect 15589 -37928 15961 -37896
rect 15589 -38172 15653 -37928
rect 15897 -38172 15961 -37928
rect 15589 -38204 15961 -38172
rect 16589 -37928 16961 -37896
rect 16589 -38172 16653 -37928
rect 16897 -38172 16961 -37928
rect 16589 -38204 16961 -38172
rect 17589 -37928 17961 -37896
rect 17589 -38172 17653 -37928
rect 17897 -38172 17961 -37928
rect 17589 -38204 17961 -38172
rect 18589 -37928 18961 -37896
rect 18589 -38172 18653 -37928
rect 18897 -38172 18961 -37928
rect 18589 -38204 18961 -38172
rect 19589 -37928 19961 -37896
rect 19589 -38172 19653 -37928
rect 19897 -38172 19961 -37928
rect 19589 -38204 19961 -38172
rect 20589 -37928 20961 -37896
rect 20589 -38172 20653 -37928
rect 20897 -38172 20961 -37928
rect 20589 -38204 20961 -38172
rect 21589 -37928 21961 -37896
rect 21589 -38172 21653 -37928
rect 21897 -38172 21961 -37928
rect 21589 -38204 21961 -38172
rect 22589 -37928 22961 -37896
rect 22589 -38172 22653 -37928
rect 22897 -38172 22961 -37928
rect 22589 -38204 22961 -38172
rect 23589 -37928 23961 -37896
rect 23589 -38172 23653 -37928
rect 23897 -38172 23961 -37928
rect 23589 -38204 23961 -38172
rect 24589 -37928 24961 -37896
rect 24589 -38172 24653 -37928
rect 24897 -38172 24961 -37928
rect 24589 -38204 24961 -38172
rect 25589 -37928 25961 -37896
rect 25589 -38172 25653 -37928
rect 25897 -38172 25961 -37928
rect 25589 -38204 25961 -38172
rect 26589 -37928 26961 -37896
rect 26589 -38172 26653 -37928
rect 26897 -38172 26961 -37928
rect 26589 -38204 26961 -38172
rect 27589 -37928 27961 -37896
rect 27589 -38172 27653 -37928
rect 27897 -38172 27961 -37928
rect 27589 -38204 27961 -38172
rect 28589 -37928 28961 -37896
rect 28589 -38172 28653 -37928
rect 28897 -38172 28961 -37928
rect 28589 -38204 28961 -38172
rect 29589 -37928 29961 -37896
rect 29589 -38172 29653 -37928
rect 29897 -38172 29961 -37928
rect 29589 -38204 29961 -38172
rect 30589 -37928 30961 -37896
rect 30589 -38172 30653 -37928
rect 30897 -38172 30961 -37928
rect 30589 -38204 30961 -38172
rect 31589 -37928 31961 -37896
rect 31589 -38172 31653 -37928
rect 31897 -38172 31961 -37928
rect 31589 -38204 31961 -38172
rect 32589 -37928 32961 -37896
rect 32589 -38172 32653 -37928
rect 32897 -38172 32961 -37928
rect 32589 -38204 32961 -38172
rect 33589 -37928 33961 -37896
rect 33589 -38172 33653 -37928
rect 33897 -38172 33961 -37928
rect 33589 -38204 33961 -38172
rect 34269 -38204 34275 -37896
rect 8275 -38210 34275 -38204
rect 8615 -38236 8935 -38210
rect 8615 -38864 8621 -38236
rect 8929 -38864 8935 -38236
rect 8615 -38890 8935 -38864
rect 9615 -38236 9935 -38210
rect 9615 -38864 9621 -38236
rect 9929 -38864 9935 -38236
rect 9615 -38890 9935 -38864
rect 10615 -38236 10935 -38210
rect 10615 -38864 10621 -38236
rect 10929 -38864 10935 -38236
rect 10615 -38890 10935 -38864
rect 11615 -38236 11935 -38210
rect 11615 -38864 11621 -38236
rect 11929 -38864 11935 -38236
rect 11615 -38890 11935 -38864
rect 12615 -38236 12935 -38210
rect 12615 -38864 12621 -38236
rect 12929 -38864 12935 -38236
rect 12615 -38890 12935 -38864
rect 13615 -38236 13935 -38210
rect 13615 -38864 13621 -38236
rect 13929 -38864 13935 -38236
rect 13615 -38890 13935 -38864
rect 14615 -38236 14935 -38210
rect 14615 -38864 14621 -38236
rect 14929 -38864 14935 -38236
rect 14615 -38890 14935 -38864
rect 15615 -38236 15935 -38210
rect 15615 -38864 15621 -38236
rect 15929 -38864 15935 -38236
rect 15615 -38890 15935 -38864
rect 16615 -38236 16935 -38210
rect 16615 -38864 16621 -38236
rect 16929 -38864 16935 -38236
rect 16615 -38890 16935 -38864
rect 17615 -38236 17935 -38210
rect 17615 -38864 17621 -38236
rect 17929 -38864 17935 -38236
rect 17615 -38890 17935 -38864
rect 18615 -38236 18935 -38210
rect 18615 -38864 18621 -38236
rect 18929 -38864 18935 -38236
rect 18615 -38890 18935 -38864
rect 19615 -38236 19935 -38210
rect 19615 -38864 19621 -38236
rect 19929 -38864 19935 -38236
rect 19615 -38890 19935 -38864
rect 20615 -38236 20935 -38210
rect 20615 -38864 20621 -38236
rect 20929 -38864 20935 -38236
rect 20615 -38890 20935 -38864
rect 21615 -38236 21935 -38210
rect 21615 -38864 21621 -38236
rect 21929 -38864 21935 -38236
rect 21615 -38890 21935 -38864
rect 22615 -38236 22935 -38210
rect 22615 -38864 22621 -38236
rect 22929 -38864 22935 -38236
rect 22615 -38890 22935 -38864
rect 23615 -38236 23935 -38210
rect 23615 -38864 23621 -38236
rect 23929 -38864 23935 -38236
rect 23615 -38890 23935 -38864
rect 24615 -38236 24935 -38210
rect 24615 -38864 24621 -38236
rect 24929 -38864 24935 -38236
rect 24615 -38890 24935 -38864
rect 25615 -38236 25935 -38210
rect 25615 -38864 25621 -38236
rect 25929 -38864 25935 -38236
rect 25615 -38890 25935 -38864
rect 26615 -38236 26935 -38210
rect 26615 -38864 26621 -38236
rect 26929 -38864 26935 -38236
rect 26615 -38890 26935 -38864
rect 27615 -38236 27935 -38210
rect 27615 -38864 27621 -38236
rect 27929 -38864 27935 -38236
rect 27615 -38890 27935 -38864
rect 28615 -38236 28935 -38210
rect 28615 -38864 28621 -38236
rect 28929 -38864 28935 -38236
rect 28615 -38890 28935 -38864
rect 29615 -38236 29935 -38210
rect 29615 -38864 29621 -38236
rect 29929 -38864 29935 -38236
rect 29615 -38890 29935 -38864
rect 30615 -38236 30935 -38210
rect 30615 -38864 30621 -38236
rect 30929 -38864 30935 -38236
rect 30615 -38890 30935 -38864
rect 31615 -38236 31935 -38210
rect 31615 -38864 31621 -38236
rect 31929 -38864 31935 -38236
rect 31615 -38890 31935 -38864
rect 32615 -38236 32935 -38210
rect 32615 -38864 32621 -38236
rect 32929 -38864 32935 -38236
rect 32615 -38890 32935 -38864
rect 33615 -38236 33935 -38210
rect 33615 -38864 33621 -38236
rect 33929 -38864 33935 -38236
rect 33615 -38890 33935 -38864
rect 8275 -38896 34275 -38890
rect 8275 -39204 8281 -38896
rect 8589 -38928 8961 -38896
rect 8589 -39172 8653 -38928
rect 8897 -39172 8961 -38928
rect 8589 -39204 8961 -39172
rect 9589 -38928 9961 -38896
rect 9589 -39172 9653 -38928
rect 9897 -39172 9961 -38928
rect 9589 -39204 9961 -39172
rect 10589 -38928 10961 -38896
rect 10589 -39172 10653 -38928
rect 10897 -39172 10961 -38928
rect 10589 -39204 10961 -39172
rect 11589 -38928 11961 -38896
rect 11589 -39172 11653 -38928
rect 11897 -39172 11961 -38928
rect 11589 -39204 11961 -39172
rect 12589 -38928 12961 -38896
rect 12589 -39172 12653 -38928
rect 12897 -39172 12961 -38928
rect 12589 -39204 12961 -39172
rect 13589 -38928 13961 -38896
rect 13589 -39172 13653 -38928
rect 13897 -39172 13961 -38928
rect 13589 -39204 13961 -39172
rect 14589 -38928 14961 -38896
rect 14589 -39172 14653 -38928
rect 14897 -39172 14961 -38928
rect 14589 -39204 14961 -39172
rect 15589 -38928 15961 -38896
rect 15589 -39172 15653 -38928
rect 15897 -39172 15961 -38928
rect 15589 -39204 15961 -39172
rect 16589 -38928 16961 -38896
rect 16589 -39172 16653 -38928
rect 16897 -39172 16961 -38928
rect 16589 -39204 16961 -39172
rect 17589 -38928 17961 -38896
rect 17589 -39172 17653 -38928
rect 17897 -39172 17961 -38928
rect 17589 -39204 17961 -39172
rect 18589 -38928 18961 -38896
rect 18589 -39172 18653 -38928
rect 18897 -39172 18961 -38928
rect 18589 -39204 18961 -39172
rect 19589 -38928 19961 -38896
rect 19589 -39172 19653 -38928
rect 19897 -39172 19961 -38928
rect 19589 -39204 19961 -39172
rect 20589 -38928 20961 -38896
rect 20589 -39172 20653 -38928
rect 20897 -39172 20961 -38928
rect 20589 -39204 20961 -39172
rect 21589 -38928 21961 -38896
rect 21589 -39172 21653 -38928
rect 21897 -39172 21961 -38928
rect 21589 -39204 21961 -39172
rect 22589 -38928 22961 -38896
rect 22589 -39172 22653 -38928
rect 22897 -39172 22961 -38928
rect 22589 -39204 22961 -39172
rect 23589 -38928 23961 -38896
rect 23589 -39172 23653 -38928
rect 23897 -39172 23961 -38928
rect 23589 -39204 23961 -39172
rect 24589 -38928 24961 -38896
rect 24589 -39172 24653 -38928
rect 24897 -39172 24961 -38928
rect 24589 -39204 24961 -39172
rect 25589 -38928 25961 -38896
rect 25589 -39172 25653 -38928
rect 25897 -39172 25961 -38928
rect 25589 -39204 25961 -39172
rect 26589 -38928 26961 -38896
rect 26589 -39172 26653 -38928
rect 26897 -39172 26961 -38928
rect 26589 -39204 26961 -39172
rect 27589 -38928 27961 -38896
rect 27589 -39172 27653 -38928
rect 27897 -39172 27961 -38928
rect 27589 -39204 27961 -39172
rect 28589 -38928 28961 -38896
rect 28589 -39172 28653 -38928
rect 28897 -39172 28961 -38928
rect 28589 -39204 28961 -39172
rect 29589 -38928 29961 -38896
rect 29589 -39172 29653 -38928
rect 29897 -39172 29961 -38928
rect 29589 -39204 29961 -39172
rect 30589 -38928 30961 -38896
rect 30589 -39172 30653 -38928
rect 30897 -39172 30961 -38928
rect 30589 -39204 30961 -39172
rect 31589 -38928 31961 -38896
rect 31589 -39172 31653 -38928
rect 31897 -39172 31961 -38928
rect 31589 -39204 31961 -39172
rect 32589 -38928 32961 -38896
rect 32589 -39172 32653 -38928
rect 32897 -39172 32961 -38928
rect 32589 -39204 32961 -39172
rect 33589 -38928 33961 -38896
rect 33589 -39172 33653 -38928
rect 33897 -39172 33961 -38928
rect 33589 -39204 33961 -39172
rect 34269 -39204 34275 -38896
rect 8275 -39210 34275 -39204
rect 8615 -39236 8935 -39210
rect 8615 -39864 8621 -39236
rect 8929 -39864 8935 -39236
rect 8615 -39890 8935 -39864
rect 9615 -39236 9935 -39210
rect 9615 -39864 9621 -39236
rect 9929 -39864 9935 -39236
rect 9615 -39890 9935 -39864
rect 10615 -39236 10935 -39210
rect 10615 -39864 10621 -39236
rect 10929 -39864 10935 -39236
rect 10615 -39890 10935 -39864
rect 11615 -39236 11935 -39210
rect 11615 -39864 11621 -39236
rect 11929 -39864 11935 -39236
rect 11615 -39890 11935 -39864
rect 12615 -39236 12935 -39210
rect 12615 -39864 12621 -39236
rect 12929 -39864 12935 -39236
rect 12615 -39890 12935 -39864
rect 13615 -39236 13935 -39210
rect 13615 -39864 13621 -39236
rect 13929 -39864 13935 -39236
rect 13615 -39890 13935 -39864
rect 14615 -39236 14935 -39210
rect 14615 -39864 14621 -39236
rect 14929 -39864 14935 -39236
rect 14615 -39890 14935 -39864
rect 15615 -39236 15935 -39210
rect 15615 -39864 15621 -39236
rect 15929 -39864 15935 -39236
rect 15615 -39890 15935 -39864
rect 16615 -39236 16935 -39210
rect 16615 -39864 16621 -39236
rect 16929 -39864 16935 -39236
rect 16615 -39890 16935 -39864
rect 17615 -39236 17935 -39210
rect 17615 -39864 17621 -39236
rect 17929 -39864 17935 -39236
rect 17615 -39890 17935 -39864
rect 18615 -39236 18935 -39210
rect 18615 -39864 18621 -39236
rect 18929 -39864 18935 -39236
rect 18615 -39890 18935 -39864
rect 19615 -39236 19935 -39210
rect 19615 -39864 19621 -39236
rect 19929 -39864 19935 -39236
rect 19615 -39890 19935 -39864
rect 20615 -39236 20935 -39210
rect 20615 -39864 20621 -39236
rect 20929 -39864 20935 -39236
rect 20615 -39890 20935 -39864
rect 21615 -39236 21935 -39210
rect 21615 -39864 21621 -39236
rect 21929 -39864 21935 -39236
rect 21615 -39890 21935 -39864
rect 22615 -39236 22935 -39210
rect 22615 -39864 22621 -39236
rect 22929 -39864 22935 -39236
rect 22615 -39890 22935 -39864
rect 23615 -39236 23935 -39210
rect 23615 -39864 23621 -39236
rect 23929 -39864 23935 -39236
rect 23615 -39890 23935 -39864
rect 24615 -39236 24935 -39210
rect 24615 -39864 24621 -39236
rect 24929 -39864 24935 -39236
rect 24615 -39890 24935 -39864
rect 25615 -39236 25935 -39210
rect 25615 -39864 25621 -39236
rect 25929 -39864 25935 -39236
rect 25615 -39890 25935 -39864
rect 26615 -39236 26935 -39210
rect 26615 -39864 26621 -39236
rect 26929 -39864 26935 -39236
rect 26615 -39890 26935 -39864
rect 27615 -39236 27935 -39210
rect 27615 -39864 27621 -39236
rect 27929 -39864 27935 -39236
rect 27615 -39890 27935 -39864
rect 28615 -39236 28935 -39210
rect 28615 -39864 28621 -39236
rect 28929 -39864 28935 -39236
rect 28615 -39890 28935 -39864
rect 29615 -39236 29935 -39210
rect 29615 -39864 29621 -39236
rect 29929 -39864 29935 -39236
rect 29615 -39890 29935 -39864
rect 30615 -39236 30935 -39210
rect 30615 -39864 30621 -39236
rect 30929 -39864 30935 -39236
rect 30615 -39890 30935 -39864
rect 31615 -39236 31935 -39210
rect 31615 -39864 31621 -39236
rect 31929 -39864 31935 -39236
rect 31615 -39890 31935 -39864
rect 32615 -39236 32935 -39210
rect 32615 -39864 32621 -39236
rect 32929 -39864 32935 -39236
rect 32615 -39890 32935 -39864
rect 33615 -39236 33935 -39210
rect 33615 -39864 33621 -39236
rect 33929 -39864 33935 -39236
rect 33615 -39890 33935 -39864
rect 8275 -39896 34275 -39890
rect 8275 -40204 8281 -39896
rect 8589 -39928 8961 -39896
rect 8589 -40172 8653 -39928
rect 8897 -40172 8961 -39928
rect 8589 -40204 8961 -40172
rect 9589 -39928 9961 -39896
rect 9589 -40172 9653 -39928
rect 9897 -40172 9961 -39928
rect 9589 -40204 9961 -40172
rect 10589 -39928 10961 -39896
rect 10589 -40172 10653 -39928
rect 10897 -40172 10961 -39928
rect 10589 -40204 10961 -40172
rect 11589 -39928 11961 -39896
rect 11589 -40172 11653 -39928
rect 11897 -40172 11961 -39928
rect 11589 -40204 11961 -40172
rect 12589 -39928 12961 -39896
rect 12589 -40172 12653 -39928
rect 12897 -40172 12961 -39928
rect 12589 -40204 12961 -40172
rect 13589 -39928 13961 -39896
rect 13589 -40172 13653 -39928
rect 13897 -40172 13961 -39928
rect 13589 -40204 13961 -40172
rect 14589 -39928 14961 -39896
rect 14589 -40172 14653 -39928
rect 14897 -40172 14961 -39928
rect 14589 -40204 14961 -40172
rect 15589 -39928 15961 -39896
rect 15589 -40172 15653 -39928
rect 15897 -40172 15961 -39928
rect 15589 -40204 15961 -40172
rect 16589 -39928 16961 -39896
rect 16589 -40172 16653 -39928
rect 16897 -40172 16961 -39928
rect 16589 -40204 16961 -40172
rect 17589 -39928 17961 -39896
rect 17589 -40172 17653 -39928
rect 17897 -40172 17961 -39928
rect 17589 -40204 17961 -40172
rect 18589 -39928 18961 -39896
rect 18589 -40172 18653 -39928
rect 18897 -40172 18961 -39928
rect 18589 -40204 18961 -40172
rect 19589 -39928 19961 -39896
rect 19589 -40172 19653 -39928
rect 19897 -40172 19961 -39928
rect 19589 -40204 19961 -40172
rect 20589 -39928 20961 -39896
rect 20589 -40172 20653 -39928
rect 20897 -40172 20961 -39928
rect 20589 -40204 20961 -40172
rect 21589 -39928 21961 -39896
rect 21589 -40172 21653 -39928
rect 21897 -40172 21961 -39928
rect 21589 -40204 21961 -40172
rect 22589 -39928 22961 -39896
rect 22589 -40172 22653 -39928
rect 22897 -40172 22961 -39928
rect 22589 -40204 22961 -40172
rect 23589 -39928 23961 -39896
rect 23589 -40172 23653 -39928
rect 23897 -40172 23961 -39928
rect 23589 -40204 23961 -40172
rect 24589 -39928 24961 -39896
rect 24589 -40172 24653 -39928
rect 24897 -40172 24961 -39928
rect 24589 -40204 24961 -40172
rect 25589 -39928 25961 -39896
rect 25589 -40172 25653 -39928
rect 25897 -40172 25961 -39928
rect 25589 -40204 25961 -40172
rect 26589 -39928 26961 -39896
rect 26589 -40172 26653 -39928
rect 26897 -40172 26961 -39928
rect 26589 -40204 26961 -40172
rect 27589 -39928 27961 -39896
rect 27589 -40172 27653 -39928
rect 27897 -40172 27961 -39928
rect 27589 -40204 27961 -40172
rect 28589 -39928 28961 -39896
rect 28589 -40172 28653 -39928
rect 28897 -40172 28961 -39928
rect 28589 -40204 28961 -40172
rect 29589 -39928 29961 -39896
rect 29589 -40172 29653 -39928
rect 29897 -40172 29961 -39928
rect 29589 -40204 29961 -40172
rect 30589 -39928 30961 -39896
rect 30589 -40172 30653 -39928
rect 30897 -40172 30961 -39928
rect 30589 -40204 30961 -40172
rect 31589 -39928 31961 -39896
rect 31589 -40172 31653 -39928
rect 31897 -40172 31961 -39928
rect 31589 -40204 31961 -40172
rect 32589 -39928 32961 -39896
rect 32589 -40172 32653 -39928
rect 32897 -40172 32961 -39928
rect 32589 -40204 32961 -40172
rect 33589 -39928 33961 -39896
rect 33589 -40172 33653 -39928
rect 33897 -40172 33961 -39928
rect 33589 -40204 33961 -40172
rect 34269 -40204 34275 -39896
rect 8275 -40210 34275 -40204
rect 8615 -40236 8935 -40210
rect 8615 -40864 8621 -40236
rect 8929 -40864 8935 -40236
rect 8615 -40890 8935 -40864
rect 9615 -40236 9935 -40210
rect 9615 -40864 9621 -40236
rect 9929 -40864 9935 -40236
rect 9615 -40890 9935 -40864
rect 10615 -40236 10935 -40210
rect 10615 -40864 10621 -40236
rect 10929 -40864 10935 -40236
rect 10615 -40890 10935 -40864
rect 11615 -40236 11935 -40210
rect 11615 -40864 11621 -40236
rect 11929 -40864 11935 -40236
rect 11615 -40890 11935 -40864
rect 12615 -40236 12935 -40210
rect 12615 -40864 12621 -40236
rect 12929 -40864 12935 -40236
rect 12615 -40890 12935 -40864
rect 13615 -40236 13935 -40210
rect 13615 -40864 13621 -40236
rect 13929 -40864 13935 -40236
rect 13615 -40890 13935 -40864
rect 14615 -40236 14935 -40210
rect 14615 -40864 14621 -40236
rect 14929 -40864 14935 -40236
rect 14615 -40890 14935 -40864
rect 15615 -40236 15935 -40210
rect 15615 -40864 15621 -40236
rect 15929 -40864 15935 -40236
rect 15615 -40890 15935 -40864
rect 16615 -40236 16935 -40210
rect 16615 -40864 16621 -40236
rect 16929 -40864 16935 -40236
rect 16615 -40890 16935 -40864
rect 17615 -40236 17935 -40210
rect 17615 -40864 17621 -40236
rect 17929 -40864 17935 -40236
rect 17615 -40890 17935 -40864
rect 18615 -40236 18935 -40210
rect 18615 -40864 18621 -40236
rect 18929 -40864 18935 -40236
rect 18615 -40890 18935 -40864
rect 19615 -40236 19935 -40210
rect 19615 -40864 19621 -40236
rect 19929 -40864 19935 -40236
rect 19615 -40890 19935 -40864
rect 20615 -40236 20935 -40210
rect 20615 -40864 20621 -40236
rect 20929 -40864 20935 -40236
rect 20615 -40890 20935 -40864
rect 21615 -40236 21935 -40210
rect 21615 -40864 21621 -40236
rect 21929 -40864 21935 -40236
rect 21615 -40890 21935 -40864
rect 22615 -40236 22935 -40210
rect 22615 -40864 22621 -40236
rect 22929 -40864 22935 -40236
rect 22615 -40890 22935 -40864
rect 23615 -40236 23935 -40210
rect 23615 -40864 23621 -40236
rect 23929 -40864 23935 -40236
rect 23615 -40890 23935 -40864
rect 24615 -40236 24935 -40210
rect 24615 -40864 24621 -40236
rect 24929 -40864 24935 -40236
rect 24615 -40890 24935 -40864
rect 25615 -40236 25935 -40210
rect 25615 -40864 25621 -40236
rect 25929 -40864 25935 -40236
rect 25615 -40890 25935 -40864
rect 26615 -40236 26935 -40210
rect 26615 -40864 26621 -40236
rect 26929 -40864 26935 -40236
rect 26615 -40890 26935 -40864
rect 27615 -40236 27935 -40210
rect 27615 -40864 27621 -40236
rect 27929 -40864 27935 -40236
rect 27615 -40890 27935 -40864
rect 28615 -40236 28935 -40210
rect 28615 -40864 28621 -40236
rect 28929 -40864 28935 -40236
rect 28615 -40890 28935 -40864
rect 29615 -40236 29935 -40210
rect 29615 -40864 29621 -40236
rect 29929 -40864 29935 -40236
rect 29615 -40890 29935 -40864
rect 30615 -40236 30935 -40210
rect 30615 -40864 30621 -40236
rect 30929 -40864 30935 -40236
rect 30615 -40890 30935 -40864
rect 31615 -40236 31935 -40210
rect 31615 -40864 31621 -40236
rect 31929 -40864 31935 -40236
rect 31615 -40890 31935 -40864
rect 32615 -40236 32935 -40210
rect 32615 -40864 32621 -40236
rect 32929 -40864 32935 -40236
rect 32615 -40890 32935 -40864
rect 33615 -40236 33935 -40210
rect 33615 -40864 33621 -40236
rect 33929 -40864 33935 -40236
rect 33615 -40890 33935 -40864
rect 8275 -40896 34275 -40890
rect 8275 -41204 8281 -40896
rect 8589 -40928 8961 -40896
rect 8589 -41172 8653 -40928
rect 8897 -41172 8961 -40928
rect 8589 -41204 8961 -41172
rect 9589 -40928 9961 -40896
rect 9589 -41172 9653 -40928
rect 9897 -41172 9961 -40928
rect 9589 -41204 9961 -41172
rect 10589 -40928 10961 -40896
rect 10589 -41172 10653 -40928
rect 10897 -41172 10961 -40928
rect 10589 -41204 10961 -41172
rect 11589 -40928 11961 -40896
rect 11589 -41172 11653 -40928
rect 11897 -41172 11961 -40928
rect 11589 -41204 11961 -41172
rect 12589 -40928 12961 -40896
rect 12589 -41172 12653 -40928
rect 12897 -41172 12961 -40928
rect 12589 -41204 12961 -41172
rect 13589 -40928 13961 -40896
rect 13589 -41172 13653 -40928
rect 13897 -41172 13961 -40928
rect 13589 -41204 13961 -41172
rect 14589 -40928 14961 -40896
rect 14589 -41172 14653 -40928
rect 14897 -41172 14961 -40928
rect 14589 -41204 14961 -41172
rect 15589 -40928 15961 -40896
rect 15589 -41172 15653 -40928
rect 15897 -41172 15961 -40928
rect 15589 -41204 15961 -41172
rect 16589 -40928 16961 -40896
rect 16589 -41172 16653 -40928
rect 16897 -41172 16961 -40928
rect 16589 -41204 16961 -41172
rect 17589 -40928 17961 -40896
rect 17589 -41172 17653 -40928
rect 17897 -41172 17961 -40928
rect 17589 -41204 17961 -41172
rect 18589 -40928 18961 -40896
rect 18589 -41172 18653 -40928
rect 18897 -41172 18961 -40928
rect 18589 -41204 18961 -41172
rect 19589 -40928 19961 -40896
rect 19589 -41172 19653 -40928
rect 19897 -41172 19961 -40928
rect 19589 -41204 19961 -41172
rect 20589 -40928 20961 -40896
rect 20589 -41172 20653 -40928
rect 20897 -41172 20961 -40928
rect 20589 -41204 20961 -41172
rect 21589 -40928 21961 -40896
rect 21589 -41172 21653 -40928
rect 21897 -41172 21961 -40928
rect 21589 -41204 21961 -41172
rect 22589 -40928 22961 -40896
rect 22589 -41172 22653 -40928
rect 22897 -41172 22961 -40928
rect 22589 -41204 22961 -41172
rect 23589 -40928 23961 -40896
rect 23589 -41172 23653 -40928
rect 23897 -41172 23961 -40928
rect 23589 -41204 23961 -41172
rect 24589 -40928 24961 -40896
rect 24589 -41172 24653 -40928
rect 24897 -41172 24961 -40928
rect 24589 -41204 24961 -41172
rect 25589 -40928 25961 -40896
rect 25589 -41172 25653 -40928
rect 25897 -41172 25961 -40928
rect 25589 -41204 25961 -41172
rect 26589 -40928 26961 -40896
rect 26589 -41172 26653 -40928
rect 26897 -41172 26961 -40928
rect 26589 -41204 26961 -41172
rect 27589 -40928 27961 -40896
rect 27589 -41172 27653 -40928
rect 27897 -41172 27961 -40928
rect 27589 -41204 27961 -41172
rect 28589 -40928 28961 -40896
rect 28589 -41172 28653 -40928
rect 28897 -41172 28961 -40928
rect 28589 -41204 28961 -41172
rect 29589 -40928 29961 -40896
rect 29589 -41172 29653 -40928
rect 29897 -41172 29961 -40928
rect 29589 -41204 29961 -41172
rect 30589 -40928 30961 -40896
rect 30589 -41172 30653 -40928
rect 30897 -41172 30961 -40928
rect 30589 -41204 30961 -41172
rect 31589 -40928 31961 -40896
rect 31589 -41172 31653 -40928
rect 31897 -41172 31961 -40928
rect 31589 -41204 31961 -41172
rect 32589 -40928 32961 -40896
rect 32589 -41172 32653 -40928
rect 32897 -41172 32961 -40928
rect 32589 -41204 32961 -41172
rect 33589 -40928 33961 -40896
rect 33589 -41172 33653 -40928
rect 33897 -41172 33961 -40928
rect 33589 -41204 33961 -41172
rect 34269 -41204 34275 -40896
rect 8275 -41210 34275 -41204
rect 8615 -41236 8935 -41210
rect 8615 -41864 8621 -41236
rect 8929 -41864 8935 -41236
rect 8615 -41890 8935 -41864
rect 9615 -41236 9935 -41210
rect 9615 -41864 9621 -41236
rect 9929 -41864 9935 -41236
rect 9615 -41890 9935 -41864
rect 10615 -41236 10935 -41210
rect 10615 -41864 10621 -41236
rect 10929 -41864 10935 -41236
rect 10615 -41890 10935 -41864
rect 11615 -41236 11935 -41210
rect 11615 -41864 11621 -41236
rect 11929 -41864 11935 -41236
rect 11615 -41890 11935 -41864
rect 12615 -41236 12935 -41210
rect 12615 -41864 12621 -41236
rect 12929 -41864 12935 -41236
rect 12615 -41890 12935 -41864
rect 13615 -41236 13935 -41210
rect 13615 -41864 13621 -41236
rect 13929 -41864 13935 -41236
rect 13615 -41890 13935 -41864
rect 14615 -41236 14935 -41210
rect 14615 -41864 14621 -41236
rect 14929 -41864 14935 -41236
rect 14615 -41890 14935 -41864
rect 15615 -41236 15935 -41210
rect 15615 -41864 15621 -41236
rect 15929 -41864 15935 -41236
rect 15615 -41890 15935 -41864
rect 16615 -41236 16935 -41210
rect 16615 -41864 16621 -41236
rect 16929 -41864 16935 -41236
rect 16615 -41890 16935 -41864
rect 17615 -41236 17935 -41210
rect 17615 -41864 17621 -41236
rect 17929 -41864 17935 -41236
rect 17615 -41890 17935 -41864
rect 18615 -41236 18935 -41210
rect 18615 -41864 18621 -41236
rect 18929 -41864 18935 -41236
rect 18615 -41890 18935 -41864
rect 19615 -41236 19935 -41210
rect 19615 -41864 19621 -41236
rect 19929 -41864 19935 -41236
rect 19615 -41890 19935 -41864
rect 20615 -41236 20935 -41210
rect 20615 -41864 20621 -41236
rect 20929 -41864 20935 -41236
rect 20615 -41890 20935 -41864
rect 21615 -41236 21935 -41210
rect 21615 -41864 21621 -41236
rect 21929 -41864 21935 -41236
rect 21615 -41890 21935 -41864
rect 22615 -41236 22935 -41210
rect 22615 -41864 22621 -41236
rect 22929 -41864 22935 -41236
rect 22615 -41890 22935 -41864
rect 23615 -41236 23935 -41210
rect 23615 -41864 23621 -41236
rect 23929 -41864 23935 -41236
rect 23615 -41890 23935 -41864
rect 24615 -41236 24935 -41210
rect 24615 -41864 24621 -41236
rect 24929 -41864 24935 -41236
rect 24615 -41890 24935 -41864
rect 25615 -41236 25935 -41210
rect 25615 -41864 25621 -41236
rect 25929 -41864 25935 -41236
rect 25615 -41890 25935 -41864
rect 26615 -41236 26935 -41210
rect 26615 -41864 26621 -41236
rect 26929 -41864 26935 -41236
rect 26615 -41890 26935 -41864
rect 27615 -41236 27935 -41210
rect 27615 -41864 27621 -41236
rect 27929 -41864 27935 -41236
rect 27615 -41890 27935 -41864
rect 28615 -41236 28935 -41210
rect 28615 -41864 28621 -41236
rect 28929 -41864 28935 -41236
rect 28615 -41890 28935 -41864
rect 29615 -41236 29935 -41210
rect 29615 -41864 29621 -41236
rect 29929 -41864 29935 -41236
rect 29615 -41890 29935 -41864
rect 30615 -41236 30935 -41210
rect 30615 -41864 30621 -41236
rect 30929 -41864 30935 -41236
rect 30615 -41890 30935 -41864
rect 31615 -41236 31935 -41210
rect 31615 -41864 31621 -41236
rect 31929 -41864 31935 -41236
rect 31615 -41890 31935 -41864
rect 32615 -41236 32935 -41210
rect 32615 -41864 32621 -41236
rect 32929 -41864 32935 -41236
rect 32615 -41890 32935 -41864
rect 33615 -41236 33935 -41210
rect 33615 -41864 33621 -41236
rect 33929 -41864 33935 -41236
rect 33615 -41890 33935 -41864
rect 8275 -41896 34275 -41890
rect 8275 -42204 8281 -41896
rect 8589 -41928 8961 -41896
rect 8589 -42172 8653 -41928
rect 8897 -42172 8961 -41928
rect 8589 -42204 8961 -42172
rect 9589 -41928 9961 -41896
rect 9589 -42172 9653 -41928
rect 9897 -42172 9961 -41928
rect 9589 -42204 9961 -42172
rect 10589 -41928 10961 -41896
rect 10589 -42172 10653 -41928
rect 10897 -42172 10961 -41928
rect 10589 -42204 10961 -42172
rect 11589 -41928 11961 -41896
rect 11589 -42172 11653 -41928
rect 11897 -42172 11961 -41928
rect 11589 -42204 11961 -42172
rect 12589 -41928 12961 -41896
rect 12589 -42172 12653 -41928
rect 12897 -42172 12961 -41928
rect 12589 -42204 12961 -42172
rect 13589 -41928 13961 -41896
rect 13589 -42172 13653 -41928
rect 13897 -42172 13961 -41928
rect 13589 -42204 13961 -42172
rect 14589 -41928 14961 -41896
rect 14589 -42172 14653 -41928
rect 14897 -42172 14961 -41928
rect 14589 -42204 14961 -42172
rect 15589 -41928 15961 -41896
rect 15589 -42172 15653 -41928
rect 15897 -42172 15961 -41928
rect 15589 -42204 15961 -42172
rect 16589 -41928 16961 -41896
rect 16589 -42172 16653 -41928
rect 16897 -42172 16961 -41928
rect 16589 -42204 16961 -42172
rect 17589 -41928 17961 -41896
rect 17589 -42172 17653 -41928
rect 17897 -42172 17961 -41928
rect 17589 -42204 17961 -42172
rect 18589 -41928 18961 -41896
rect 18589 -42172 18653 -41928
rect 18897 -42172 18961 -41928
rect 18589 -42204 18961 -42172
rect 19589 -41928 19961 -41896
rect 19589 -42172 19653 -41928
rect 19897 -42172 19961 -41928
rect 19589 -42204 19961 -42172
rect 20589 -41928 20961 -41896
rect 20589 -42172 20653 -41928
rect 20897 -42172 20961 -41928
rect 20589 -42204 20961 -42172
rect 21589 -41928 21961 -41896
rect 21589 -42172 21653 -41928
rect 21897 -42172 21961 -41928
rect 21589 -42204 21961 -42172
rect 22589 -41928 22961 -41896
rect 22589 -42172 22653 -41928
rect 22897 -42172 22961 -41928
rect 22589 -42204 22961 -42172
rect 23589 -41928 23961 -41896
rect 23589 -42172 23653 -41928
rect 23897 -42172 23961 -41928
rect 23589 -42204 23961 -42172
rect 24589 -41928 24961 -41896
rect 24589 -42172 24653 -41928
rect 24897 -42172 24961 -41928
rect 24589 -42204 24961 -42172
rect 25589 -41928 25961 -41896
rect 25589 -42172 25653 -41928
rect 25897 -42172 25961 -41928
rect 25589 -42204 25961 -42172
rect 26589 -41928 26961 -41896
rect 26589 -42172 26653 -41928
rect 26897 -42172 26961 -41928
rect 26589 -42204 26961 -42172
rect 27589 -41928 27961 -41896
rect 27589 -42172 27653 -41928
rect 27897 -42172 27961 -41928
rect 27589 -42204 27961 -42172
rect 28589 -41928 28961 -41896
rect 28589 -42172 28653 -41928
rect 28897 -42172 28961 -41928
rect 28589 -42204 28961 -42172
rect 29589 -41928 29961 -41896
rect 29589 -42172 29653 -41928
rect 29897 -42172 29961 -41928
rect 29589 -42204 29961 -42172
rect 30589 -41928 30961 -41896
rect 30589 -42172 30653 -41928
rect 30897 -42172 30961 -41928
rect 30589 -42204 30961 -42172
rect 31589 -41928 31961 -41896
rect 31589 -42172 31653 -41928
rect 31897 -42172 31961 -41928
rect 31589 -42204 31961 -42172
rect 32589 -41928 32961 -41896
rect 32589 -42172 32653 -41928
rect 32897 -42172 32961 -41928
rect 32589 -42204 32961 -42172
rect 33589 -41928 33961 -41896
rect 33589 -42172 33653 -41928
rect 33897 -42172 33961 -41928
rect 33589 -42204 33961 -42172
rect 34269 -42204 34275 -41896
rect 8275 -42210 34275 -42204
rect 8615 -42236 8935 -42210
rect 8615 -42864 8621 -42236
rect 8929 -42864 8935 -42236
rect 8615 -42890 8935 -42864
rect 9615 -42236 9935 -42210
rect 9615 -42864 9621 -42236
rect 9929 -42864 9935 -42236
rect 9615 -42890 9935 -42864
rect 10615 -42236 10935 -42210
rect 10615 -42864 10621 -42236
rect 10929 -42864 10935 -42236
rect 10615 -42890 10935 -42864
rect 11615 -42236 11935 -42210
rect 11615 -42864 11621 -42236
rect 11929 -42864 11935 -42236
rect 11615 -42890 11935 -42864
rect 12615 -42236 12935 -42210
rect 12615 -42864 12621 -42236
rect 12929 -42864 12935 -42236
rect 12615 -42890 12935 -42864
rect 13615 -42236 13935 -42210
rect 13615 -42864 13621 -42236
rect 13929 -42864 13935 -42236
rect 13615 -42890 13935 -42864
rect 14615 -42236 14935 -42210
rect 14615 -42864 14621 -42236
rect 14929 -42864 14935 -42236
rect 14615 -42890 14935 -42864
rect 15615 -42236 15935 -42210
rect 15615 -42864 15621 -42236
rect 15929 -42864 15935 -42236
rect 15615 -42890 15935 -42864
rect 16615 -42236 16935 -42210
rect 16615 -42864 16621 -42236
rect 16929 -42864 16935 -42236
rect 16615 -42890 16935 -42864
rect 17615 -42236 17935 -42210
rect 17615 -42864 17621 -42236
rect 17929 -42864 17935 -42236
rect 17615 -42890 17935 -42864
rect 18615 -42236 18935 -42210
rect 18615 -42864 18621 -42236
rect 18929 -42864 18935 -42236
rect 18615 -42890 18935 -42864
rect 19615 -42236 19935 -42210
rect 19615 -42864 19621 -42236
rect 19929 -42864 19935 -42236
rect 19615 -42890 19935 -42864
rect 20615 -42236 20935 -42210
rect 20615 -42864 20621 -42236
rect 20929 -42864 20935 -42236
rect 20615 -42890 20935 -42864
rect 21615 -42236 21935 -42210
rect 21615 -42864 21621 -42236
rect 21929 -42864 21935 -42236
rect 21615 -42890 21935 -42864
rect 22615 -42236 22935 -42210
rect 22615 -42864 22621 -42236
rect 22929 -42864 22935 -42236
rect 22615 -42890 22935 -42864
rect 23615 -42236 23935 -42210
rect 23615 -42864 23621 -42236
rect 23929 -42864 23935 -42236
rect 23615 -42890 23935 -42864
rect 24615 -42236 24935 -42210
rect 24615 -42864 24621 -42236
rect 24929 -42864 24935 -42236
rect 24615 -42890 24935 -42864
rect 25615 -42236 25935 -42210
rect 25615 -42864 25621 -42236
rect 25929 -42864 25935 -42236
rect 25615 -42890 25935 -42864
rect 26615 -42236 26935 -42210
rect 26615 -42864 26621 -42236
rect 26929 -42864 26935 -42236
rect 26615 -42890 26935 -42864
rect 27615 -42236 27935 -42210
rect 27615 -42864 27621 -42236
rect 27929 -42864 27935 -42236
rect 27615 -42890 27935 -42864
rect 28615 -42236 28935 -42210
rect 28615 -42864 28621 -42236
rect 28929 -42864 28935 -42236
rect 28615 -42890 28935 -42864
rect 29615 -42236 29935 -42210
rect 29615 -42864 29621 -42236
rect 29929 -42864 29935 -42236
rect 29615 -42890 29935 -42864
rect 30615 -42236 30935 -42210
rect 30615 -42864 30621 -42236
rect 30929 -42864 30935 -42236
rect 30615 -42890 30935 -42864
rect 31615 -42236 31935 -42210
rect 31615 -42864 31621 -42236
rect 31929 -42864 31935 -42236
rect 31615 -42890 31935 -42864
rect 32615 -42236 32935 -42210
rect 32615 -42864 32621 -42236
rect 32929 -42864 32935 -42236
rect 32615 -42890 32935 -42864
rect 33615 -42236 33935 -42210
rect 33615 -42864 33621 -42236
rect 33929 -42864 33935 -42236
rect 33615 -42890 33935 -42864
rect 8275 -42896 34275 -42890
rect 8275 -43204 8281 -42896
rect 8589 -42928 8961 -42896
rect 8589 -43172 8653 -42928
rect 8897 -43172 8961 -42928
rect 8589 -43204 8961 -43172
rect 9589 -42928 9961 -42896
rect 9589 -43172 9653 -42928
rect 9897 -43172 9961 -42928
rect 9589 -43204 9961 -43172
rect 10589 -42928 10961 -42896
rect 10589 -43172 10653 -42928
rect 10897 -43172 10961 -42928
rect 10589 -43204 10961 -43172
rect 11589 -42928 11961 -42896
rect 11589 -43172 11653 -42928
rect 11897 -43172 11961 -42928
rect 11589 -43204 11961 -43172
rect 12589 -42928 12961 -42896
rect 12589 -43172 12653 -42928
rect 12897 -43172 12961 -42928
rect 12589 -43204 12961 -43172
rect 13589 -42928 13961 -42896
rect 13589 -43172 13653 -42928
rect 13897 -43172 13961 -42928
rect 13589 -43204 13961 -43172
rect 14589 -42928 14961 -42896
rect 14589 -43172 14653 -42928
rect 14897 -43172 14961 -42928
rect 14589 -43204 14961 -43172
rect 15589 -42928 15961 -42896
rect 15589 -43172 15653 -42928
rect 15897 -43172 15961 -42928
rect 15589 -43204 15961 -43172
rect 16589 -42928 16961 -42896
rect 16589 -43172 16653 -42928
rect 16897 -43172 16961 -42928
rect 16589 -43204 16961 -43172
rect 17589 -42928 17961 -42896
rect 17589 -43172 17653 -42928
rect 17897 -43172 17961 -42928
rect 17589 -43204 17961 -43172
rect 18589 -42928 18961 -42896
rect 18589 -43172 18653 -42928
rect 18897 -43172 18961 -42928
rect 18589 -43204 18961 -43172
rect 19589 -42928 19961 -42896
rect 19589 -43172 19653 -42928
rect 19897 -43172 19961 -42928
rect 19589 -43204 19961 -43172
rect 20589 -42928 20961 -42896
rect 20589 -43172 20653 -42928
rect 20897 -43172 20961 -42928
rect 20589 -43204 20961 -43172
rect 21589 -42928 21961 -42896
rect 21589 -43172 21653 -42928
rect 21897 -43172 21961 -42928
rect 21589 -43204 21961 -43172
rect 22589 -42928 22961 -42896
rect 22589 -43172 22653 -42928
rect 22897 -43172 22961 -42928
rect 22589 -43204 22961 -43172
rect 23589 -42928 23961 -42896
rect 23589 -43172 23653 -42928
rect 23897 -43172 23961 -42928
rect 23589 -43204 23961 -43172
rect 24589 -42928 24961 -42896
rect 24589 -43172 24653 -42928
rect 24897 -43172 24961 -42928
rect 24589 -43204 24961 -43172
rect 25589 -42928 25961 -42896
rect 25589 -43172 25653 -42928
rect 25897 -43172 25961 -42928
rect 25589 -43204 25961 -43172
rect 26589 -42928 26961 -42896
rect 26589 -43172 26653 -42928
rect 26897 -43172 26961 -42928
rect 26589 -43204 26961 -43172
rect 27589 -42928 27961 -42896
rect 27589 -43172 27653 -42928
rect 27897 -43172 27961 -42928
rect 27589 -43204 27961 -43172
rect 28589 -42928 28961 -42896
rect 28589 -43172 28653 -42928
rect 28897 -43172 28961 -42928
rect 28589 -43204 28961 -43172
rect 29589 -42928 29961 -42896
rect 29589 -43172 29653 -42928
rect 29897 -43172 29961 -42928
rect 29589 -43204 29961 -43172
rect 30589 -42928 30961 -42896
rect 30589 -43172 30653 -42928
rect 30897 -43172 30961 -42928
rect 30589 -43204 30961 -43172
rect 31589 -42928 31961 -42896
rect 31589 -43172 31653 -42928
rect 31897 -43172 31961 -42928
rect 31589 -43204 31961 -43172
rect 32589 -42928 32961 -42896
rect 32589 -43172 32653 -42928
rect 32897 -43172 32961 -42928
rect 32589 -43204 32961 -43172
rect 33589 -42928 33961 -42896
rect 33589 -43172 33653 -42928
rect 33897 -43172 33961 -42928
rect 33589 -43204 33961 -43172
rect 34269 -43204 34275 -42896
rect 8275 -43210 34275 -43204
rect 8615 -43236 8935 -43210
rect 8615 -43864 8621 -43236
rect 8929 -43864 8935 -43236
rect 8615 -43890 8935 -43864
rect 9615 -43236 9935 -43210
rect 9615 -43864 9621 -43236
rect 9929 -43864 9935 -43236
rect 9615 -43890 9935 -43864
rect 10615 -43236 10935 -43210
rect 10615 -43864 10621 -43236
rect 10929 -43864 10935 -43236
rect 10615 -43890 10935 -43864
rect 11615 -43236 11935 -43210
rect 11615 -43864 11621 -43236
rect 11929 -43864 11935 -43236
rect 11615 -43890 11935 -43864
rect 12615 -43236 12935 -43210
rect 12615 -43864 12621 -43236
rect 12929 -43864 12935 -43236
rect 12615 -43890 12935 -43864
rect 13615 -43236 13935 -43210
rect 13615 -43864 13621 -43236
rect 13929 -43864 13935 -43236
rect 13615 -43890 13935 -43864
rect 14615 -43236 14935 -43210
rect 14615 -43864 14621 -43236
rect 14929 -43864 14935 -43236
rect 14615 -43890 14935 -43864
rect 15615 -43236 15935 -43210
rect 15615 -43864 15621 -43236
rect 15929 -43864 15935 -43236
rect 15615 -43890 15935 -43864
rect 16615 -43236 16935 -43210
rect 16615 -43864 16621 -43236
rect 16929 -43864 16935 -43236
rect 16615 -43890 16935 -43864
rect 17615 -43236 17935 -43210
rect 17615 -43864 17621 -43236
rect 17929 -43864 17935 -43236
rect 17615 -43890 17935 -43864
rect 18615 -43236 18935 -43210
rect 18615 -43864 18621 -43236
rect 18929 -43864 18935 -43236
rect 18615 -43890 18935 -43864
rect 19615 -43236 19935 -43210
rect 19615 -43864 19621 -43236
rect 19929 -43864 19935 -43236
rect 19615 -43890 19935 -43864
rect 20615 -43236 20935 -43210
rect 20615 -43864 20621 -43236
rect 20929 -43864 20935 -43236
rect 20615 -43890 20935 -43864
rect 21615 -43236 21935 -43210
rect 21615 -43864 21621 -43236
rect 21929 -43864 21935 -43236
rect 21615 -43890 21935 -43864
rect 22615 -43236 22935 -43210
rect 22615 -43864 22621 -43236
rect 22929 -43864 22935 -43236
rect 22615 -43890 22935 -43864
rect 23615 -43236 23935 -43210
rect 23615 -43864 23621 -43236
rect 23929 -43864 23935 -43236
rect 23615 -43890 23935 -43864
rect 24615 -43236 24935 -43210
rect 24615 -43864 24621 -43236
rect 24929 -43864 24935 -43236
rect 24615 -43890 24935 -43864
rect 25615 -43236 25935 -43210
rect 25615 -43864 25621 -43236
rect 25929 -43864 25935 -43236
rect 25615 -43890 25935 -43864
rect 26615 -43236 26935 -43210
rect 26615 -43864 26621 -43236
rect 26929 -43864 26935 -43236
rect 26615 -43890 26935 -43864
rect 27615 -43236 27935 -43210
rect 27615 -43864 27621 -43236
rect 27929 -43864 27935 -43236
rect 27615 -43890 27935 -43864
rect 28615 -43236 28935 -43210
rect 28615 -43864 28621 -43236
rect 28929 -43864 28935 -43236
rect 28615 -43890 28935 -43864
rect 29615 -43236 29935 -43210
rect 29615 -43864 29621 -43236
rect 29929 -43864 29935 -43236
rect 29615 -43890 29935 -43864
rect 30615 -43236 30935 -43210
rect 30615 -43864 30621 -43236
rect 30929 -43864 30935 -43236
rect 30615 -43890 30935 -43864
rect 31615 -43236 31935 -43210
rect 31615 -43864 31621 -43236
rect 31929 -43864 31935 -43236
rect 31615 -43890 31935 -43864
rect 32615 -43236 32935 -43210
rect 32615 -43864 32621 -43236
rect 32929 -43864 32935 -43236
rect 32615 -43890 32935 -43864
rect 33615 -43236 33935 -43210
rect 33615 -43864 33621 -43236
rect 33929 -43864 33935 -43236
rect 33615 -43890 33935 -43864
rect 8275 -43896 34275 -43890
rect 8275 -44204 8281 -43896
rect 8589 -43928 8961 -43896
rect 8589 -44172 8653 -43928
rect 8897 -44172 8961 -43928
rect 8589 -44204 8961 -44172
rect 9589 -43928 9961 -43896
rect 9589 -44172 9653 -43928
rect 9897 -44172 9961 -43928
rect 9589 -44204 9961 -44172
rect 10589 -43928 10961 -43896
rect 10589 -44172 10653 -43928
rect 10897 -44172 10961 -43928
rect 10589 -44204 10961 -44172
rect 11589 -43928 11961 -43896
rect 11589 -44172 11653 -43928
rect 11897 -44172 11961 -43928
rect 11589 -44204 11961 -44172
rect 12589 -43928 12961 -43896
rect 12589 -44172 12653 -43928
rect 12897 -44172 12961 -43928
rect 12589 -44204 12961 -44172
rect 13589 -43928 13961 -43896
rect 13589 -44172 13653 -43928
rect 13897 -44172 13961 -43928
rect 13589 -44204 13961 -44172
rect 14589 -43928 14961 -43896
rect 14589 -44172 14653 -43928
rect 14897 -44172 14961 -43928
rect 14589 -44204 14961 -44172
rect 15589 -43928 15961 -43896
rect 15589 -44172 15653 -43928
rect 15897 -44172 15961 -43928
rect 15589 -44204 15961 -44172
rect 16589 -43928 16961 -43896
rect 16589 -44172 16653 -43928
rect 16897 -44172 16961 -43928
rect 16589 -44204 16961 -44172
rect 17589 -43928 17961 -43896
rect 17589 -44172 17653 -43928
rect 17897 -44172 17961 -43928
rect 17589 -44204 17961 -44172
rect 18589 -43928 18961 -43896
rect 18589 -44172 18653 -43928
rect 18897 -44172 18961 -43928
rect 18589 -44204 18961 -44172
rect 19589 -43928 19961 -43896
rect 19589 -44172 19653 -43928
rect 19897 -44172 19961 -43928
rect 19589 -44204 19961 -44172
rect 20589 -43928 20961 -43896
rect 20589 -44172 20653 -43928
rect 20897 -44172 20961 -43928
rect 20589 -44204 20961 -44172
rect 21589 -43928 21961 -43896
rect 21589 -44172 21653 -43928
rect 21897 -44172 21961 -43928
rect 21589 -44204 21961 -44172
rect 22589 -43928 22961 -43896
rect 22589 -44172 22653 -43928
rect 22897 -44172 22961 -43928
rect 22589 -44204 22961 -44172
rect 23589 -43928 23961 -43896
rect 23589 -44172 23653 -43928
rect 23897 -44172 23961 -43928
rect 23589 -44204 23961 -44172
rect 24589 -43928 24961 -43896
rect 24589 -44172 24653 -43928
rect 24897 -44172 24961 -43928
rect 24589 -44204 24961 -44172
rect 25589 -43928 25961 -43896
rect 25589 -44172 25653 -43928
rect 25897 -44172 25961 -43928
rect 25589 -44204 25961 -44172
rect 26589 -43928 26961 -43896
rect 26589 -44172 26653 -43928
rect 26897 -44172 26961 -43928
rect 26589 -44204 26961 -44172
rect 27589 -43928 27961 -43896
rect 27589 -44172 27653 -43928
rect 27897 -44172 27961 -43928
rect 27589 -44204 27961 -44172
rect 28589 -43928 28961 -43896
rect 28589 -44172 28653 -43928
rect 28897 -44172 28961 -43928
rect 28589 -44204 28961 -44172
rect 29589 -43928 29961 -43896
rect 29589 -44172 29653 -43928
rect 29897 -44172 29961 -43928
rect 29589 -44204 29961 -44172
rect 30589 -43928 30961 -43896
rect 30589 -44172 30653 -43928
rect 30897 -44172 30961 -43928
rect 30589 -44204 30961 -44172
rect 31589 -43928 31961 -43896
rect 31589 -44172 31653 -43928
rect 31897 -44172 31961 -43928
rect 31589 -44204 31961 -44172
rect 32589 -43928 32961 -43896
rect 32589 -44172 32653 -43928
rect 32897 -44172 32961 -43928
rect 32589 -44204 32961 -44172
rect 33589 -43928 33961 -43896
rect 33589 -44172 33653 -43928
rect 33897 -44172 33961 -43928
rect 33589 -44204 33961 -44172
rect 34269 -44204 34275 -43896
rect 8275 -44210 34275 -44204
rect -46275 -44550 5725 -44496
rect 8615 -44236 8935 -44210
rect -49485 -44890 -49165 -44864
rect 8615 -44864 8621 -44236
rect 8929 -44864 8935 -44236
rect 8615 -44890 8935 -44864
rect 9615 -44236 9935 -44210
rect 9615 -44864 9621 -44236
rect 9929 -44864 9935 -44236
rect 9615 -44890 9935 -44864
rect 10615 -44236 10935 -44210
rect 10615 -44864 10621 -44236
rect 10929 -44864 10935 -44236
rect 10615 -44890 10935 -44864
rect 11615 -44236 11935 -44210
rect 11615 -44864 11621 -44236
rect 11929 -44864 11935 -44236
rect 11615 -44890 11935 -44864
rect 12615 -44236 12935 -44210
rect 12615 -44864 12621 -44236
rect 12929 -44864 12935 -44236
rect 12615 -44890 12935 -44864
rect 13615 -44236 13935 -44210
rect 13615 -44864 13621 -44236
rect 13929 -44864 13935 -44236
rect 13615 -44890 13935 -44864
rect 14615 -44236 14935 -44210
rect 14615 -44864 14621 -44236
rect 14929 -44864 14935 -44236
rect 14615 -44890 14935 -44864
rect 15615 -44236 15935 -44210
rect 15615 -44864 15621 -44236
rect 15929 -44864 15935 -44236
rect 15615 -44890 15935 -44864
rect 16615 -44236 16935 -44210
rect 16615 -44864 16621 -44236
rect 16929 -44864 16935 -44236
rect 16615 -44890 16935 -44864
rect 17615 -44236 17935 -44210
rect 17615 -44864 17621 -44236
rect 17929 -44864 17935 -44236
rect 17615 -44890 17935 -44864
rect 18615 -44236 18935 -44210
rect 18615 -44864 18621 -44236
rect 18929 -44864 18935 -44236
rect 18615 -44890 18935 -44864
rect 19615 -44236 19935 -44210
rect 19615 -44864 19621 -44236
rect 19929 -44864 19935 -44236
rect 19615 -44890 19935 -44864
rect 20615 -44236 20935 -44210
rect 20615 -44864 20621 -44236
rect 20929 -44864 20935 -44236
rect 20615 -44890 20935 -44864
rect 21615 -44236 21935 -44210
rect 21615 -44864 21621 -44236
rect 21929 -44864 21935 -44236
rect 21615 -44890 21935 -44864
rect 22615 -44236 22935 -44210
rect 22615 -44864 22621 -44236
rect 22929 -44864 22935 -44236
rect 22615 -44890 22935 -44864
rect 23615 -44236 23935 -44210
rect 23615 -44864 23621 -44236
rect 23929 -44864 23935 -44236
rect 23615 -44890 23935 -44864
rect 24615 -44236 24935 -44210
rect 24615 -44864 24621 -44236
rect 24929 -44864 24935 -44236
rect 24615 -44890 24935 -44864
rect 25615 -44236 25935 -44210
rect 25615 -44864 25621 -44236
rect 25929 -44864 25935 -44236
rect 25615 -44890 25935 -44864
rect 26615 -44236 26935 -44210
rect 26615 -44864 26621 -44236
rect 26929 -44864 26935 -44236
rect 26615 -44890 26935 -44864
rect 27615 -44236 27935 -44210
rect 27615 -44864 27621 -44236
rect 27929 -44864 27935 -44236
rect 27615 -44890 27935 -44864
rect 28615 -44236 28935 -44210
rect 28615 -44864 28621 -44236
rect 28929 -44864 28935 -44236
rect 28615 -44890 28935 -44864
rect 29615 -44236 29935 -44210
rect 29615 -44864 29621 -44236
rect 29929 -44864 29935 -44236
rect 29615 -44890 29935 -44864
rect 30615 -44236 30935 -44210
rect 30615 -44864 30621 -44236
rect 30929 -44864 30935 -44236
rect 30615 -44890 30935 -44864
rect 31615 -44236 31935 -44210
rect 31615 -44864 31621 -44236
rect 31929 -44864 31935 -44236
rect 31615 -44890 31935 -44864
rect 32615 -44236 32935 -44210
rect 32615 -44864 32621 -44236
rect 32929 -44864 32935 -44236
rect 32615 -44890 32935 -44864
rect 33615 -44236 33935 -44210
rect 33615 -44864 33621 -44236
rect 33929 -44864 33935 -44236
rect 33615 -44890 33935 -44864
rect -74825 -44896 -48825 -44890
rect -74825 -45204 -74819 -44896
rect -74511 -44928 -74139 -44896
rect -74511 -45172 -74447 -44928
rect -74203 -45172 -74139 -44928
rect -74511 -45204 -74139 -45172
rect -73511 -44928 -73139 -44896
rect -73511 -45172 -73447 -44928
rect -73203 -45172 -73139 -44928
rect -73511 -45204 -73139 -45172
rect -72511 -44928 -72139 -44896
rect -72511 -45172 -72447 -44928
rect -72203 -45172 -72139 -44928
rect -72511 -45204 -72139 -45172
rect -71511 -44928 -71139 -44896
rect -71511 -45172 -71447 -44928
rect -71203 -45172 -71139 -44928
rect -71511 -45204 -71139 -45172
rect -70511 -44928 -70139 -44896
rect -70511 -45172 -70447 -44928
rect -70203 -45172 -70139 -44928
rect -70511 -45204 -70139 -45172
rect -69511 -44928 -69139 -44896
rect -69511 -45172 -69447 -44928
rect -69203 -45172 -69139 -44928
rect -69511 -45204 -69139 -45172
rect -68511 -44928 -68139 -44896
rect -68511 -45172 -68447 -44928
rect -68203 -45172 -68139 -44928
rect -68511 -45204 -68139 -45172
rect -67511 -44928 -67139 -44896
rect -67511 -45172 -67447 -44928
rect -67203 -45172 -67139 -44928
rect -67511 -45204 -67139 -45172
rect -66511 -44928 -66139 -44896
rect -66511 -45172 -66447 -44928
rect -66203 -45172 -66139 -44928
rect -66511 -45204 -66139 -45172
rect -65511 -44928 -65139 -44896
rect -65511 -45172 -65447 -44928
rect -65203 -45172 -65139 -44928
rect -65511 -45204 -65139 -45172
rect -64511 -44928 -64139 -44896
rect -64511 -45172 -64447 -44928
rect -64203 -45172 -64139 -44928
rect -64511 -45204 -64139 -45172
rect -63511 -44928 -63139 -44896
rect -63511 -45172 -63447 -44928
rect -63203 -45172 -63139 -44928
rect -63511 -45204 -63139 -45172
rect -62511 -44928 -62139 -44896
rect -62511 -45172 -62447 -44928
rect -62203 -45172 -62139 -44928
rect -62511 -45204 -62139 -45172
rect -61511 -44928 -61139 -44896
rect -61511 -45172 -61447 -44928
rect -61203 -45172 -61139 -44928
rect -61511 -45204 -61139 -45172
rect -60511 -44928 -60139 -44896
rect -60511 -45172 -60447 -44928
rect -60203 -45172 -60139 -44928
rect -60511 -45204 -60139 -45172
rect -59511 -44928 -59139 -44896
rect -59511 -45172 -59447 -44928
rect -59203 -45172 -59139 -44928
rect -59511 -45204 -59139 -45172
rect -58511 -44928 -58139 -44896
rect -58511 -45172 -58447 -44928
rect -58203 -45172 -58139 -44928
rect -58511 -45204 -58139 -45172
rect -57511 -44928 -57139 -44896
rect -57511 -45172 -57447 -44928
rect -57203 -45172 -57139 -44928
rect -57511 -45204 -57139 -45172
rect -56511 -44928 -56139 -44896
rect -56511 -45172 -56447 -44928
rect -56203 -45172 -56139 -44928
rect -56511 -45204 -56139 -45172
rect -55511 -44928 -55139 -44896
rect -55511 -45172 -55447 -44928
rect -55203 -45172 -55139 -44928
rect -55511 -45204 -55139 -45172
rect -54511 -44928 -54139 -44896
rect -54511 -45172 -54447 -44928
rect -54203 -45172 -54139 -44928
rect -54511 -45204 -54139 -45172
rect -53511 -44928 -53139 -44896
rect -53511 -45172 -53447 -44928
rect -53203 -45172 -53139 -44928
rect -53511 -45204 -53139 -45172
rect -52511 -44928 -52139 -44896
rect -52511 -45172 -52447 -44928
rect -52203 -45172 -52139 -44928
rect -52511 -45204 -52139 -45172
rect -51511 -44928 -51139 -44896
rect -51511 -45172 -51447 -44928
rect -51203 -45172 -51139 -44928
rect -51511 -45204 -51139 -45172
rect -50511 -44928 -50139 -44896
rect -50511 -45172 -50447 -44928
rect -50203 -45172 -50139 -44928
rect -50511 -45204 -50139 -45172
rect -49511 -44928 -49139 -44896
rect -49511 -45172 -49447 -44928
rect -49203 -45172 -49139 -44928
rect -49511 -45204 -49139 -45172
rect -48831 -45204 -48825 -44896
rect -74825 -45210 -48825 -45204
rect 8275 -44896 34275 -44890
rect 8275 -45204 8281 -44896
rect 8589 -44928 8961 -44896
rect 8589 -45172 8653 -44928
rect 8897 -45172 8961 -44928
rect 8589 -45204 8961 -45172
rect 9589 -44928 9961 -44896
rect 9589 -45172 9653 -44928
rect 9897 -45172 9961 -44928
rect 9589 -45204 9961 -45172
rect 10589 -44928 10961 -44896
rect 10589 -45172 10653 -44928
rect 10897 -45172 10961 -44928
rect 10589 -45204 10961 -45172
rect 11589 -44928 11961 -44896
rect 11589 -45172 11653 -44928
rect 11897 -45172 11961 -44928
rect 11589 -45204 11961 -45172
rect 12589 -44928 12961 -44896
rect 12589 -45172 12653 -44928
rect 12897 -45172 12961 -44928
rect 12589 -45204 12961 -45172
rect 13589 -44928 13961 -44896
rect 13589 -45172 13653 -44928
rect 13897 -45172 13961 -44928
rect 13589 -45204 13961 -45172
rect 14589 -44928 14961 -44896
rect 14589 -45172 14653 -44928
rect 14897 -45172 14961 -44928
rect 14589 -45204 14961 -45172
rect 15589 -44928 15961 -44896
rect 15589 -45172 15653 -44928
rect 15897 -45172 15961 -44928
rect 15589 -45204 15961 -45172
rect 16589 -44928 16961 -44896
rect 16589 -45172 16653 -44928
rect 16897 -45172 16961 -44928
rect 16589 -45204 16961 -45172
rect 17589 -44928 17961 -44896
rect 17589 -45172 17653 -44928
rect 17897 -45172 17961 -44928
rect 17589 -45204 17961 -45172
rect 18589 -44928 18961 -44896
rect 18589 -45172 18653 -44928
rect 18897 -45172 18961 -44928
rect 18589 -45204 18961 -45172
rect 19589 -44928 19961 -44896
rect 19589 -45172 19653 -44928
rect 19897 -45172 19961 -44928
rect 19589 -45204 19961 -45172
rect 20589 -44928 20961 -44896
rect 20589 -45172 20653 -44928
rect 20897 -45172 20961 -44928
rect 20589 -45204 20961 -45172
rect 21589 -44928 21961 -44896
rect 21589 -45172 21653 -44928
rect 21897 -45172 21961 -44928
rect 21589 -45204 21961 -45172
rect 22589 -44928 22961 -44896
rect 22589 -45172 22653 -44928
rect 22897 -45172 22961 -44928
rect 22589 -45204 22961 -45172
rect 23589 -44928 23961 -44896
rect 23589 -45172 23653 -44928
rect 23897 -45172 23961 -44928
rect 23589 -45204 23961 -45172
rect 24589 -44928 24961 -44896
rect 24589 -45172 24653 -44928
rect 24897 -45172 24961 -44928
rect 24589 -45204 24961 -45172
rect 25589 -44928 25961 -44896
rect 25589 -45172 25653 -44928
rect 25897 -45172 25961 -44928
rect 25589 -45204 25961 -45172
rect 26589 -44928 26961 -44896
rect 26589 -45172 26653 -44928
rect 26897 -45172 26961 -44928
rect 26589 -45204 26961 -45172
rect 27589 -44928 27961 -44896
rect 27589 -45172 27653 -44928
rect 27897 -45172 27961 -44928
rect 27589 -45204 27961 -45172
rect 28589 -44928 28961 -44896
rect 28589 -45172 28653 -44928
rect 28897 -45172 28961 -44928
rect 28589 -45204 28961 -45172
rect 29589 -44928 29961 -44896
rect 29589 -45172 29653 -44928
rect 29897 -45172 29961 -44928
rect 29589 -45204 29961 -45172
rect 30589 -44928 30961 -44896
rect 30589 -45172 30653 -44928
rect 30897 -45172 30961 -44928
rect 30589 -45204 30961 -45172
rect 31589 -44928 31961 -44896
rect 31589 -45172 31653 -44928
rect 31897 -45172 31961 -44928
rect 31589 -45204 31961 -45172
rect 32589 -44928 32961 -44896
rect 32589 -45172 32653 -44928
rect 32897 -45172 32961 -44928
rect 32589 -45204 32961 -45172
rect 33589 -44928 33961 -44896
rect 33589 -45172 33653 -44928
rect 33897 -45172 33961 -44928
rect 33589 -45204 33961 -45172
rect 34269 -45204 34275 -44896
rect 8275 -45210 34275 -45204
rect -74485 -45236 -74165 -45210
rect -74485 -45864 -74479 -45236
rect -74171 -45864 -74165 -45236
rect -74485 -45890 -74165 -45864
rect -73485 -45236 -73165 -45210
rect -73485 -45864 -73479 -45236
rect -73171 -45864 -73165 -45236
rect -73485 -45890 -73165 -45864
rect -72485 -45236 -72165 -45210
rect -72485 -45864 -72479 -45236
rect -72171 -45864 -72165 -45236
rect -72485 -45890 -72165 -45864
rect -71485 -45236 -71165 -45210
rect -71485 -45864 -71479 -45236
rect -71171 -45864 -71165 -45236
rect -71485 -45890 -71165 -45864
rect -70485 -45236 -70165 -45210
rect -70485 -45864 -70479 -45236
rect -70171 -45864 -70165 -45236
rect -70485 -45890 -70165 -45864
rect -69485 -45236 -69165 -45210
rect -69485 -45864 -69479 -45236
rect -69171 -45864 -69165 -45236
rect -69485 -45890 -69165 -45864
rect -68485 -45236 -68165 -45210
rect -68485 -45864 -68479 -45236
rect -68171 -45864 -68165 -45236
rect -68485 -45890 -68165 -45864
rect -67485 -45236 -67165 -45210
rect -67485 -45864 -67479 -45236
rect -67171 -45864 -67165 -45236
rect -67485 -45890 -67165 -45864
rect -66485 -45236 -66165 -45210
rect -66485 -45864 -66479 -45236
rect -66171 -45864 -66165 -45236
rect -66485 -45890 -66165 -45864
rect -65485 -45236 -65165 -45210
rect -65485 -45864 -65479 -45236
rect -65171 -45864 -65165 -45236
rect -65485 -45890 -65165 -45864
rect -64485 -45236 -64165 -45210
rect -64485 -45864 -64479 -45236
rect -64171 -45864 -64165 -45236
rect -64485 -45890 -64165 -45864
rect -63485 -45236 -63165 -45210
rect -63485 -45864 -63479 -45236
rect -63171 -45864 -63165 -45236
rect -63485 -45890 -63165 -45864
rect -62485 -45236 -62165 -45210
rect -62485 -45864 -62479 -45236
rect -62171 -45864 -62165 -45236
rect -62485 -45890 -62165 -45864
rect -61485 -45236 -61165 -45210
rect -61485 -45864 -61479 -45236
rect -61171 -45864 -61165 -45236
rect -61485 -45890 -61165 -45864
rect -60485 -45236 -60165 -45210
rect -60485 -45864 -60479 -45236
rect -60171 -45864 -60165 -45236
rect -60485 -45890 -60165 -45864
rect -59485 -45236 -59165 -45210
rect -59485 -45864 -59479 -45236
rect -59171 -45864 -59165 -45236
rect -59485 -45890 -59165 -45864
rect -58485 -45236 -58165 -45210
rect -58485 -45864 -58479 -45236
rect -58171 -45864 -58165 -45236
rect -58485 -45890 -58165 -45864
rect -57485 -45236 -57165 -45210
rect -57485 -45864 -57479 -45236
rect -57171 -45864 -57165 -45236
rect -57485 -45890 -57165 -45864
rect -56485 -45236 -56165 -45210
rect -56485 -45864 -56479 -45236
rect -56171 -45864 -56165 -45236
rect -56485 -45890 -56165 -45864
rect -55485 -45236 -55165 -45210
rect -55485 -45864 -55479 -45236
rect -55171 -45864 -55165 -45236
rect -55485 -45890 -55165 -45864
rect -54485 -45236 -54165 -45210
rect -54485 -45864 -54479 -45236
rect -54171 -45864 -54165 -45236
rect -54485 -45890 -54165 -45864
rect -53485 -45236 -53165 -45210
rect -53485 -45864 -53479 -45236
rect -53171 -45864 -53165 -45236
rect -53485 -45890 -53165 -45864
rect -52485 -45236 -52165 -45210
rect -52485 -45864 -52479 -45236
rect -52171 -45864 -52165 -45236
rect -52485 -45890 -52165 -45864
rect -51485 -45236 -51165 -45210
rect -51485 -45864 -51479 -45236
rect -51171 -45864 -51165 -45236
rect -51485 -45890 -51165 -45864
rect -50485 -45236 -50165 -45210
rect -50485 -45864 -50479 -45236
rect -50171 -45864 -50165 -45236
rect -50485 -45890 -50165 -45864
rect -49485 -45236 -49165 -45210
rect -49485 -45864 -49479 -45236
rect -49171 -45864 -49165 -45236
rect -49485 -45890 -49165 -45864
rect 8615 -45236 8935 -45210
rect 8615 -45864 8621 -45236
rect 8929 -45864 8935 -45236
rect 8615 -45890 8935 -45864
rect 9615 -45236 9935 -45210
rect 9615 -45864 9621 -45236
rect 9929 -45864 9935 -45236
rect 9615 -45890 9935 -45864
rect 10615 -45236 10935 -45210
rect 10615 -45864 10621 -45236
rect 10929 -45864 10935 -45236
rect 10615 -45890 10935 -45864
rect 11615 -45236 11935 -45210
rect 11615 -45864 11621 -45236
rect 11929 -45864 11935 -45236
rect 11615 -45890 11935 -45864
rect 12615 -45236 12935 -45210
rect 12615 -45864 12621 -45236
rect 12929 -45864 12935 -45236
rect 12615 -45890 12935 -45864
rect 13615 -45236 13935 -45210
rect 13615 -45864 13621 -45236
rect 13929 -45864 13935 -45236
rect 13615 -45890 13935 -45864
rect 14615 -45236 14935 -45210
rect 14615 -45864 14621 -45236
rect 14929 -45864 14935 -45236
rect 14615 -45890 14935 -45864
rect 15615 -45236 15935 -45210
rect 15615 -45864 15621 -45236
rect 15929 -45864 15935 -45236
rect 15615 -45890 15935 -45864
rect 16615 -45236 16935 -45210
rect 16615 -45864 16621 -45236
rect 16929 -45864 16935 -45236
rect 16615 -45890 16935 -45864
rect 17615 -45236 17935 -45210
rect 17615 -45864 17621 -45236
rect 17929 -45864 17935 -45236
rect 17615 -45890 17935 -45864
rect 18615 -45236 18935 -45210
rect 18615 -45864 18621 -45236
rect 18929 -45864 18935 -45236
rect 18615 -45890 18935 -45864
rect 19615 -45236 19935 -45210
rect 19615 -45864 19621 -45236
rect 19929 -45864 19935 -45236
rect 19615 -45890 19935 -45864
rect 20615 -45236 20935 -45210
rect 20615 -45864 20621 -45236
rect 20929 -45864 20935 -45236
rect 20615 -45890 20935 -45864
rect 21615 -45236 21935 -45210
rect 21615 -45864 21621 -45236
rect 21929 -45864 21935 -45236
rect 21615 -45890 21935 -45864
rect 22615 -45236 22935 -45210
rect 22615 -45864 22621 -45236
rect 22929 -45864 22935 -45236
rect 22615 -45890 22935 -45864
rect 23615 -45236 23935 -45210
rect 23615 -45864 23621 -45236
rect 23929 -45864 23935 -45236
rect 23615 -45890 23935 -45864
rect 24615 -45236 24935 -45210
rect 24615 -45864 24621 -45236
rect 24929 -45864 24935 -45236
rect 24615 -45890 24935 -45864
rect 25615 -45236 25935 -45210
rect 25615 -45864 25621 -45236
rect 25929 -45864 25935 -45236
rect 25615 -45890 25935 -45864
rect 26615 -45236 26935 -45210
rect 26615 -45864 26621 -45236
rect 26929 -45864 26935 -45236
rect 26615 -45890 26935 -45864
rect 27615 -45236 27935 -45210
rect 27615 -45864 27621 -45236
rect 27929 -45864 27935 -45236
rect 27615 -45890 27935 -45864
rect 28615 -45236 28935 -45210
rect 28615 -45864 28621 -45236
rect 28929 -45864 28935 -45236
rect 28615 -45890 28935 -45864
rect 29615 -45236 29935 -45210
rect 29615 -45864 29621 -45236
rect 29929 -45864 29935 -45236
rect 29615 -45890 29935 -45864
rect 30615 -45236 30935 -45210
rect 30615 -45864 30621 -45236
rect 30929 -45864 30935 -45236
rect 30615 -45890 30935 -45864
rect 31615 -45236 31935 -45210
rect 31615 -45864 31621 -45236
rect 31929 -45864 31935 -45236
rect 31615 -45890 31935 -45864
rect 32615 -45236 32935 -45210
rect 32615 -45864 32621 -45236
rect 32929 -45864 32935 -45236
rect 32615 -45890 32935 -45864
rect 33615 -45236 33935 -45210
rect 33615 -45864 33621 -45236
rect 33929 -45864 33935 -45236
rect 33615 -45890 33935 -45864
rect -74825 -45896 -48825 -45890
rect -74825 -46204 -74819 -45896
rect -74511 -45928 -74139 -45896
rect -74511 -46172 -74447 -45928
rect -74203 -46172 -74139 -45928
rect -74511 -46204 -74139 -46172
rect -73511 -45928 -73139 -45896
rect -73511 -46172 -73447 -45928
rect -73203 -46172 -73139 -45928
rect -73511 -46204 -73139 -46172
rect -72511 -45928 -72139 -45896
rect -72511 -46172 -72447 -45928
rect -72203 -46172 -72139 -45928
rect -72511 -46204 -72139 -46172
rect -71511 -45928 -71139 -45896
rect -71511 -46172 -71447 -45928
rect -71203 -46172 -71139 -45928
rect -71511 -46204 -71139 -46172
rect -70511 -45928 -70139 -45896
rect -70511 -46172 -70447 -45928
rect -70203 -46172 -70139 -45928
rect -70511 -46204 -70139 -46172
rect -69511 -45928 -69139 -45896
rect -69511 -46172 -69447 -45928
rect -69203 -46172 -69139 -45928
rect -69511 -46204 -69139 -46172
rect -68511 -45928 -68139 -45896
rect -68511 -46172 -68447 -45928
rect -68203 -46172 -68139 -45928
rect -68511 -46204 -68139 -46172
rect -67511 -45928 -67139 -45896
rect -67511 -46172 -67447 -45928
rect -67203 -46172 -67139 -45928
rect -67511 -46204 -67139 -46172
rect -66511 -45928 -66139 -45896
rect -66511 -46172 -66447 -45928
rect -66203 -46172 -66139 -45928
rect -66511 -46204 -66139 -46172
rect -65511 -45928 -65139 -45896
rect -65511 -46172 -65447 -45928
rect -65203 -46172 -65139 -45928
rect -65511 -46204 -65139 -46172
rect -64511 -45928 -64139 -45896
rect -64511 -46172 -64447 -45928
rect -64203 -46172 -64139 -45928
rect -64511 -46204 -64139 -46172
rect -63511 -45928 -63139 -45896
rect -63511 -46172 -63447 -45928
rect -63203 -46172 -63139 -45928
rect -63511 -46204 -63139 -46172
rect -62511 -45928 -62139 -45896
rect -62511 -46172 -62447 -45928
rect -62203 -46172 -62139 -45928
rect -62511 -46204 -62139 -46172
rect -61511 -45928 -61139 -45896
rect -61511 -46172 -61447 -45928
rect -61203 -46172 -61139 -45928
rect -61511 -46204 -61139 -46172
rect -60511 -45928 -60139 -45896
rect -60511 -46172 -60447 -45928
rect -60203 -46172 -60139 -45928
rect -60511 -46204 -60139 -46172
rect -59511 -45928 -59139 -45896
rect -59511 -46172 -59447 -45928
rect -59203 -46172 -59139 -45928
rect -59511 -46204 -59139 -46172
rect -58511 -45928 -58139 -45896
rect -58511 -46172 -58447 -45928
rect -58203 -46172 -58139 -45928
rect -58511 -46204 -58139 -46172
rect -57511 -45928 -57139 -45896
rect -57511 -46172 -57447 -45928
rect -57203 -46172 -57139 -45928
rect -57511 -46204 -57139 -46172
rect -56511 -45928 -56139 -45896
rect -56511 -46172 -56447 -45928
rect -56203 -46172 -56139 -45928
rect -56511 -46204 -56139 -46172
rect -55511 -45928 -55139 -45896
rect -55511 -46172 -55447 -45928
rect -55203 -46172 -55139 -45928
rect -55511 -46204 -55139 -46172
rect -54511 -45928 -54139 -45896
rect -54511 -46172 -54447 -45928
rect -54203 -46172 -54139 -45928
rect -54511 -46204 -54139 -46172
rect -53511 -45928 -53139 -45896
rect -53511 -46172 -53447 -45928
rect -53203 -46172 -53139 -45928
rect -53511 -46204 -53139 -46172
rect -52511 -45928 -52139 -45896
rect -52511 -46172 -52447 -45928
rect -52203 -46172 -52139 -45928
rect -52511 -46204 -52139 -46172
rect -51511 -45928 -51139 -45896
rect -51511 -46172 -51447 -45928
rect -51203 -46172 -51139 -45928
rect -51511 -46204 -51139 -46172
rect -50511 -45928 -50139 -45896
rect -50511 -46172 -50447 -45928
rect -50203 -46172 -50139 -45928
rect -50511 -46204 -50139 -46172
rect -49511 -45928 -49139 -45896
rect -49511 -46172 -49447 -45928
rect -49203 -46172 -49139 -45928
rect -49511 -46204 -49139 -46172
rect -48831 -46204 -48825 -45896
rect -74825 -46210 -48825 -46204
rect 8275 -45896 34275 -45890
rect 8275 -46204 8281 -45896
rect 8589 -45928 8961 -45896
rect 8589 -46172 8653 -45928
rect 8897 -46172 8961 -45928
rect 8589 -46204 8961 -46172
rect 9589 -45928 9961 -45896
rect 9589 -46172 9653 -45928
rect 9897 -46172 9961 -45928
rect 9589 -46204 9961 -46172
rect 10589 -45928 10961 -45896
rect 10589 -46172 10653 -45928
rect 10897 -46172 10961 -45928
rect 10589 -46204 10961 -46172
rect 11589 -45928 11961 -45896
rect 11589 -46172 11653 -45928
rect 11897 -46172 11961 -45928
rect 11589 -46204 11961 -46172
rect 12589 -45928 12961 -45896
rect 12589 -46172 12653 -45928
rect 12897 -46172 12961 -45928
rect 12589 -46204 12961 -46172
rect 13589 -45928 13961 -45896
rect 13589 -46172 13653 -45928
rect 13897 -46172 13961 -45928
rect 13589 -46204 13961 -46172
rect 14589 -45928 14961 -45896
rect 14589 -46172 14653 -45928
rect 14897 -46172 14961 -45928
rect 14589 -46204 14961 -46172
rect 15589 -45928 15961 -45896
rect 15589 -46172 15653 -45928
rect 15897 -46172 15961 -45928
rect 15589 -46204 15961 -46172
rect 16589 -45928 16961 -45896
rect 16589 -46172 16653 -45928
rect 16897 -46172 16961 -45928
rect 16589 -46204 16961 -46172
rect 17589 -45928 17961 -45896
rect 17589 -46172 17653 -45928
rect 17897 -46172 17961 -45928
rect 17589 -46204 17961 -46172
rect 18589 -45928 18961 -45896
rect 18589 -46172 18653 -45928
rect 18897 -46172 18961 -45928
rect 18589 -46204 18961 -46172
rect 19589 -45928 19961 -45896
rect 19589 -46172 19653 -45928
rect 19897 -46172 19961 -45928
rect 19589 -46204 19961 -46172
rect 20589 -45928 20961 -45896
rect 20589 -46172 20653 -45928
rect 20897 -46172 20961 -45928
rect 20589 -46204 20961 -46172
rect 21589 -45928 21961 -45896
rect 21589 -46172 21653 -45928
rect 21897 -46172 21961 -45928
rect 21589 -46204 21961 -46172
rect 22589 -45928 22961 -45896
rect 22589 -46172 22653 -45928
rect 22897 -46172 22961 -45928
rect 22589 -46204 22961 -46172
rect 23589 -45928 23961 -45896
rect 23589 -46172 23653 -45928
rect 23897 -46172 23961 -45928
rect 23589 -46204 23961 -46172
rect 24589 -45928 24961 -45896
rect 24589 -46172 24653 -45928
rect 24897 -46172 24961 -45928
rect 24589 -46204 24961 -46172
rect 25589 -45928 25961 -45896
rect 25589 -46172 25653 -45928
rect 25897 -46172 25961 -45928
rect 25589 -46204 25961 -46172
rect 26589 -45928 26961 -45896
rect 26589 -46172 26653 -45928
rect 26897 -46172 26961 -45928
rect 26589 -46204 26961 -46172
rect 27589 -45928 27961 -45896
rect 27589 -46172 27653 -45928
rect 27897 -46172 27961 -45928
rect 27589 -46204 27961 -46172
rect 28589 -45928 28961 -45896
rect 28589 -46172 28653 -45928
rect 28897 -46172 28961 -45928
rect 28589 -46204 28961 -46172
rect 29589 -45928 29961 -45896
rect 29589 -46172 29653 -45928
rect 29897 -46172 29961 -45928
rect 29589 -46204 29961 -46172
rect 30589 -45928 30961 -45896
rect 30589 -46172 30653 -45928
rect 30897 -46172 30961 -45928
rect 30589 -46204 30961 -46172
rect 31589 -45928 31961 -45896
rect 31589 -46172 31653 -45928
rect 31897 -46172 31961 -45928
rect 31589 -46204 31961 -46172
rect 32589 -45928 32961 -45896
rect 32589 -46172 32653 -45928
rect 32897 -46172 32961 -45928
rect 32589 -46204 32961 -46172
rect 33589 -45928 33961 -45896
rect 33589 -46172 33653 -45928
rect 33897 -46172 33961 -45928
rect 33589 -46204 33961 -46172
rect 34269 -46204 34275 -45896
rect 8275 -46210 34275 -46204
rect -74485 -46236 -74165 -46210
rect -74485 -46544 -74479 -46236
rect -74171 -46544 -74165 -46236
rect -74485 -46550 -74165 -46544
rect -73485 -46236 -73165 -46210
rect -73485 -46544 -73479 -46236
rect -73171 -46544 -73165 -46236
rect -73485 -46550 -73165 -46544
rect -72485 -46236 -72165 -46210
rect -72485 -46544 -72479 -46236
rect -72171 -46544 -72165 -46236
rect -72485 -46550 -72165 -46544
rect -71485 -46236 -71165 -46210
rect -71485 -46544 -71479 -46236
rect -71171 -46544 -71165 -46236
rect -71485 -46550 -71165 -46544
rect -70485 -46236 -70165 -46210
rect -70485 -46544 -70479 -46236
rect -70171 -46544 -70165 -46236
rect -70485 -46550 -70165 -46544
rect -69485 -46236 -69165 -46210
rect -69485 -46544 -69479 -46236
rect -69171 -46544 -69165 -46236
rect -69485 -46550 -69165 -46544
rect -68485 -46236 -68165 -46210
rect -68485 -46544 -68479 -46236
rect -68171 -46544 -68165 -46236
rect -68485 -46550 -68165 -46544
rect -67485 -46236 -67165 -46210
rect -67485 -46544 -67479 -46236
rect -67171 -46544 -67165 -46236
rect -67485 -46550 -67165 -46544
rect -66485 -46236 -66165 -46210
rect -66485 -46544 -66479 -46236
rect -66171 -46544 -66165 -46236
rect -66485 -46550 -66165 -46544
rect -65485 -46236 -65165 -46210
rect -65485 -46544 -65479 -46236
rect -65171 -46544 -65165 -46236
rect -65485 -46550 -65165 -46544
rect -64485 -46236 -64165 -46210
rect -64485 -46544 -64479 -46236
rect -64171 -46544 -64165 -46236
rect -64485 -46550 -64165 -46544
rect -63485 -46236 -63165 -46210
rect -63485 -46544 -63479 -46236
rect -63171 -46544 -63165 -46236
rect -63485 -46550 -63165 -46544
rect -62485 -46236 -62165 -46210
rect -62485 -46544 -62479 -46236
rect -62171 -46544 -62165 -46236
rect -62485 -46550 -62165 -46544
rect -61485 -46236 -61165 -46210
rect -61485 -46544 -61479 -46236
rect -61171 -46544 -61165 -46236
rect -61485 -46550 -61165 -46544
rect -60485 -46236 -60165 -46210
rect -60485 -46544 -60479 -46236
rect -60171 -46544 -60165 -46236
rect -60485 -46550 -60165 -46544
rect -59485 -46236 -59165 -46210
rect -59485 -46544 -59479 -46236
rect -59171 -46544 -59165 -46236
rect -59485 -46550 -59165 -46544
rect -58485 -46236 -58165 -46210
rect -58485 -46544 -58479 -46236
rect -58171 -46544 -58165 -46236
rect -58485 -46550 -58165 -46544
rect -57485 -46236 -57165 -46210
rect -57485 -46544 -57479 -46236
rect -57171 -46544 -57165 -46236
rect -57485 -46550 -57165 -46544
rect -56485 -46236 -56165 -46210
rect -56485 -46544 -56479 -46236
rect -56171 -46544 -56165 -46236
rect -56485 -46550 -56165 -46544
rect -55485 -46236 -55165 -46210
rect -55485 -46544 -55479 -46236
rect -55171 -46544 -55165 -46236
rect -55485 -46550 -55165 -46544
rect -54485 -46236 -54165 -46210
rect -54485 -46544 -54479 -46236
rect -54171 -46544 -54165 -46236
rect -54485 -46550 -54165 -46544
rect -53485 -46236 -53165 -46210
rect -53485 -46544 -53479 -46236
rect -53171 -46544 -53165 -46236
rect -53485 -46550 -53165 -46544
rect -52485 -46236 -52165 -46210
rect -52485 -46544 -52479 -46236
rect -52171 -46544 -52165 -46236
rect -52485 -46550 -52165 -46544
rect -51485 -46236 -51165 -46210
rect -51485 -46544 -51479 -46236
rect -51171 -46544 -51165 -46236
rect -51485 -46550 -51165 -46544
rect -50485 -46236 -50165 -46210
rect -50485 -46544 -50479 -46236
rect -50171 -46544 -50165 -46236
rect -50485 -46550 -50165 -46544
rect -49485 -46236 -49165 -46210
rect -49485 -46544 -49479 -46236
rect -49171 -46544 -49165 -46236
rect -49485 -46550 -49165 -46544
rect 8615 -46236 8935 -46210
rect 8615 -46544 8621 -46236
rect 8929 -46544 8935 -46236
rect 8615 -46550 8935 -46544
rect 9615 -46236 9935 -46210
rect 9615 -46544 9621 -46236
rect 9929 -46544 9935 -46236
rect 9615 -46550 9935 -46544
rect 10615 -46236 10935 -46210
rect 10615 -46544 10621 -46236
rect 10929 -46544 10935 -46236
rect 10615 -46550 10935 -46544
rect 11615 -46236 11935 -46210
rect 11615 -46544 11621 -46236
rect 11929 -46544 11935 -46236
rect 11615 -46550 11935 -46544
rect 12615 -46236 12935 -46210
rect 12615 -46544 12621 -46236
rect 12929 -46544 12935 -46236
rect 12615 -46550 12935 -46544
rect 13615 -46236 13935 -46210
rect 13615 -46544 13621 -46236
rect 13929 -46544 13935 -46236
rect 13615 -46550 13935 -46544
rect 14615 -46236 14935 -46210
rect 14615 -46544 14621 -46236
rect 14929 -46544 14935 -46236
rect 14615 -46550 14935 -46544
rect 15615 -46236 15935 -46210
rect 15615 -46544 15621 -46236
rect 15929 -46544 15935 -46236
rect 15615 -46550 15935 -46544
rect 16615 -46236 16935 -46210
rect 16615 -46544 16621 -46236
rect 16929 -46544 16935 -46236
rect 16615 -46550 16935 -46544
rect 17615 -46236 17935 -46210
rect 17615 -46544 17621 -46236
rect 17929 -46544 17935 -46236
rect 17615 -46550 17935 -46544
rect 18615 -46236 18935 -46210
rect 18615 -46544 18621 -46236
rect 18929 -46544 18935 -46236
rect 18615 -46550 18935 -46544
rect 19615 -46236 19935 -46210
rect 19615 -46544 19621 -46236
rect 19929 -46544 19935 -46236
rect 19615 -46550 19935 -46544
rect 20615 -46236 20935 -46210
rect 20615 -46544 20621 -46236
rect 20929 -46544 20935 -46236
rect 20615 -46550 20935 -46544
rect 21615 -46236 21935 -46210
rect 21615 -46544 21621 -46236
rect 21929 -46544 21935 -46236
rect 21615 -46550 21935 -46544
rect 22615 -46236 22935 -46210
rect 22615 -46544 22621 -46236
rect 22929 -46544 22935 -46236
rect 22615 -46550 22935 -46544
rect 23615 -46236 23935 -46210
rect 23615 -46544 23621 -46236
rect 23929 -46544 23935 -46236
rect 23615 -46550 23935 -46544
rect 24615 -46236 24935 -46210
rect 24615 -46544 24621 -46236
rect 24929 -46544 24935 -46236
rect 24615 -46550 24935 -46544
rect 25615 -46236 25935 -46210
rect 25615 -46544 25621 -46236
rect 25929 -46544 25935 -46236
rect 25615 -46550 25935 -46544
rect 26615 -46236 26935 -46210
rect 26615 -46544 26621 -46236
rect 26929 -46544 26935 -46236
rect 26615 -46550 26935 -46544
rect 27615 -46236 27935 -46210
rect 27615 -46544 27621 -46236
rect 27929 -46544 27935 -46236
rect 27615 -46550 27935 -46544
rect 28615 -46236 28935 -46210
rect 28615 -46544 28621 -46236
rect 28929 -46544 28935 -46236
rect 28615 -46550 28935 -46544
rect 29615 -46236 29935 -46210
rect 29615 -46544 29621 -46236
rect 29929 -46544 29935 -46236
rect 29615 -46550 29935 -46544
rect 30615 -46236 30935 -46210
rect 30615 -46544 30621 -46236
rect 30929 -46544 30935 -46236
rect 30615 -46550 30935 -46544
rect 31615 -46236 31935 -46210
rect 31615 -46544 31621 -46236
rect 31929 -46544 31935 -46236
rect 31615 -46550 31935 -46544
rect 32615 -46236 32935 -46210
rect 32615 -46544 32621 -46236
rect 32929 -46544 32935 -46236
rect 32615 -46550 32935 -46544
rect 33615 -46236 33935 -46210
rect 33615 -46544 33621 -46236
rect 33929 -46544 33935 -46236
rect 33615 -46550 33935 -46544
<< via1 >>
rect -74479 38236 -74171 38544
rect -73479 38236 -73171 38544
rect -72479 38236 -72171 38544
rect -71479 38236 -71171 38544
rect -70479 38236 -70171 38544
rect -69479 38236 -69171 38544
rect -68479 38236 -68171 38544
rect -67479 38236 -67171 38544
rect -66479 38236 -66171 38544
rect -65479 38236 -65171 38544
rect -64479 38236 -64171 38544
rect -63479 38236 -63171 38544
rect -62479 38236 -62171 38544
rect -61479 38236 -61171 38544
rect -60479 38236 -60171 38544
rect -59479 38236 -59171 38544
rect 10000 38236 10308 38544
rect 11000 38236 11308 38544
rect 12000 38236 12308 38544
rect 13000 38236 13308 38544
rect 14000 38236 14308 38544
rect 15000 38236 15308 38544
rect 16000 38236 16308 38544
rect 17000 38236 17308 38544
rect 18000 38236 18308 38544
rect 19000 38236 19308 38544
rect 20000 38236 20308 38544
rect 21000 38236 21308 38544
rect 22000 38236 22308 38544
rect 23000 38236 23308 38544
rect 24000 38236 24308 38544
rect 25000 38236 25308 38544
rect 26000 38236 26308 38544
rect 27000 38236 27308 38544
rect 28000 38236 28308 38544
rect 29000 38236 29308 38544
rect 30000 38236 30308 38544
rect 31000 38236 31308 38544
rect 32000 38236 32308 38544
rect 33000 38236 33308 38544
rect 34000 38236 34308 38544
rect -74819 37896 -74511 38204
rect -74447 37928 -74203 38172
rect -74139 37896 -73511 38204
rect -73447 37928 -73203 38172
rect -73139 37896 -72511 38204
rect -72447 37928 -72203 38172
rect -72139 37896 -71511 38204
rect -71447 37928 -71203 38172
rect -71139 37896 -70511 38204
rect -70447 37928 -70203 38172
rect -70139 37896 -69511 38204
rect -69447 37928 -69203 38172
rect -69139 37896 -68511 38204
rect -68447 37928 -68203 38172
rect -68139 37896 -67511 38204
rect -67447 37928 -67203 38172
rect -67139 37896 -66511 38204
rect -66447 37928 -66203 38172
rect -66139 37896 -65511 38204
rect -65447 37928 -65203 38172
rect -65139 37896 -64511 38204
rect -64447 37928 -64203 38172
rect -64139 37896 -63511 38204
rect -63447 37928 -63203 38172
rect -63139 37896 -62511 38204
rect -62447 37928 -62203 38172
rect -62139 37896 -61511 38204
rect -61447 37928 -61203 38172
rect -61139 37896 -60511 38204
rect -60447 37928 -60203 38172
rect -60139 37896 -59511 38204
rect -59447 37928 -59203 38172
rect -59139 37896 -58831 38204
rect 9660 37896 9968 38204
rect 10032 37928 10276 38172
rect 10340 37896 10968 38204
rect 11032 37928 11276 38172
rect 11340 37896 11968 38204
rect 12032 37928 12276 38172
rect 12340 37896 12968 38204
rect 13032 37928 13276 38172
rect 13340 37896 13968 38204
rect 14032 37928 14276 38172
rect 14340 37896 14968 38204
rect 15032 37928 15276 38172
rect 15340 37896 15968 38204
rect 16032 37928 16276 38172
rect 16340 37896 16968 38204
rect 17032 37928 17276 38172
rect 17340 37896 17968 38204
rect 18032 37928 18276 38172
rect 18340 37896 18968 38204
rect 19032 37928 19276 38172
rect 19340 37896 19968 38204
rect 20032 37928 20276 38172
rect 20340 37896 20968 38204
rect 21032 37928 21276 38172
rect 21340 37896 21968 38204
rect 22032 37928 22276 38172
rect 22340 37896 22968 38204
rect 23032 37928 23276 38172
rect 23340 37896 23968 38204
rect 24032 37928 24276 38172
rect 24340 37896 24968 38204
rect 25032 37928 25276 38172
rect 25340 37896 25968 38204
rect 26032 37928 26276 38172
rect 26340 37896 26968 38204
rect 27032 37928 27276 38172
rect 27340 37896 27968 38204
rect 28032 37928 28276 38172
rect 28340 37896 28968 38204
rect 29032 37928 29276 38172
rect 29340 37896 29968 38204
rect 30032 37928 30276 38172
rect 30340 37896 30968 38204
rect 31032 37928 31276 38172
rect 31340 37896 31968 38204
rect 32032 37928 32276 38172
rect 32340 37896 32968 38204
rect 33032 37928 33276 38172
rect 33340 37896 33968 38204
rect 34032 37928 34276 38172
rect 34340 37896 34648 38204
rect -74479 37236 -74171 37864
rect -73479 37236 -73171 37864
rect -72479 37236 -72171 37864
rect -71479 37236 -71171 37864
rect -70479 37236 -70171 37864
rect -69479 37236 -69171 37864
rect -68479 37236 -68171 37864
rect -67479 37236 -67171 37864
rect -66479 37236 -66171 37864
rect -65479 37236 -65171 37864
rect -64479 37236 -64171 37864
rect -63479 37236 -63171 37864
rect -62479 37236 -62171 37864
rect -61479 37236 -61171 37864
rect -60479 37236 -60171 37864
rect -59479 37236 -59171 37864
rect 10000 37236 10308 37864
rect 11000 37236 11308 37864
rect 12000 37236 12308 37864
rect 13000 37236 13308 37864
rect 14000 37236 14308 37864
rect 15000 37236 15308 37864
rect 16000 37236 16308 37864
rect 17000 37236 17308 37864
rect 18000 37236 18308 37864
rect 19000 37236 19308 37864
rect 20000 37236 20308 37864
rect 21000 37236 21308 37864
rect 22000 37236 22308 37864
rect 23000 37236 23308 37864
rect 24000 37236 24308 37864
rect 25000 37236 25308 37864
rect 26000 37236 26308 37864
rect 27000 37236 27308 37864
rect 28000 37236 28308 37864
rect 29000 37236 29308 37864
rect 30000 37236 30308 37864
rect 31000 37236 31308 37864
rect 32000 37236 32308 37864
rect 33000 37236 33308 37864
rect 34000 37236 34308 37864
rect -74819 36896 -74511 37204
rect -74447 36928 -74203 37172
rect -74139 36896 -73511 37204
rect -73447 36928 -73203 37172
rect -73139 36896 -72511 37204
rect -72447 36928 -72203 37172
rect -72139 36896 -71511 37204
rect -71447 36928 -71203 37172
rect -71139 36896 -70511 37204
rect -70447 36928 -70203 37172
rect -70139 36896 -69511 37204
rect -69447 36928 -69203 37172
rect -69139 36896 -68511 37204
rect -68447 36928 -68203 37172
rect -68139 36896 -67511 37204
rect -67447 36928 -67203 37172
rect -67139 36896 -66511 37204
rect -66447 36928 -66203 37172
rect -66139 36896 -65511 37204
rect -65447 36928 -65203 37172
rect -65139 36896 -64511 37204
rect -64447 36928 -64203 37172
rect -64139 36896 -63511 37204
rect -63447 36928 -63203 37172
rect -63139 36896 -62511 37204
rect -62447 36928 -62203 37172
rect -62139 36896 -61511 37204
rect -61447 36928 -61203 37172
rect -61139 36896 -60511 37204
rect -60447 36928 -60203 37172
rect -60139 36896 -59511 37204
rect -59447 36928 -59203 37172
rect -59139 36896 -58831 37204
rect 9660 36896 9968 37204
rect 10032 36928 10276 37172
rect 10340 36896 10968 37204
rect 11032 36928 11276 37172
rect 11340 36896 11968 37204
rect 12032 36928 12276 37172
rect 12340 36896 12968 37204
rect 13032 36928 13276 37172
rect 13340 36896 13968 37204
rect 14032 36928 14276 37172
rect 14340 36896 14968 37204
rect 15032 36928 15276 37172
rect 15340 36896 15968 37204
rect 16032 36928 16276 37172
rect 16340 36896 16968 37204
rect 17032 36928 17276 37172
rect 17340 36896 17968 37204
rect 18032 36928 18276 37172
rect 18340 36896 18968 37204
rect 19032 36928 19276 37172
rect 19340 36896 19968 37204
rect 20032 36928 20276 37172
rect 20340 36896 20968 37204
rect 21032 36928 21276 37172
rect 21340 36896 21968 37204
rect 22032 36928 22276 37172
rect 22340 36896 22968 37204
rect 23032 36928 23276 37172
rect 23340 36896 23968 37204
rect 24032 36928 24276 37172
rect 24340 36896 24968 37204
rect 25032 36928 25276 37172
rect 25340 36896 25968 37204
rect 26032 36928 26276 37172
rect 26340 36896 26968 37204
rect 27032 36928 27276 37172
rect 27340 36896 27968 37204
rect 28032 36928 28276 37172
rect 28340 36896 28968 37204
rect 29032 36928 29276 37172
rect 29340 36896 29968 37204
rect 30032 36928 30276 37172
rect 30340 36896 30968 37204
rect 31032 36928 31276 37172
rect 31340 36896 31968 37204
rect 32032 36928 32276 37172
rect 32340 36896 32968 37204
rect 33032 36928 33276 37172
rect 33340 36896 33968 37204
rect 34032 36928 34276 37172
rect 34340 36896 34648 37204
rect -74479 36236 -74171 36864
rect -73479 36236 -73171 36864
rect -72479 36236 -72171 36864
rect -71479 36236 -71171 36864
rect -70479 36236 -70171 36864
rect -69479 36236 -69171 36864
rect -68479 36236 -68171 36864
rect -67479 36236 -67171 36864
rect -66479 36236 -66171 36864
rect -65479 36236 -65171 36864
rect -64479 36236 -64171 36864
rect -63479 36236 -63171 36864
rect -62479 36236 -62171 36864
rect -61479 36236 -61171 36864
rect -60479 36236 -60171 36864
rect -59479 36236 -59171 36864
rect 10000 36236 10308 36864
rect 11000 36236 11308 36864
rect 12000 36236 12308 36864
rect 13000 36236 13308 36864
rect 14000 36236 14308 36864
rect 15000 36236 15308 36864
rect 16000 36236 16308 36864
rect 17000 36236 17308 36864
rect 18000 36236 18308 36864
rect 19000 36236 19308 36864
rect 20000 36236 20308 36864
rect 21000 36236 21308 36864
rect 22000 36236 22308 36864
rect 23000 36236 23308 36864
rect 24000 36236 24308 36864
rect 25000 36236 25308 36864
rect 26000 36236 26308 36864
rect 27000 36236 27308 36864
rect 28000 36236 28308 36864
rect 29000 36236 29308 36864
rect 30000 36236 30308 36864
rect 31000 36236 31308 36864
rect 32000 36236 32308 36864
rect 33000 36236 33308 36864
rect 34000 36236 34308 36864
rect -74819 35896 -74511 36204
rect -74447 35928 -74203 36172
rect -74139 35896 -73511 36204
rect -73447 35928 -73203 36172
rect -73139 35896 -72511 36204
rect -72447 35928 -72203 36172
rect -72139 35896 -71511 36204
rect -71447 35928 -71203 36172
rect -71139 35896 -70511 36204
rect -70447 35928 -70203 36172
rect -70139 35896 -69511 36204
rect -69447 35928 -69203 36172
rect -69139 35896 -68511 36204
rect -68447 35928 -68203 36172
rect -68139 35896 -67511 36204
rect -67447 35928 -67203 36172
rect -67139 35896 -66511 36204
rect -66447 35928 -66203 36172
rect -66139 35896 -65511 36204
rect -65447 35928 -65203 36172
rect -65139 35896 -64511 36204
rect -64447 35928 -64203 36172
rect -64139 35896 -63511 36204
rect -63447 35928 -63203 36172
rect -63139 35896 -62511 36204
rect -62447 35928 -62203 36172
rect -62139 35896 -61511 36204
rect -61447 35928 -61203 36172
rect -61139 35896 -60511 36204
rect -60447 35928 -60203 36172
rect -60139 35896 -59511 36204
rect -59447 35928 -59203 36172
rect -59139 35896 -58831 36204
rect 9660 35896 9968 36204
rect 10032 35928 10276 36172
rect 10340 35896 10968 36204
rect 11032 35928 11276 36172
rect 11340 35896 11968 36204
rect 12032 35928 12276 36172
rect 12340 35896 12968 36204
rect 13032 35928 13276 36172
rect 13340 35896 13968 36204
rect 14032 35928 14276 36172
rect 14340 35896 14968 36204
rect 15032 35928 15276 36172
rect 15340 35896 15968 36204
rect 16032 35928 16276 36172
rect 16340 35896 16968 36204
rect 17032 35928 17276 36172
rect 17340 35896 17968 36204
rect 18032 35928 18276 36172
rect 18340 35896 18968 36204
rect 19032 35928 19276 36172
rect 19340 35896 19968 36204
rect 20032 35928 20276 36172
rect 20340 35896 20968 36204
rect 21032 35928 21276 36172
rect 21340 35896 21968 36204
rect 22032 35928 22276 36172
rect 22340 35896 22968 36204
rect 23032 35928 23276 36172
rect 23340 35896 23968 36204
rect 24032 35928 24276 36172
rect 24340 35896 24968 36204
rect 25032 35928 25276 36172
rect 25340 35896 25968 36204
rect 26032 35928 26276 36172
rect 26340 35896 26968 36204
rect 27032 35928 27276 36172
rect 27340 35896 27968 36204
rect 28032 35928 28276 36172
rect 28340 35896 28968 36204
rect 29032 35928 29276 36172
rect 29340 35896 29968 36204
rect 30032 35928 30276 36172
rect 30340 35896 30968 36204
rect 31032 35928 31276 36172
rect 31340 35896 31968 36204
rect 32032 35928 32276 36172
rect 32340 35896 32968 36204
rect 33032 35928 33276 36172
rect 33340 35896 33968 36204
rect 34032 35928 34276 36172
rect 34340 35896 34648 36204
rect -74479 35236 -74171 35864
rect -73479 35236 -73171 35864
rect -72479 35236 -72171 35864
rect -71479 35236 -71171 35864
rect -70479 35236 -70171 35864
rect -69479 35236 -69171 35864
rect -68479 35236 -68171 35864
rect -67479 35236 -67171 35864
rect -66479 35236 -66171 35864
rect -65479 35236 -65171 35864
rect -64479 35236 -64171 35864
rect -63479 35236 -63171 35864
rect -62479 35236 -62171 35864
rect -61479 35236 -61171 35864
rect -60479 35236 -60171 35864
rect -59479 35236 -59171 35864
rect 10000 35236 10308 35864
rect 11000 35236 11308 35864
rect 12000 35236 12308 35864
rect 13000 35236 13308 35864
rect 14000 35236 14308 35864
rect 15000 35236 15308 35864
rect 16000 35236 16308 35864
rect 17000 35236 17308 35864
rect 18000 35236 18308 35864
rect 19000 35236 19308 35864
rect 20000 35236 20308 35864
rect 21000 35236 21308 35864
rect 22000 35236 22308 35864
rect 23000 35236 23308 35864
rect 24000 35236 24308 35864
rect 25000 35236 25308 35864
rect 26000 35236 26308 35864
rect 27000 35236 27308 35864
rect 28000 35236 28308 35864
rect 29000 35236 29308 35864
rect 30000 35236 30308 35864
rect 31000 35236 31308 35864
rect 32000 35236 32308 35864
rect 33000 35236 33308 35864
rect 34000 35236 34308 35864
rect -74819 34896 -74511 35204
rect -74447 34928 -74203 35172
rect -74139 34896 -73511 35204
rect -73447 34928 -73203 35172
rect -73139 34896 -72511 35204
rect -72447 34928 -72203 35172
rect -72139 34896 -71511 35204
rect -71447 34928 -71203 35172
rect -71139 34896 -70511 35204
rect -70447 34928 -70203 35172
rect -70139 34896 -69511 35204
rect -69447 34928 -69203 35172
rect -69139 34896 -68511 35204
rect -68447 34928 -68203 35172
rect -68139 34896 -67511 35204
rect -67447 34928 -67203 35172
rect -67139 34896 -66511 35204
rect -66447 34928 -66203 35172
rect -66139 34896 -65511 35204
rect -65447 34928 -65203 35172
rect -65139 34896 -64511 35204
rect -64447 34928 -64203 35172
rect -64139 34896 -63511 35204
rect -63447 34928 -63203 35172
rect -63139 34896 -62511 35204
rect -62447 34928 -62203 35172
rect -62139 34896 -61511 35204
rect -61447 34928 -61203 35172
rect -61139 34896 -60511 35204
rect -60447 34928 -60203 35172
rect -60139 34896 -59511 35204
rect -59447 34928 -59203 35172
rect -59139 34896 -58831 35204
rect 9660 34896 9968 35204
rect 10032 34928 10276 35172
rect 10340 34896 10968 35204
rect 11032 34928 11276 35172
rect 11340 34896 11968 35204
rect 12032 34928 12276 35172
rect 12340 34896 12968 35204
rect 13032 34928 13276 35172
rect 13340 34896 13968 35204
rect 14032 34928 14276 35172
rect 14340 34896 14968 35204
rect 15032 34928 15276 35172
rect 15340 34896 15968 35204
rect 16032 34928 16276 35172
rect 16340 34896 16968 35204
rect 17032 34928 17276 35172
rect 17340 34896 17968 35204
rect 18032 34928 18276 35172
rect 18340 34896 18968 35204
rect 19032 34928 19276 35172
rect 19340 34896 19968 35204
rect 20032 34928 20276 35172
rect 20340 34896 20968 35204
rect 21032 34928 21276 35172
rect 21340 34896 21968 35204
rect 22032 34928 22276 35172
rect 22340 34896 22968 35204
rect 23032 34928 23276 35172
rect 23340 34896 23968 35204
rect 24032 34928 24276 35172
rect 24340 34896 24968 35204
rect 25032 34928 25276 35172
rect 25340 34896 25968 35204
rect 26032 34928 26276 35172
rect 26340 34896 26968 35204
rect 27032 34928 27276 35172
rect 27340 34896 27968 35204
rect 28032 34928 28276 35172
rect 28340 34896 28968 35204
rect 29032 34928 29276 35172
rect 29340 34896 29968 35204
rect 30032 34928 30276 35172
rect 30340 34896 30968 35204
rect 31032 34928 31276 35172
rect 31340 34896 31968 35204
rect 32032 34928 32276 35172
rect 32340 34896 32968 35204
rect 33032 34928 33276 35172
rect 33340 34896 33968 35204
rect 34032 34928 34276 35172
rect 34340 34896 34648 35204
rect -74479 34236 -74171 34864
rect -73479 34236 -73171 34864
rect -72479 34236 -72171 34864
rect -71479 34236 -71171 34864
rect -70479 34236 -70171 34864
rect -69479 34236 -69171 34864
rect -68479 34236 -68171 34864
rect -67479 34236 -67171 34864
rect -66479 34236 -66171 34864
rect -65479 34236 -65171 34864
rect -64479 34236 -64171 34864
rect -63479 34236 -63171 34864
rect -62479 34236 -62171 34864
rect -61479 34236 -61171 34864
rect -60479 34236 -60171 34864
rect -59479 34236 -59171 34864
rect 10000 34236 10308 34864
rect 11000 34236 11308 34864
rect 12000 34236 12308 34864
rect 13000 34236 13308 34864
rect 14000 34236 14308 34864
rect 15000 34236 15308 34864
rect 16000 34236 16308 34864
rect 17000 34236 17308 34864
rect 18000 34236 18308 34864
rect 19000 34236 19308 34864
rect 20000 34236 20308 34864
rect 21000 34236 21308 34864
rect 22000 34236 22308 34864
rect 23000 34236 23308 34864
rect 24000 34236 24308 34864
rect 25000 34236 25308 34864
rect 26000 34236 26308 34864
rect 27000 34236 27308 34864
rect 28000 34236 28308 34864
rect 29000 34236 29308 34864
rect 30000 34236 30308 34864
rect 31000 34236 31308 34864
rect 32000 34236 32308 34864
rect 33000 34236 33308 34864
rect 34000 34236 34308 34864
rect -74819 33896 -74511 34204
rect -74447 33928 -74203 34172
rect -74139 33896 -73511 34204
rect -73447 33928 -73203 34172
rect -73139 33896 -72511 34204
rect -72447 33928 -72203 34172
rect -72139 33896 -71511 34204
rect -71447 33928 -71203 34172
rect -71139 33896 -70511 34204
rect -70447 33928 -70203 34172
rect -70139 33896 -69511 34204
rect -69447 33928 -69203 34172
rect -69139 33896 -68511 34204
rect -68447 33928 -68203 34172
rect -68139 33896 -67511 34204
rect -67447 33928 -67203 34172
rect -67139 33896 -66511 34204
rect -66447 33928 -66203 34172
rect -66139 33896 -65511 34204
rect -65447 33928 -65203 34172
rect -65139 33896 -64511 34204
rect -64447 33928 -64203 34172
rect -64139 33896 -63511 34204
rect -63447 33928 -63203 34172
rect -63139 33896 -62511 34204
rect -62447 33928 -62203 34172
rect -62139 33896 -61511 34204
rect -61447 33928 -61203 34172
rect -61139 33896 -60511 34204
rect -60447 33928 -60203 34172
rect -60139 33896 -59511 34204
rect -59447 33928 -59203 34172
rect -59139 33896 -58831 34204
rect -74479 33236 -74171 33864
rect -73479 33236 -73171 33864
rect -72479 33236 -72171 33864
rect -71479 33236 -71171 33864
rect -70479 33236 -70171 33864
rect -69479 33236 -69171 33864
rect -68479 33236 -68171 33864
rect -67479 33236 -67171 33864
rect -66479 33236 -66171 33864
rect -65479 33236 -65171 33864
rect -64479 33236 -64171 33864
rect -63479 33236 -63171 33864
rect -62479 33236 -62171 33864
rect -61479 33236 -61171 33864
rect -60479 33236 -60171 33864
rect -59479 33236 -59171 33864
rect -50466 33542 -48814 34170
rect 2881 33542 4533 34170
rect 9660 33896 9968 34204
rect 10032 33928 10276 34172
rect 10340 33896 10968 34204
rect 11032 33928 11276 34172
rect 11340 33896 11968 34204
rect 12032 33928 12276 34172
rect 12340 33896 12968 34204
rect 13032 33928 13276 34172
rect 13340 33896 13968 34204
rect 14032 33928 14276 34172
rect 14340 33896 14968 34204
rect 15032 33928 15276 34172
rect 15340 33896 15968 34204
rect 16032 33928 16276 34172
rect 16340 33896 16968 34204
rect 17032 33928 17276 34172
rect 17340 33896 17968 34204
rect 18032 33928 18276 34172
rect 18340 33896 18968 34204
rect 19032 33928 19276 34172
rect 19340 33896 19968 34204
rect 20032 33928 20276 34172
rect 20340 33896 20968 34204
rect 21032 33928 21276 34172
rect 21340 33896 21968 34204
rect 22032 33928 22276 34172
rect 22340 33896 22968 34204
rect 23032 33928 23276 34172
rect 23340 33896 23968 34204
rect 24032 33928 24276 34172
rect 24340 33896 24968 34204
rect 25032 33928 25276 34172
rect 25340 33896 25968 34204
rect 26032 33928 26276 34172
rect 26340 33896 26968 34204
rect 27032 33928 27276 34172
rect 27340 33896 27968 34204
rect 28032 33928 28276 34172
rect 28340 33896 28968 34204
rect 29032 33928 29276 34172
rect 29340 33896 29968 34204
rect 30032 33928 30276 34172
rect 30340 33896 30968 34204
rect 31032 33928 31276 34172
rect 31340 33896 31968 34204
rect 32032 33928 32276 34172
rect 32340 33896 32968 34204
rect 33032 33928 33276 34172
rect 33340 33896 33968 34204
rect 34032 33928 34276 34172
rect 34340 33896 34648 34204
rect -74819 32896 -74511 33204
rect -74447 32928 -74203 33172
rect -74139 32896 -73511 33204
rect -73447 32928 -73203 33172
rect -73139 32896 -72511 33204
rect -72447 32928 -72203 33172
rect -72139 32896 -71511 33204
rect -71447 32928 -71203 33172
rect -71139 32896 -70511 33204
rect -70447 32928 -70203 33172
rect -70139 32896 -69511 33204
rect -69447 32928 -69203 33172
rect -69139 32896 -68511 33204
rect -68447 32928 -68203 33172
rect -68139 32896 -67511 33204
rect -67447 32928 -67203 33172
rect -67139 32896 -66511 33204
rect -66447 32928 -66203 33172
rect -66139 32896 -65511 33204
rect -65447 32928 -65203 33172
rect -65139 32896 -64511 33204
rect -64447 32928 -64203 33172
rect -64139 32896 -63511 33204
rect -63447 32928 -63203 33172
rect -63139 32896 -62511 33204
rect -62447 32928 -62203 33172
rect -62139 32896 -61511 33204
rect -61447 32928 -61203 33172
rect -61139 32896 -60511 33204
rect -60447 32928 -60203 33172
rect -60139 32896 -59511 33204
rect -59447 32928 -59203 33172
rect -59139 32896 -58831 33204
rect -74479 32236 -74171 32864
rect -73479 32236 -73171 32864
rect -72479 32236 -72171 32864
rect -71479 32236 -71171 32864
rect -70479 32236 -70171 32864
rect -69479 32236 -69171 32864
rect -68479 32236 -68171 32864
rect -67479 32236 -67171 32864
rect -66479 32236 -66171 32864
rect -65479 32236 -65171 32864
rect -64479 32236 -64171 32864
rect -63479 32236 -63171 32864
rect -62479 32236 -62171 32864
rect -61479 32236 -61171 32864
rect -60479 32236 -60171 32864
rect -59479 32236 -59171 32864
rect -50951 32940 -50579 32965
rect -50951 32618 -50926 32940
rect -50926 32618 -50604 32940
rect -50604 32618 -50579 32940
rect -50951 32593 -50579 32618
rect -50298 33273 -50246 33298
rect -50298 33246 -50289 33273
rect -50289 33246 -50255 33273
rect -50255 33246 -50246 33273
rect -50298 33201 -50246 33234
rect -50298 33182 -50289 33201
rect -50289 33182 -50255 33201
rect -50255 33182 -50246 33201
rect -50298 33167 -50289 33170
rect -50289 33167 -50255 33170
rect -50255 33167 -50246 33170
rect -50298 33129 -50246 33167
rect -50298 33118 -50289 33129
rect -50289 33118 -50255 33129
rect -50255 33118 -50246 33129
rect -50298 33095 -50289 33106
rect -50289 33095 -50255 33106
rect -50255 33095 -50246 33106
rect -50298 33057 -50246 33095
rect -50298 33054 -50289 33057
rect -50289 33054 -50255 33057
rect -50255 33054 -50246 33057
rect -50298 33023 -50289 33042
rect -50289 33023 -50255 33042
rect -50255 33023 -50246 33042
rect -50298 32990 -50246 33023
rect -50298 32951 -50289 32978
rect -50289 32951 -50255 32978
rect -50255 32951 -50246 32978
rect -50298 32926 -50246 32951
rect -49982 33273 -49930 33298
rect -49982 33246 -49973 33273
rect -49973 33246 -49939 33273
rect -49939 33246 -49930 33273
rect -49982 33201 -49930 33234
rect -49982 33182 -49973 33201
rect -49973 33182 -49939 33201
rect -49939 33182 -49930 33201
rect -49982 33167 -49973 33170
rect -49973 33167 -49939 33170
rect -49939 33167 -49930 33170
rect -49982 33129 -49930 33167
rect -49982 33118 -49973 33129
rect -49973 33118 -49939 33129
rect -49939 33118 -49930 33129
rect -49982 33095 -49973 33106
rect -49973 33095 -49939 33106
rect -49939 33095 -49930 33106
rect -49982 33057 -49930 33095
rect -49982 33054 -49973 33057
rect -49973 33054 -49939 33057
rect -49939 33054 -49930 33057
rect -49982 33023 -49973 33042
rect -49973 33023 -49939 33042
rect -49939 33023 -49930 33042
rect -49982 32990 -49930 33023
rect -49982 32951 -49973 32978
rect -49973 32951 -49939 32978
rect -49939 32951 -49930 32978
rect -49982 32926 -49930 32951
rect -49666 33273 -49614 33298
rect -49666 33246 -49657 33273
rect -49657 33246 -49623 33273
rect -49623 33246 -49614 33273
rect -49666 33201 -49614 33234
rect -49666 33182 -49657 33201
rect -49657 33182 -49623 33201
rect -49623 33182 -49614 33201
rect -49666 33167 -49657 33170
rect -49657 33167 -49623 33170
rect -49623 33167 -49614 33170
rect -49666 33129 -49614 33167
rect -49666 33118 -49657 33129
rect -49657 33118 -49623 33129
rect -49623 33118 -49614 33129
rect -49666 33095 -49657 33106
rect -49657 33095 -49623 33106
rect -49623 33095 -49614 33106
rect -49666 33057 -49614 33095
rect -49666 33054 -49657 33057
rect -49657 33054 -49623 33057
rect -49623 33054 -49614 33057
rect -49666 33023 -49657 33042
rect -49657 33023 -49623 33042
rect -49623 33023 -49614 33042
rect -49666 32990 -49614 33023
rect -49666 32951 -49657 32978
rect -49657 32951 -49623 32978
rect -49623 32951 -49614 32978
rect -49666 32926 -49614 32951
rect -49350 33273 -49298 33298
rect -49350 33246 -49341 33273
rect -49341 33246 -49307 33273
rect -49307 33246 -49298 33273
rect -49350 33201 -49298 33234
rect -49350 33182 -49341 33201
rect -49341 33182 -49307 33201
rect -49307 33182 -49298 33201
rect -49350 33167 -49341 33170
rect -49341 33167 -49307 33170
rect -49307 33167 -49298 33170
rect -49350 33129 -49298 33167
rect -49350 33118 -49341 33129
rect -49341 33118 -49307 33129
rect -49307 33118 -49298 33129
rect -49350 33095 -49341 33106
rect -49341 33095 -49307 33106
rect -49307 33095 -49298 33106
rect -49350 33057 -49298 33095
rect -49350 33054 -49341 33057
rect -49341 33054 -49307 33057
rect -49307 33054 -49298 33057
rect -49350 33023 -49341 33042
rect -49341 33023 -49307 33042
rect -49307 33023 -49298 33042
rect -49350 32990 -49298 33023
rect -49350 32951 -49341 32978
rect -49341 32951 -49307 32978
rect -49307 32951 -49298 32978
rect -49350 32926 -49298 32951
rect -49034 33273 -48982 33298
rect -49034 33246 -49025 33273
rect -49025 33246 -48991 33273
rect -48991 33246 -48982 33273
rect -49034 33201 -48982 33234
rect -49034 33182 -49025 33201
rect -49025 33182 -48991 33201
rect -48991 33182 -48982 33201
rect -49034 33167 -49025 33170
rect -49025 33167 -48991 33170
rect -48991 33167 -48982 33170
rect -49034 33129 -48982 33167
rect -49034 33118 -49025 33129
rect -49025 33118 -48991 33129
rect -48991 33118 -48982 33129
rect -49034 33095 -49025 33106
rect -49025 33095 -48991 33106
rect -48991 33095 -48982 33106
rect -49034 33057 -48982 33095
rect -49034 33054 -49025 33057
rect -49025 33054 -48991 33057
rect -48991 33054 -48982 33057
rect -49034 33023 -49025 33042
rect -49025 33023 -48991 33042
rect -48991 33023 -48982 33042
rect -49034 32990 -48982 33023
rect -49034 32951 -49025 32978
rect -49025 32951 -48991 32978
rect -48991 32951 -48982 32978
rect -49034 32926 -48982 32951
rect 2396 32940 2768 32965
rect -74819 31896 -74511 32204
rect -74447 31928 -74203 32172
rect -74139 31896 -73511 32204
rect -73447 31928 -73203 32172
rect -73139 31896 -72511 32204
rect -72447 31928 -72203 32172
rect -72139 31896 -71511 32204
rect -71447 31928 -71203 32172
rect -71139 31896 -70511 32204
rect -70447 31928 -70203 32172
rect -70139 31896 -69511 32204
rect -69447 31928 -69203 32172
rect -69139 31896 -68511 32204
rect -68447 31928 -68203 32172
rect -68139 31896 -67511 32204
rect -67447 31928 -67203 32172
rect -67139 31896 -66511 32204
rect -66447 31928 -66203 32172
rect -66139 31896 -65511 32204
rect -65447 31928 -65203 32172
rect -65139 31896 -64511 32204
rect -64447 31928 -64203 32172
rect -64139 31896 -63511 32204
rect -63447 31928 -63203 32172
rect -63139 31896 -62511 32204
rect -62447 31928 -62203 32172
rect -62139 31896 -61511 32204
rect -61447 31928 -61203 32172
rect -61139 31896 -60511 32204
rect -60447 31928 -60203 32172
rect -60139 31896 -59511 32204
rect -59447 31928 -59203 32172
rect -59139 31896 -58831 32204
rect -50298 32608 -50246 32645
rect -50298 32593 -50289 32608
rect -50289 32593 -50255 32608
rect -50255 32593 -50246 32608
rect -50298 32574 -50289 32581
rect -50289 32574 -50255 32581
rect -50255 32574 -50246 32581
rect -50298 32536 -50246 32574
rect -50298 32529 -50289 32536
rect -50289 32529 -50255 32536
rect -50255 32529 -50246 32536
rect -50298 32502 -50289 32517
rect -50289 32502 -50255 32517
rect -50255 32502 -50246 32517
rect -50298 32465 -50246 32502
rect -49982 32608 -49930 32645
rect -49982 32593 -49973 32608
rect -49973 32593 -49939 32608
rect -49939 32593 -49930 32608
rect -49982 32574 -49973 32581
rect -49973 32574 -49939 32581
rect -49939 32574 -49930 32581
rect -49982 32536 -49930 32574
rect -49982 32529 -49973 32536
rect -49973 32529 -49939 32536
rect -49939 32529 -49930 32536
rect -49982 32502 -49973 32517
rect -49973 32502 -49939 32517
rect -49939 32502 -49930 32517
rect -49982 32465 -49930 32502
rect -49666 32608 -49614 32645
rect -49666 32593 -49657 32608
rect -49657 32593 -49623 32608
rect -49623 32593 -49614 32608
rect -49666 32574 -49657 32581
rect -49657 32574 -49623 32581
rect -49623 32574 -49614 32581
rect -49666 32536 -49614 32574
rect -49666 32529 -49657 32536
rect -49657 32529 -49623 32536
rect -49623 32529 -49614 32536
rect -49666 32502 -49657 32517
rect -49657 32502 -49623 32517
rect -49623 32502 -49614 32517
rect -49666 32465 -49614 32502
rect -49350 32608 -49298 32645
rect -49350 32593 -49341 32608
rect -49341 32593 -49307 32608
rect -49307 32593 -49298 32608
rect -49350 32574 -49341 32581
rect -49341 32574 -49307 32581
rect -49307 32574 -49298 32581
rect -49350 32536 -49298 32574
rect -49350 32529 -49341 32536
rect -49341 32529 -49307 32536
rect -49307 32529 -49298 32536
rect -49350 32502 -49341 32517
rect -49341 32502 -49307 32517
rect -49307 32502 -49298 32517
rect -49350 32465 -49298 32502
rect -49034 32608 -48982 32645
rect -49034 32593 -49025 32608
rect -49025 32593 -48991 32608
rect -48991 32593 -48982 32608
rect -49034 32574 -49025 32581
rect -49025 32574 -48991 32581
rect -48991 32574 -48982 32581
rect -49034 32536 -48982 32574
rect -49034 32529 -49025 32536
rect -49025 32529 -48991 32536
rect -48991 32529 -48982 32536
rect -49034 32502 -49025 32517
rect -49025 32502 -48991 32517
rect -48991 32502 -48982 32517
rect -49034 32465 -48982 32502
rect 2396 32618 2421 32940
rect 2421 32618 2743 32940
rect 2743 32618 2768 32940
rect 2396 32593 2768 32618
rect 3049 33273 3101 33298
rect 3049 33246 3058 33273
rect 3058 33246 3092 33273
rect 3092 33246 3101 33273
rect 3049 33201 3101 33234
rect 3049 33182 3058 33201
rect 3058 33182 3092 33201
rect 3092 33182 3101 33201
rect 3049 33167 3058 33170
rect 3058 33167 3092 33170
rect 3092 33167 3101 33170
rect 3049 33129 3101 33167
rect 3049 33118 3058 33129
rect 3058 33118 3092 33129
rect 3092 33118 3101 33129
rect 3049 33095 3058 33106
rect 3058 33095 3092 33106
rect 3092 33095 3101 33106
rect 3049 33057 3101 33095
rect 3049 33054 3058 33057
rect 3058 33054 3092 33057
rect 3092 33054 3101 33057
rect 3049 33023 3058 33042
rect 3058 33023 3092 33042
rect 3092 33023 3101 33042
rect 3049 32990 3101 33023
rect 3049 32951 3058 32978
rect 3058 32951 3092 32978
rect 3092 32951 3101 32978
rect 3049 32926 3101 32951
rect 3365 33273 3417 33298
rect 3365 33246 3374 33273
rect 3374 33246 3408 33273
rect 3408 33246 3417 33273
rect 3365 33201 3417 33234
rect 3365 33182 3374 33201
rect 3374 33182 3408 33201
rect 3408 33182 3417 33201
rect 3365 33167 3374 33170
rect 3374 33167 3408 33170
rect 3408 33167 3417 33170
rect 3365 33129 3417 33167
rect 3365 33118 3374 33129
rect 3374 33118 3408 33129
rect 3408 33118 3417 33129
rect 3365 33095 3374 33106
rect 3374 33095 3408 33106
rect 3408 33095 3417 33106
rect 3365 33057 3417 33095
rect 3365 33054 3374 33057
rect 3374 33054 3408 33057
rect 3408 33054 3417 33057
rect 3365 33023 3374 33042
rect 3374 33023 3408 33042
rect 3408 33023 3417 33042
rect 3365 32990 3417 33023
rect 3365 32951 3374 32978
rect 3374 32951 3408 32978
rect 3408 32951 3417 32978
rect 3365 32926 3417 32951
rect 3681 33273 3733 33298
rect 3681 33246 3690 33273
rect 3690 33246 3724 33273
rect 3724 33246 3733 33273
rect 3681 33201 3733 33234
rect 3681 33182 3690 33201
rect 3690 33182 3724 33201
rect 3724 33182 3733 33201
rect 3681 33167 3690 33170
rect 3690 33167 3724 33170
rect 3724 33167 3733 33170
rect 3681 33129 3733 33167
rect 3681 33118 3690 33129
rect 3690 33118 3724 33129
rect 3724 33118 3733 33129
rect 3681 33095 3690 33106
rect 3690 33095 3724 33106
rect 3724 33095 3733 33106
rect 3681 33057 3733 33095
rect 3681 33054 3690 33057
rect 3690 33054 3724 33057
rect 3724 33054 3733 33057
rect 3681 33023 3690 33042
rect 3690 33023 3724 33042
rect 3724 33023 3733 33042
rect 3681 32990 3733 33023
rect 3681 32951 3690 32978
rect 3690 32951 3724 32978
rect 3724 32951 3733 32978
rect 3681 32926 3733 32951
rect 3997 33273 4049 33298
rect 3997 33246 4006 33273
rect 4006 33246 4040 33273
rect 4040 33246 4049 33273
rect 3997 33201 4049 33234
rect 3997 33182 4006 33201
rect 4006 33182 4040 33201
rect 4040 33182 4049 33201
rect 3997 33167 4006 33170
rect 4006 33167 4040 33170
rect 4040 33167 4049 33170
rect 3997 33129 4049 33167
rect 3997 33118 4006 33129
rect 4006 33118 4040 33129
rect 4040 33118 4049 33129
rect 3997 33095 4006 33106
rect 4006 33095 4040 33106
rect 4040 33095 4049 33106
rect 3997 33057 4049 33095
rect 3997 33054 4006 33057
rect 4006 33054 4040 33057
rect 4040 33054 4049 33057
rect 3997 33023 4006 33042
rect 4006 33023 4040 33042
rect 4040 33023 4049 33042
rect 3997 32990 4049 33023
rect 3997 32951 4006 32978
rect 4006 32951 4040 32978
rect 4040 32951 4049 32978
rect 3997 32926 4049 32951
rect 4313 33273 4365 33298
rect 4313 33246 4322 33273
rect 4322 33246 4356 33273
rect 4356 33246 4365 33273
rect 4313 33201 4365 33234
rect 4313 33182 4322 33201
rect 4322 33182 4356 33201
rect 4356 33182 4365 33201
rect 4313 33167 4322 33170
rect 4322 33167 4356 33170
rect 4356 33167 4365 33170
rect 4313 33129 4365 33167
rect 4313 33118 4322 33129
rect 4322 33118 4356 33129
rect 4356 33118 4365 33129
rect 4313 33095 4322 33106
rect 4322 33095 4356 33106
rect 4356 33095 4365 33106
rect 4313 33057 4365 33095
rect 4313 33054 4322 33057
rect 4322 33054 4356 33057
rect 4356 33054 4365 33057
rect 4313 33023 4322 33042
rect 4322 33023 4356 33042
rect 4356 33023 4365 33042
rect 4313 32990 4365 33023
rect 4313 32951 4322 32978
rect 4322 32951 4356 32978
rect 4356 32951 4365 32978
rect 4313 32926 4365 32951
rect 10000 33236 10308 33864
rect 11000 33236 11308 33864
rect 12000 33236 12308 33864
rect 13000 33236 13308 33864
rect 14000 33236 14308 33864
rect 15000 33236 15308 33864
rect 16000 33236 16308 33864
rect 17000 33236 17308 33864
rect 18000 33236 18308 33864
rect 19000 33236 19308 33864
rect 20000 33236 20308 33864
rect 21000 33236 21308 33864
rect 22000 33236 22308 33864
rect 23000 33236 23308 33864
rect 24000 33236 24308 33864
rect 25000 33236 25308 33864
rect 26000 33236 26308 33864
rect 27000 33236 27308 33864
rect 28000 33236 28308 33864
rect 29000 33236 29308 33864
rect 30000 33236 30308 33864
rect 31000 33236 31308 33864
rect 32000 33236 32308 33864
rect 33000 33236 33308 33864
rect 34000 33236 34308 33864
rect 9660 32896 9968 33204
rect 10032 32928 10276 33172
rect 10340 32896 10968 33204
rect 11032 32928 11276 33172
rect 11340 32896 11968 33204
rect 12032 32928 12276 33172
rect 12340 32896 12968 33204
rect 13032 32928 13276 33172
rect 13340 32896 13968 33204
rect 14032 32928 14276 33172
rect 14340 32896 14968 33204
rect 15032 32928 15276 33172
rect 15340 32896 15968 33204
rect 16032 32928 16276 33172
rect 16340 32896 16968 33204
rect 17032 32928 17276 33172
rect 17340 32896 17968 33204
rect 18032 32928 18276 33172
rect 18340 32896 18968 33204
rect 19032 32928 19276 33172
rect 19340 32896 19968 33204
rect 20032 32928 20276 33172
rect 20340 32896 20968 33204
rect 21032 32928 21276 33172
rect 21340 32896 21968 33204
rect 22032 32928 22276 33172
rect 22340 32896 22968 33204
rect 23032 32928 23276 33172
rect 23340 32896 23968 33204
rect 24032 32928 24276 33172
rect 24340 32896 24968 33204
rect 25032 32928 25276 33172
rect 25340 32896 25968 33204
rect 26032 32928 26276 33172
rect 26340 32896 26968 33204
rect 27032 32928 27276 33172
rect 27340 32896 27968 33204
rect 28032 32928 28276 33172
rect 28340 32896 28968 33204
rect 29032 32928 29276 33172
rect 29340 32896 29968 33204
rect 30032 32928 30276 33172
rect 30340 32896 30968 33204
rect 31032 32928 31276 33172
rect 31340 32896 31968 33204
rect 32032 32928 32276 33172
rect 32340 32896 32968 33204
rect 33032 32928 33276 33172
rect 33340 32896 33968 33204
rect 34032 32928 34276 33172
rect 34340 32896 34648 33204
rect 3049 32608 3101 32645
rect 3049 32593 3058 32608
rect 3058 32593 3092 32608
rect 3092 32593 3101 32608
rect 3049 32574 3058 32581
rect 3058 32574 3092 32581
rect 3092 32574 3101 32581
rect 3049 32536 3101 32574
rect 3049 32529 3058 32536
rect 3058 32529 3092 32536
rect 3092 32529 3101 32536
rect 3049 32502 3058 32517
rect 3058 32502 3092 32517
rect 3092 32502 3101 32517
rect 3049 32465 3101 32502
rect 3365 32608 3417 32645
rect 3365 32593 3374 32608
rect 3374 32593 3408 32608
rect 3408 32593 3417 32608
rect 3365 32574 3374 32581
rect 3374 32574 3408 32581
rect 3408 32574 3417 32581
rect 3365 32536 3417 32574
rect 3365 32529 3374 32536
rect 3374 32529 3408 32536
rect 3408 32529 3417 32536
rect 3365 32502 3374 32517
rect 3374 32502 3408 32517
rect 3408 32502 3417 32517
rect 3365 32465 3417 32502
rect 3681 32608 3733 32645
rect 3681 32593 3690 32608
rect 3690 32593 3724 32608
rect 3724 32593 3733 32608
rect 3681 32574 3690 32581
rect 3690 32574 3724 32581
rect 3724 32574 3733 32581
rect 3681 32536 3733 32574
rect 3681 32529 3690 32536
rect 3690 32529 3724 32536
rect 3724 32529 3733 32536
rect 3681 32502 3690 32517
rect 3690 32502 3724 32517
rect 3724 32502 3733 32517
rect 3681 32465 3733 32502
rect 3997 32608 4049 32645
rect 3997 32593 4006 32608
rect 4006 32593 4040 32608
rect 4040 32593 4049 32608
rect 3997 32574 4006 32581
rect 4006 32574 4040 32581
rect 4040 32574 4049 32581
rect 3997 32536 4049 32574
rect 3997 32529 4006 32536
rect 4006 32529 4040 32536
rect 4040 32529 4049 32536
rect 3997 32502 4006 32517
rect 4006 32502 4040 32517
rect 4040 32502 4049 32517
rect 3997 32465 4049 32502
rect 4313 32608 4365 32645
rect 4313 32593 4322 32608
rect 4322 32593 4356 32608
rect 4356 32593 4365 32608
rect 4313 32574 4322 32581
rect 4322 32574 4356 32581
rect 4356 32574 4365 32581
rect 4313 32536 4365 32574
rect 4313 32529 4322 32536
rect 4322 32529 4356 32536
rect 4356 32529 4365 32536
rect 4313 32502 4322 32517
rect 4322 32502 4356 32517
rect 4356 32502 4365 32517
rect 4313 32465 4365 32502
rect 10000 32236 10308 32864
rect 11000 32236 11308 32864
rect 12000 32236 12308 32864
rect 13000 32236 13308 32864
rect 14000 32236 14308 32864
rect 15000 32236 15308 32864
rect 16000 32236 16308 32864
rect 17000 32236 17308 32864
rect 18000 32236 18308 32864
rect 19000 32236 19308 32864
rect 20000 32236 20308 32864
rect 21000 32236 21308 32864
rect 22000 32236 22308 32864
rect 23000 32236 23308 32864
rect 24000 32236 24308 32864
rect 25000 32236 25308 32864
rect 26000 32236 26308 32864
rect 27000 32236 27308 32864
rect 28000 32236 28308 32864
rect 29000 32236 29308 32864
rect 30000 32236 30308 32864
rect 31000 32236 31308 32864
rect 32000 32236 32308 32864
rect 33000 32236 33308 32864
rect 34000 32236 34308 32864
rect -74479 31236 -74171 31864
rect -73479 31236 -73171 31864
rect -72479 31236 -72171 31864
rect -71479 31236 -71171 31864
rect -70479 31236 -70171 31864
rect -69479 31236 -69171 31864
rect -68479 31236 -68171 31864
rect -67479 31236 -67171 31864
rect -66479 31236 -66171 31864
rect -65479 31236 -65171 31864
rect -64479 31236 -64171 31864
rect -63479 31236 -63171 31864
rect -62479 31236 -62171 31864
rect -61479 31236 -61171 31864
rect -60479 31236 -60171 31864
rect -59479 31236 -59171 31864
rect 9660 31896 9968 32204
rect 10032 31928 10276 32172
rect 10340 31896 10968 32204
rect 11032 31928 11276 32172
rect 11340 31896 11968 32204
rect 12032 31928 12276 32172
rect 12340 31896 12968 32204
rect 13032 31928 13276 32172
rect 13340 31896 13968 32204
rect 14032 31928 14276 32172
rect 14340 31896 14968 32204
rect 15032 31928 15276 32172
rect 15340 31896 15968 32204
rect 16032 31928 16276 32172
rect 16340 31896 16968 32204
rect 17032 31928 17276 32172
rect 17340 31896 17968 32204
rect 18032 31928 18276 32172
rect 18340 31896 18968 32204
rect 19032 31928 19276 32172
rect 19340 31896 19968 32204
rect 20032 31928 20276 32172
rect 20340 31896 20968 32204
rect 21032 31928 21276 32172
rect 21340 31896 21968 32204
rect 22032 31928 22276 32172
rect 22340 31896 22968 32204
rect 23032 31928 23276 32172
rect 23340 31896 23968 32204
rect 24032 31928 24276 32172
rect 24340 31896 24968 32204
rect 25032 31928 25276 32172
rect 25340 31896 25968 32204
rect 26032 31928 26276 32172
rect 26340 31896 26968 32204
rect 27032 31928 27276 32172
rect 27340 31896 27968 32204
rect 28032 31928 28276 32172
rect 28340 31896 28968 32204
rect 29032 31928 29276 32172
rect 29340 31896 29968 32204
rect 30032 31928 30276 32172
rect 30340 31896 30968 32204
rect 31032 31928 31276 32172
rect 31340 31896 31968 32204
rect 32032 31928 32276 32172
rect 32340 31896 32968 32204
rect 33032 31928 33276 32172
rect 33340 31896 33968 32204
rect 34032 31928 34276 32172
rect 34340 31896 34648 32204
rect 10000 31236 10308 31864
rect 11000 31236 11308 31864
rect 12000 31236 12308 31864
rect 13000 31236 13308 31864
rect 14000 31236 14308 31864
rect 15000 31236 15308 31864
rect 16000 31236 16308 31864
rect 17000 31236 17308 31864
rect 18000 31236 18308 31864
rect 19000 31236 19308 31864
rect 20000 31236 20308 31864
rect 21000 31236 21308 31864
rect 22000 31236 22308 31864
rect 23000 31236 23308 31864
rect 24000 31236 24308 31864
rect 25000 31236 25308 31864
rect 26000 31236 26308 31864
rect 27000 31236 27308 31864
rect 28000 31236 28308 31864
rect 29000 31236 29308 31864
rect 30000 31236 30308 31864
rect 31000 31236 31308 31864
rect 32000 31236 32308 31864
rect 33000 31236 33308 31864
rect 34000 31236 34308 31864
rect -74819 30896 -74511 31204
rect -74447 30928 -74203 31172
rect -74139 30896 -73511 31204
rect -73447 30928 -73203 31172
rect -73139 30896 -72511 31204
rect -72447 30928 -72203 31172
rect -72139 30896 -71511 31204
rect -71447 30928 -71203 31172
rect -71139 30896 -70511 31204
rect -70447 30928 -70203 31172
rect -70139 30896 -69511 31204
rect -69447 30928 -69203 31172
rect -69139 30896 -68511 31204
rect -68447 30928 -68203 31172
rect -68139 30896 -67511 31204
rect -67447 30928 -67203 31172
rect -67139 30896 -66511 31204
rect -66447 30928 -66203 31172
rect -66139 30896 -65511 31204
rect -65447 30928 -65203 31172
rect -65139 30896 -64511 31204
rect -64447 30928 -64203 31172
rect -64139 30896 -63511 31204
rect -63447 30928 -63203 31172
rect -63139 30896 -62511 31204
rect -62447 30928 -62203 31172
rect -62139 30896 -61511 31204
rect -61447 30928 -61203 31172
rect -61139 30896 -60511 31204
rect -60447 30928 -60203 31172
rect -60139 30896 -59511 31204
rect -59447 30928 -59203 31172
rect -59139 30896 -58831 31204
rect 9660 30896 9968 31204
rect 10032 30928 10276 31172
rect 10340 30896 10968 31204
rect 11032 30928 11276 31172
rect 11340 30896 11968 31204
rect 12032 30928 12276 31172
rect 12340 30896 12968 31204
rect 13032 30928 13276 31172
rect 13340 30896 13968 31204
rect 14032 30928 14276 31172
rect 14340 30896 14968 31204
rect 15032 30928 15276 31172
rect 15340 30896 15968 31204
rect 16032 30928 16276 31172
rect 16340 30896 16968 31204
rect 17032 30928 17276 31172
rect 17340 30896 17968 31204
rect 18032 30928 18276 31172
rect 18340 30896 18968 31204
rect 19032 30928 19276 31172
rect 19340 30896 19968 31204
rect 20032 30928 20276 31172
rect 20340 30896 20968 31204
rect 21032 30928 21276 31172
rect 21340 30896 21968 31204
rect 22032 30928 22276 31172
rect 22340 30896 22968 31204
rect 23032 30928 23276 31172
rect 23340 30896 23968 31204
rect 24032 30928 24276 31172
rect 24340 30896 24968 31204
rect 25032 30928 25276 31172
rect 25340 30896 25968 31204
rect 26032 30928 26276 31172
rect 26340 30896 26968 31204
rect 27032 30928 27276 31172
rect 27340 30896 27968 31204
rect 28032 30928 28276 31172
rect 28340 30896 28968 31204
rect 29032 30928 29276 31172
rect 29340 30896 29968 31204
rect 30032 30928 30276 31172
rect 30340 30896 30968 31204
rect 31032 30928 31276 31172
rect 31340 30896 31968 31204
rect 32032 30928 32276 31172
rect 32340 30896 32968 31204
rect 33032 30928 33276 31172
rect 33340 30896 33968 31204
rect 34032 30928 34276 31172
rect 34340 30896 34648 31204
rect -74479 30236 -74171 30864
rect -73479 30236 -73171 30864
rect -72479 30236 -72171 30864
rect -71479 30236 -71171 30864
rect -70479 30236 -70171 30864
rect -69479 30236 -69171 30864
rect -68479 30236 -68171 30864
rect -67479 30236 -67171 30864
rect -66479 30236 -66171 30864
rect -65479 30236 -65171 30864
rect -64479 30236 -64171 30864
rect -63479 30236 -63171 30864
rect -62479 30236 -62171 30864
rect -61479 30236 -61171 30864
rect -60479 30236 -60171 30864
rect -59479 30236 -59171 30864
rect 10000 30236 10308 30864
rect 11000 30236 11308 30864
rect 12000 30236 12308 30864
rect 13000 30236 13308 30864
rect 14000 30236 14308 30864
rect 15000 30236 15308 30864
rect 16000 30236 16308 30864
rect 17000 30236 17308 30864
rect 18000 30236 18308 30864
rect 19000 30236 19308 30864
rect 20000 30236 20308 30864
rect 21000 30236 21308 30864
rect 22000 30236 22308 30864
rect 23000 30236 23308 30864
rect 24000 30236 24308 30864
rect 25000 30236 25308 30864
rect 26000 30236 26308 30864
rect 27000 30236 27308 30864
rect 28000 30236 28308 30864
rect 29000 30236 29308 30864
rect 30000 30236 30308 30864
rect 31000 30236 31308 30864
rect 32000 30236 32308 30864
rect 33000 30236 33308 30864
rect 34000 30236 34308 30864
rect -74819 29896 -74511 30204
rect -74447 29928 -74203 30172
rect -74139 29896 -73511 30204
rect -73447 29928 -73203 30172
rect -73139 29896 -72511 30204
rect -72447 29928 -72203 30172
rect -72139 29896 -71511 30204
rect -71447 29928 -71203 30172
rect -71139 29896 -70511 30204
rect -70447 29928 -70203 30172
rect -70139 29896 -69511 30204
rect -69447 29928 -69203 30172
rect -69139 29896 -68511 30204
rect -68447 29928 -68203 30172
rect -68139 29896 -67511 30204
rect -67447 29928 -67203 30172
rect -67139 29896 -66511 30204
rect -66447 29928 -66203 30172
rect -66139 29896 -65511 30204
rect -65447 29928 -65203 30172
rect -65139 29896 -64511 30204
rect -64447 29928 -64203 30172
rect -64139 29896 -63511 30204
rect -63447 29928 -63203 30172
rect -63139 29896 -62511 30204
rect -62447 29928 -62203 30172
rect -62139 29896 -61511 30204
rect -61447 29928 -61203 30172
rect -61139 29896 -60511 30204
rect -60447 29928 -60203 30172
rect -60139 29896 -59511 30204
rect -59447 29928 -59203 30172
rect -59139 29896 -58831 30204
rect 9660 29896 9968 30204
rect 10032 29928 10276 30172
rect 10340 29896 10968 30204
rect 11032 29928 11276 30172
rect 11340 29896 11968 30204
rect 12032 29928 12276 30172
rect 12340 29896 12968 30204
rect 13032 29928 13276 30172
rect 13340 29896 13968 30204
rect 14032 29928 14276 30172
rect 14340 29896 14968 30204
rect 15032 29928 15276 30172
rect 15340 29896 15968 30204
rect 16032 29928 16276 30172
rect 16340 29896 16968 30204
rect 17032 29928 17276 30172
rect 17340 29896 17968 30204
rect 18032 29928 18276 30172
rect 18340 29896 18968 30204
rect 19032 29928 19276 30172
rect 19340 29896 19968 30204
rect 20032 29928 20276 30172
rect 20340 29896 20968 30204
rect 21032 29928 21276 30172
rect 21340 29896 21968 30204
rect 22032 29928 22276 30172
rect 22340 29896 22968 30204
rect 23032 29928 23276 30172
rect 23340 29896 23968 30204
rect 24032 29928 24276 30172
rect 24340 29896 24968 30204
rect 25032 29928 25276 30172
rect 25340 29896 25968 30204
rect 26032 29928 26276 30172
rect 26340 29896 26968 30204
rect 27032 29928 27276 30172
rect 27340 29896 27968 30204
rect 28032 29928 28276 30172
rect 28340 29896 28968 30204
rect 29032 29928 29276 30172
rect 29340 29896 29968 30204
rect 30032 29928 30276 30172
rect 30340 29896 30968 30204
rect 31032 29928 31276 30172
rect 31340 29896 31968 30204
rect 32032 29928 32276 30172
rect 32340 29896 32968 30204
rect 33032 29928 33276 30172
rect 33340 29896 33968 30204
rect 34032 29928 34276 30172
rect 34340 29896 34648 30204
rect -74479 29236 -74171 29864
rect -73479 29236 -73171 29864
rect -72479 29236 -72171 29864
rect -71479 29236 -71171 29864
rect -70479 29236 -70171 29864
rect -69479 29236 -69171 29864
rect -68479 29236 -68171 29864
rect -67479 29236 -67171 29864
rect -66479 29236 -66171 29864
rect -65479 29236 -65171 29864
rect -64479 29236 -64171 29864
rect -63479 29236 -63171 29864
rect -62479 29236 -62171 29864
rect -61479 29236 -61171 29864
rect -60479 29236 -60171 29864
rect -59479 29236 -59171 29864
rect 10000 29236 10308 29864
rect 11000 29236 11308 29864
rect 12000 29236 12308 29864
rect 13000 29236 13308 29864
rect 14000 29236 14308 29864
rect 15000 29236 15308 29864
rect 16000 29236 16308 29864
rect 17000 29236 17308 29864
rect 18000 29236 18308 29864
rect 19000 29236 19308 29864
rect 20000 29236 20308 29864
rect 21000 29236 21308 29864
rect 22000 29236 22308 29864
rect 23000 29236 23308 29864
rect 24000 29236 24308 29864
rect 25000 29236 25308 29864
rect 26000 29236 26308 29864
rect 27000 29236 27308 29864
rect 28000 29236 28308 29864
rect 29000 29236 29308 29864
rect 30000 29236 30308 29864
rect 31000 29236 31308 29864
rect 32000 29236 32308 29864
rect 33000 29236 33308 29864
rect 34000 29236 34308 29864
rect -74819 28896 -74511 29204
rect -74447 28928 -74203 29172
rect -74139 28896 -73511 29204
rect -73447 28928 -73203 29172
rect -73139 28896 -72511 29204
rect -72447 28928 -72203 29172
rect -72139 28896 -71511 29204
rect -71447 28928 -71203 29172
rect -71139 28896 -70511 29204
rect -70447 28928 -70203 29172
rect -70139 28896 -69511 29204
rect -69447 28928 -69203 29172
rect -69139 28896 -68511 29204
rect -68447 28928 -68203 29172
rect -68139 28896 -67511 29204
rect -67447 28928 -67203 29172
rect -67139 28896 -66511 29204
rect -66447 28928 -66203 29172
rect -66139 28896 -65511 29204
rect -65447 28928 -65203 29172
rect -65139 28896 -64511 29204
rect -64447 28928 -64203 29172
rect -64139 28896 -63511 29204
rect -63447 28928 -63203 29172
rect -63139 28896 -62511 29204
rect -62447 28928 -62203 29172
rect -62139 28896 -61511 29204
rect -61447 28928 -61203 29172
rect -61139 28896 -60511 29204
rect -60447 28928 -60203 29172
rect -60139 28896 -59511 29204
rect -59447 28928 -59203 29172
rect -59139 28896 -58831 29204
rect 9660 28896 9968 29204
rect 10032 28928 10276 29172
rect 10340 28896 10968 29204
rect 11032 28928 11276 29172
rect 11340 28896 11968 29204
rect 12032 28928 12276 29172
rect 12340 28896 12968 29204
rect 13032 28928 13276 29172
rect 13340 28896 13968 29204
rect 14032 28928 14276 29172
rect 14340 28896 14968 29204
rect 15032 28928 15276 29172
rect 15340 28896 15968 29204
rect 16032 28928 16276 29172
rect 16340 28896 16968 29204
rect 17032 28928 17276 29172
rect 17340 28896 17968 29204
rect 18032 28928 18276 29172
rect 18340 28896 18968 29204
rect 19032 28928 19276 29172
rect 19340 28896 19968 29204
rect 20032 28928 20276 29172
rect 20340 28896 20968 29204
rect 21032 28928 21276 29172
rect 21340 28896 21968 29204
rect 22032 28928 22276 29172
rect 22340 28896 22968 29204
rect 23032 28928 23276 29172
rect 23340 28896 23968 29204
rect 24032 28928 24276 29172
rect 24340 28896 24968 29204
rect 25032 28928 25276 29172
rect 25340 28896 25968 29204
rect 26032 28928 26276 29172
rect 26340 28896 26968 29204
rect 27032 28928 27276 29172
rect 27340 28896 27968 29204
rect 28032 28928 28276 29172
rect 28340 28896 28968 29204
rect 29032 28928 29276 29172
rect 29340 28896 29968 29204
rect 30032 28928 30276 29172
rect 30340 28896 30968 29204
rect 31032 28928 31276 29172
rect 31340 28896 31968 29204
rect 32032 28928 32276 29172
rect 32340 28896 32968 29204
rect 33032 28928 33276 29172
rect 33340 28896 33968 29204
rect 34032 28928 34276 29172
rect 34340 28896 34648 29204
rect -74479 28556 -74171 28864
rect -73479 28556 -73171 28864
rect -72479 28556 -72171 28864
rect -71479 28556 -71171 28864
rect -70479 28556 -70171 28864
rect -69479 28556 -69171 28864
rect -68479 28556 -68171 28864
rect -67479 28556 -67171 28864
rect -66479 28556 -66171 28864
rect -65479 28556 -65171 28864
rect -64479 28556 -64171 28864
rect -63479 28556 -63171 28864
rect -62479 28556 -62171 28864
rect -61479 28556 -61171 28864
rect -60479 28556 -60171 28864
rect -59479 28556 -59171 28864
rect 10000 28556 10308 28864
rect 11000 28556 11308 28864
rect 12000 28556 12308 28864
rect 13000 28556 13308 28864
rect 14000 28556 14308 28864
rect 15000 28556 15308 28864
rect 16000 28556 16308 28864
rect 17000 28556 17308 28864
rect 18000 28556 18308 28864
rect 19000 28556 19308 28864
rect 20000 28556 20308 28864
rect 21000 28556 21308 28864
rect 22000 28556 22308 28864
rect 23000 28556 23308 28864
rect 24000 28556 24308 28864
rect 25000 28556 25308 28864
rect 26000 28556 26308 28864
rect 27000 28556 27308 28864
rect 28000 28556 28308 28864
rect 29000 28556 29308 28864
rect 30000 28556 30308 28864
rect 31000 28556 31308 28864
rect 32000 28556 32308 28864
rect 33000 28556 33308 28864
rect 34000 28556 34308 28864
rect -72776 16041 -60884 25949
rect -47607 25523 -47043 26087
rect 6638 25567 7202 26131
rect -21212 13856 -19304 15124
rect 20324 16046 32216 25954
rect -42408 7880 -40692 13820
rect 142 7880 1858 13820
rect -42408 -2298 -40692 2298
rect 142 -2298 1858 2298
rect -42408 -13820 -40692 -7880
rect 142 -13820 1858 -7880
rect -72776 -25954 -60884 -16046
rect 20324 -25954 32216 -16046
rect -74479 -28864 -74171 -28556
rect -73479 -28864 -73171 -28556
rect -72479 -28864 -72171 -28556
rect -71479 -28864 -71171 -28556
rect -70479 -28864 -70171 -28556
rect -69479 -28864 -69171 -28556
rect -68479 -28864 -68171 -28556
rect -67479 -28864 -67171 -28556
rect -66479 -28864 -66171 -28556
rect -65479 -28864 -65171 -28556
rect -64479 -28864 -64171 -28556
rect -63479 -28864 -63171 -28556
rect -62479 -28864 -62171 -28556
rect -61479 -28864 -61171 -28556
rect -60479 -28864 -60171 -28556
rect -59479 -28864 -59171 -28556
rect -58479 -28864 -58171 -28556
rect -57479 -28864 -57171 -28556
rect -56479 -28864 -56171 -28556
rect -55479 -28864 -55171 -28556
rect -54479 -28864 -54171 -28556
rect -53479 -28864 -53171 -28556
rect -52479 -28864 -52171 -28556
rect -51479 -28864 -51171 -28556
rect -50479 -28864 -50171 -28556
rect -49479 -28864 -49171 -28556
rect 8621 -28864 8929 -28556
rect 9621 -28864 9929 -28556
rect 10621 -28864 10929 -28556
rect 11621 -28864 11929 -28556
rect 12621 -28864 12929 -28556
rect 13621 -28864 13929 -28556
rect 14621 -28864 14929 -28556
rect 15621 -28864 15929 -28556
rect 16621 -28864 16929 -28556
rect 17621 -28864 17929 -28556
rect 18621 -28864 18929 -28556
rect 19621 -28864 19929 -28556
rect 20621 -28864 20929 -28556
rect 21621 -28864 21929 -28556
rect 22621 -28864 22929 -28556
rect 23621 -28864 23929 -28556
rect 24621 -28864 24929 -28556
rect 25621 -28864 25929 -28556
rect 26621 -28864 26929 -28556
rect 27621 -28864 27929 -28556
rect 28621 -28864 28929 -28556
rect 29621 -28864 29929 -28556
rect 30621 -28864 30929 -28556
rect 31621 -28864 31929 -28556
rect 32621 -28864 32929 -28556
rect 33621 -28864 33929 -28556
rect -74819 -29204 -74511 -28896
rect -74447 -29172 -74203 -28928
rect -74139 -29204 -73511 -28896
rect -73447 -29172 -73203 -28928
rect -73139 -29204 -72511 -28896
rect -72447 -29172 -72203 -28928
rect -72139 -29204 -71511 -28896
rect -71447 -29172 -71203 -28928
rect -71139 -29204 -70511 -28896
rect -70447 -29172 -70203 -28928
rect -70139 -29204 -69511 -28896
rect -69447 -29172 -69203 -28928
rect -69139 -29204 -68511 -28896
rect -68447 -29172 -68203 -28928
rect -68139 -29204 -67511 -28896
rect -67447 -29172 -67203 -28928
rect -67139 -29204 -66511 -28896
rect -66447 -29172 -66203 -28928
rect -66139 -29204 -65511 -28896
rect -65447 -29172 -65203 -28928
rect -65139 -29204 -64511 -28896
rect -64447 -29172 -64203 -28928
rect -64139 -29204 -63511 -28896
rect -63447 -29172 -63203 -28928
rect -63139 -29204 -62511 -28896
rect -62447 -29172 -62203 -28928
rect -62139 -29204 -61511 -28896
rect -61447 -29172 -61203 -28928
rect -61139 -29204 -60511 -28896
rect -60447 -29172 -60203 -28928
rect -60139 -29204 -59511 -28896
rect -59447 -29172 -59203 -28928
rect -59139 -29204 -58511 -28896
rect -58447 -29172 -58203 -28928
rect -58139 -29204 -57511 -28896
rect -57447 -29172 -57203 -28928
rect -57139 -29204 -56511 -28896
rect -56447 -29172 -56203 -28928
rect -56139 -29204 -55511 -28896
rect -55447 -29172 -55203 -28928
rect -55139 -29204 -54511 -28896
rect -54447 -29172 -54203 -28928
rect -54139 -29204 -53511 -28896
rect -53447 -29172 -53203 -28928
rect -53139 -29204 -52511 -28896
rect -52447 -29172 -52203 -28928
rect -52139 -29204 -51511 -28896
rect -51447 -29172 -51203 -28928
rect -51139 -29204 -50511 -28896
rect -50447 -29172 -50203 -28928
rect -50139 -29204 -49511 -28896
rect -49447 -29172 -49203 -28928
rect -49139 -29204 -48831 -28896
rect 8281 -29204 8589 -28896
rect 8653 -29172 8897 -28928
rect 8961 -29204 9589 -28896
rect 9653 -29172 9897 -28928
rect 9961 -29204 10589 -28896
rect 10653 -29172 10897 -28928
rect 10961 -29204 11589 -28896
rect 11653 -29172 11897 -28928
rect 11961 -29204 12589 -28896
rect 12653 -29172 12897 -28928
rect 12961 -29204 13589 -28896
rect 13653 -29172 13897 -28928
rect 13961 -29204 14589 -28896
rect 14653 -29172 14897 -28928
rect 14961 -29204 15589 -28896
rect 15653 -29172 15897 -28928
rect 15961 -29204 16589 -28896
rect 16653 -29172 16897 -28928
rect 16961 -29204 17589 -28896
rect 17653 -29172 17897 -28928
rect 17961 -29204 18589 -28896
rect 18653 -29172 18897 -28928
rect 18961 -29204 19589 -28896
rect 19653 -29172 19897 -28928
rect 19961 -29204 20589 -28896
rect 20653 -29172 20897 -28928
rect 20961 -29204 21589 -28896
rect 21653 -29172 21897 -28928
rect 21961 -29204 22589 -28896
rect 22653 -29172 22897 -28928
rect 22961 -29204 23589 -28896
rect 23653 -29172 23897 -28928
rect 23961 -29204 24589 -28896
rect 24653 -29172 24897 -28928
rect 24961 -29204 25589 -28896
rect 25653 -29172 25897 -28928
rect 25961 -29204 26589 -28896
rect 26653 -29172 26897 -28928
rect 26961 -29204 27589 -28896
rect 27653 -29172 27897 -28928
rect 27961 -29204 28589 -28896
rect 28653 -29172 28897 -28928
rect 28961 -29204 29589 -28896
rect 29653 -29172 29897 -28928
rect 29961 -29204 30589 -28896
rect 30653 -29172 30897 -28928
rect 30961 -29204 31589 -28896
rect 31653 -29172 31897 -28928
rect 31961 -29204 32589 -28896
rect 32653 -29172 32897 -28928
rect 32961 -29204 33589 -28896
rect 33653 -29172 33897 -28928
rect 33961 -29204 34269 -28896
rect -74479 -29864 -74171 -29236
rect -73479 -29864 -73171 -29236
rect -72479 -29864 -72171 -29236
rect -71479 -29864 -71171 -29236
rect -70479 -29864 -70171 -29236
rect -69479 -29864 -69171 -29236
rect -68479 -29864 -68171 -29236
rect -67479 -29864 -67171 -29236
rect -66479 -29864 -66171 -29236
rect -65479 -29864 -65171 -29236
rect -64479 -29864 -64171 -29236
rect -63479 -29864 -63171 -29236
rect -62479 -29864 -62171 -29236
rect -61479 -29864 -61171 -29236
rect -60479 -29864 -60171 -29236
rect -59479 -29864 -59171 -29236
rect -58479 -29864 -58171 -29236
rect -57479 -29864 -57171 -29236
rect -56479 -29864 -56171 -29236
rect -55479 -29864 -55171 -29236
rect -54479 -29864 -54171 -29236
rect -53479 -29864 -53171 -29236
rect -52479 -29864 -52171 -29236
rect -51479 -29864 -51171 -29236
rect -50479 -29864 -50171 -29236
rect -49479 -29864 -49171 -29236
rect 8621 -29864 8929 -29236
rect 9621 -29864 9929 -29236
rect 10621 -29864 10929 -29236
rect 11621 -29864 11929 -29236
rect 12621 -29864 12929 -29236
rect 13621 -29864 13929 -29236
rect 14621 -29864 14929 -29236
rect 15621 -29864 15929 -29236
rect 16621 -29864 16929 -29236
rect 17621 -29864 17929 -29236
rect 18621 -29864 18929 -29236
rect 19621 -29864 19929 -29236
rect 20621 -29864 20929 -29236
rect 21621 -29864 21929 -29236
rect 22621 -29864 22929 -29236
rect 23621 -29864 23929 -29236
rect 24621 -29864 24929 -29236
rect 25621 -29864 25929 -29236
rect 26621 -29864 26929 -29236
rect 27621 -29864 27929 -29236
rect 28621 -29864 28929 -29236
rect 29621 -29864 29929 -29236
rect 30621 -29864 30929 -29236
rect 31621 -29864 31929 -29236
rect 32621 -29864 32929 -29236
rect 33621 -29864 33929 -29236
rect -74819 -30204 -74511 -29896
rect -74447 -30172 -74203 -29928
rect -74139 -30204 -73511 -29896
rect -73447 -30172 -73203 -29928
rect -73139 -30204 -72511 -29896
rect -72447 -30172 -72203 -29928
rect -72139 -30204 -71511 -29896
rect -71447 -30172 -71203 -29928
rect -71139 -30204 -70511 -29896
rect -70447 -30172 -70203 -29928
rect -70139 -30204 -69511 -29896
rect -69447 -30172 -69203 -29928
rect -69139 -30204 -68511 -29896
rect -68447 -30172 -68203 -29928
rect -68139 -30204 -67511 -29896
rect -67447 -30172 -67203 -29928
rect -67139 -30204 -66511 -29896
rect -66447 -30172 -66203 -29928
rect -66139 -30204 -65511 -29896
rect -65447 -30172 -65203 -29928
rect -65139 -30204 -64511 -29896
rect -64447 -30172 -64203 -29928
rect -64139 -30204 -63511 -29896
rect -63447 -30172 -63203 -29928
rect -63139 -30204 -62511 -29896
rect -62447 -30172 -62203 -29928
rect -62139 -30204 -61511 -29896
rect -61447 -30172 -61203 -29928
rect -61139 -30204 -60511 -29896
rect -60447 -30172 -60203 -29928
rect -60139 -30204 -59511 -29896
rect -59447 -30172 -59203 -29928
rect -59139 -30204 -58511 -29896
rect -58447 -30172 -58203 -29928
rect -58139 -30204 -57511 -29896
rect -57447 -30172 -57203 -29928
rect -57139 -30204 -56511 -29896
rect -56447 -30172 -56203 -29928
rect -56139 -30204 -55511 -29896
rect -55447 -30172 -55203 -29928
rect -55139 -30204 -54511 -29896
rect -54447 -30172 -54203 -29928
rect -54139 -30204 -53511 -29896
rect -53447 -30172 -53203 -29928
rect -53139 -30204 -52511 -29896
rect -52447 -30172 -52203 -29928
rect -52139 -30204 -51511 -29896
rect -51447 -30172 -51203 -29928
rect -51139 -30204 -50511 -29896
rect -50447 -30172 -50203 -29928
rect -50139 -30204 -49511 -29896
rect -49447 -30172 -49203 -29928
rect -49139 -30204 -48831 -29896
rect 8281 -30204 8589 -29896
rect 8653 -30172 8897 -29928
rect 8961 -30204 9589 -29896
rect 9653 -30172 9897 -29928
rect 9961 -30204 10589 -29896
rect 10653 -30172 10897 -29928
rect 10961 -30204 11589 -29896
rect 11653 -30172 11897 -29928
rect 11961 -30204 12589 -29896
rect 12653 -30172 12897 -29928
rect 12961 -30204 13589 -29896
rect 13653 -30172 13897 -29928
rect 13961 -30204 14589 -29896
rect 14653 -30172 14897 -29928
rect 14961 -30204 15589 -29896
rect 15653 -30172 15897 -29928
rect 15961 -30204 16589 -29896
rect 16653 -30172 16897 -29928
rect 16961 -30204 17589 -29896
rect 17653 -30172 17897 -29928
rect 17961 -30204 18589 -29896
rect 18653 -30172 18897 -29928
rect 18961 -30204 19589 -29896
rect 19653 -30172 19897 -29928
rect 19961 -30204 20589 -29896
rect 20653 -30172 20897 -29928
rect 20961 -30204 21589 -29896
rect 21653 -30172 21897 -29928
rect 21961 -30204 22589 -29896
rect 22653 -30172 22897 -29928
rect 22961 -30204 23589 -29896
rect 23653 -30172 23897 -29928
rect 23961 -30204 24589 -29896
rect 24653 -30172 24897 -29928
rect 24961 -30204 25589 -29896
rect 25653 -30172 25897 -29928
rect 25961 -30204 26589 -29896
rect 26653 -30172 26897 -29928
rect 26961 -30204 27589 -29896
rect 27653 -30172 27897 -29928
rect 27961 -30204 28589 -29896
rect 28653 -30172 28897 -29928
rect 28961 -30204 29589 -29896
rect 29653 -30172 29897 -29928
rect 29961 -30204 30589 -29896
rect 30653 -30172 30897 -29928
rect 30961 -30204 31589 -29896
rect 31653 -30172 31897 -29928
rect 31961 -30204 32589 -29896
rect 32653 -30172 32897 -29928
rect 32961 -30204 33589 -29896
rect 33653 -30172 33897 -29928
rect 33961 -30204 34269 -29896
rect -74479 -30864 -74171 -30236
rect -73479 -30864 -73171 -30236
rect -72479 -30864 -72171 -30236
rect -71479 -30864 -71171 -30236
rect -70479 -30864 -70171 -30236
rect -69479 -30864 -69171 -30236
rect -68479 -30864 -68171 -30236
rect -67479 -30864 -67171 -30236
rect -66479 -30864 -66171 -30236
rect -65479 -30864 -65171 -30236
rect -64479 -30864 -64171 -30236
rect -63479 -30864 -63171 -30236
rect -62479 -30864 -62171 -30236
rect -61479 -30864 -61171 -30236
rect -60479 -30864 -60171 -30236
rect -59479 -30864 -59171 -30236
rect -58479 -30864 -58171 -30236
rect -57479 -30864 -57171 -30236
rect -56479 -30864 -56171 -30236
rect -55479 -30864 -55171 -30236
rect -54479 -30864 -54171 -30236
rect -53479 -30864 -53171 -30236
rect -52479 -30864 -52171 -30236
rect -51479 -30864 -51171 -30236
rect -50479 -30864 -50171 -30236
rect -49479 -30864 -49171 -30236
rect 8621 -30864 8929 -30236
rect 9621 -30864 9929 -30236
rect 10621 -30864 10929 -30236
rect 11621 -30864 11929 -30236
rect 12621 -30864 12929 -30236
rect 13621 -30864 13929 -30236
rect 14621 -30864 14929 -30236
rect 15621 -30864 15929 -30236
rect 16621 -30864 16929 -30236
rect 17621 -30864 17929 -30236
rect 18621 -30864 18929 -30236
rect 19621 -30864 19929 -30236
rect 20621 -30864 20929 -30236
rect 21621 -30864 21929 -30236
rect 22621 -30864 22929 -30236
rect 23621 -30864 23929 -30236
rect 24621 -30864 24929 -30236
rect 25621 -30864 25929 -30236
rect 26621 -30864 26929 -30236
rect 27621 -30864 27929 -30236
rect 28621 -30864 28929 -30236
rect 29621 -30864 29929 -30236
rect 30621 -30864 30929 -30236
rect 31621 -30864 31929 -30236
rect 32621 -30864 32929 -30236
rect 33621 -30864 33929 -30236
rect -74819 -31204 -74511 -30896
rect -74447 -31172 -74203 -30928
rect -74139 -31204 -73511 -30896
rect -73447 -31172 -73203 -30928
rect -73139 -31204 -72511 -30896
rect -72447 -31172 -72203 -30928
rect -72139 -31204 -71511 -30896
rect -71447 -31172 -71203 -30928
rect -71139 -31204 -70511 -30896
rect -70447 -31172 -70203 -30928
rect -70139 -31204 -69511 -30896
rect -69447 -31172 -69203 -30928
rect -69139 -31204 -68511 -30896
rect -68447 -31172 -68203 -30928
rect -68139 -31204 -67511 -30896
rect -67447 -31172 -67203 -30928
rect -67139 -31204 -66511 -30896
rect -66447 -31172 -66203 -30928
rect -66139 -31204 -65511 -30896
rect -65447 -31172 -65203 -30928
rect -65139 -31204 -64511 -30896
rect -64447 -31172 -64203 -30928
rect -64139 -31204 -63511 -30896
rect -63447 -31172 -63203 -30928
rect -63139 -31204 -62511 -30896
rect -62447 -31172 -62203 -30928
rect -62139 -31204 -61511 -30896
rect -61447 -31172 -61203 -30928
rect -61139 -31204 -60511 -30896
rect -60447 -31172 -60203 -30928
rect -60139 -31204 -59511 -30896
rect -59447 -31172 -59203 -30928
rect -59139 -31204 -58511 -30896
rect -58447 -31172 -58203 -30928
rect -58139 -31204 -57511 -30896
rect -57447 -31172 -57203 -30928
rect -57139 -31204 -56511 -30896
rect -56447 -31172 -56203 -30928
rect -56139 -31204 -55511 -30896
rect -55447 -31172 -55203 -30928
rect -55139 -31204 -54511 -30896
rect -54447 -31172 -54203 -30928
rect -54139 -31204 -53511 -30896
rect -53447 -31172 -53203 -30928
rect -53139 -31204 -52511 -30896
rect -52447 -31172 -52203 -30928
rect -52139 -31204 -51511 -30896
rect -51447 -31172 -51203 -30928
rect -51139 -31204 -50511 -30896
rect -50447 -31172 -50203 -30928
rect -50139 -31204 -49511 -30896
rect -49447 -31172 -49203 -30928
rect -49139 -31204 -48831 -30896
rect 8281 -31204 8589 -30896
rect 8653 -31172 8897 -30928
rect 8961 -31204 9589 -30896
rect 9653 -31172 9897 -30928
rect 9961 -31204 10589 -30896
rect 10653 -31172 10897 -30928
rect 10961 -31204 11589 -30896
rect 11653 -31172 11897 -30928
rect 11961 -31204 12589 -30896
rect 12653 -31172 12897 -30928
rect 12961 -31204 13589 -30896
rect 13653 -31172 13897 -30928
rect 13961 -31204 14589 -30896
rect 14653 -31172 14897 -30928
rect 14961 -31204 15589 -30896
rect 15653 -31172 15897 -30928
rect 15961 -31204 16589 -30896
rect 16653 -31172 16897 -30928
rect 16961 -31204 17589 -30896
rect 17653 -31172 17897 -30928
rect 17961 -31204 18589 -30896
rect 18653 -31172 18897 -30928
rect 18961 -31204 19589 -30896
rect 19653 -31172 19897 -30928
rect 19961 -31204 20589 -30896
rect 20653 -31172 20897 -30928
rect 20961 -31204 21589 -30896
rect 21653 -31172 21897 -30928
rect 21961 -31204 22589 -30896
rect 22653 -31172 22897 -30928
rect 22961 -31204 23589 -30896
rect 23653 -31172 23897 -30928
rect 23961 -31204 24589 -30896
rect 24653 -31172 24897 -30928
rect 24961 -31204 25589 -30896
rect 25653 -31172 25897 -30928
rect 25961 -31204 26589 -30896
rect 26653 -31172 26897 -30928
rect 26961 -31204 27589 -30896
rect 27653 -31172 27897 -30928
rect 27961 -31204 28589 -30896
rect 28653 -31172 28897 -30928
rect 28961 -31204 29589 -30896
rect 29653 -31172 29897 -30928
rect 29961 -31204 30589 -30896
rect 30653 -31172 30897 -30928
rect 30961 -31204 31589 -30896
rect 31653 -31172 31897 -30928
rect 31961 -31204 32589 -30896
rect 32653 -31172 32897 -30928
rect 32961 -31204 33589 -30896
rect 33653 -31172 33897 -30928
rect 33961 -31204 34269 -30896
rect -74479 -31864 -74171 -31236
rect -73479 -31864 -73171 -31236
rect -72479 -31864 -72171 -31236
rect -71479 -31864 -71171 -31236
rect -70479 -31864 -70171 -31236
rect -69479 -31864 -69171 -31236
rect -68479 -31864 -68171 -31236
rect -67479 -31864 -67171 -31236
rect -66479 -31864 -66171 -31236
rect -65479 -31864 -65171 -31236
rect -64479 -31864 -64171 -31236
rect -63479 -31864 -63171 -31236
rect -62479 -31864 -62171 -31236
rect -61479 -31864 -61171 -31236
rect -60479 -31864 -60171 -31236
rect -59479 -31864 -59171 -31236
rect -58479 -31864 -58171 -31236
rect -57479 -31864 -57171 -31236
rect -56479 -31864 -56171 -31236
rect -55479 -31864 -55171 -31236
rect -54479 -31864 -54171 -31236
rect -53479 -31864 -53171 -31236
rect -52479 -31864 -52171 -31236
rect -51479 -31864 -51171 -31236
rect -50479 -31864 -50171 -31236
rect -49479 -31864 -49171 -31236
rect 8621 -31864 8929 -31236
rect 9621 -31864 9929 -31236
rect 10621 -31864 10929 -31236
rect 11621 -31864 11929 -31236
rect 12621 -31864 12929 -31236
rect 13621 -31864 13929 -31236
rect 14621 -31864 14929 -31236
rect 15621 -31864 15929 -31236
rect 16621 -31864 16929 -31236
rect 17621 -31864 17929 -31236
rect 18621 -31864 18929 -31236
rect 19621 -31864 19929 -31236
rect 20621 -31864 20929 -31236
rect 21621 -31864 21929 -31236
rect 22621 -31864 22929 -31236
rect 23621 -31864 23929 -31236
rect 24621 -31864 24929 -31236
rect 25621 -31864 25929 -31236
rect 26621 -31864 26929 -31236
rect 27621 -31864 27929 -31236
rect 28621 -31864 28929 -31236
rect 29621 -31864 29929 -31236
rect 30621 -31864 30929 -31236
rect 31621 -31864 31929 -31236
rect 32621 -31864 32929 -31236
rect 33621 -31864 33929 -31236
rect -74819 -32204 -74511 -31896
rect -74447 -32172 -74203 -31928
rect -74139 -32204 -73511 -31896
rect -73447 -32172 -73203 -31928
rect -73139 -32204 -72511 -31896
rect -72447 -32172 -72203 -31928
rect -72139 -32204 -71511 -31896
rect -71447 -32172 -71203 -31928
rect -71139 -32204 -70511 -31896
rect -70447 -32172 -70203 -31928
rect -70139 -32204 -69511 -31896
rect -69447 -32172 -69203 -31928
rect -69139 -32204 -68511 -31896
rect -68447 -32172 -68203 -31928
rect -68139 -32204 -67511 -31896
rect -67447 -32172 -67203 -31928
rect -67139 -32204 -66511 -31896
rect -66447 -32172 -66203 -31928
rect -66139 -32204 -65511 -31896
rect -65447 -32172 -65203 -31928
rect -65139 -32204 -64511 -31896
rect -64447 -32172 -64203 -31928
rect -64139 -32204 -63511 -31896
rect -63447 -32172 -63203 -31928
rect -63139 -32204 -62511 -31896
rect -62447 -32172 -62203 -31928
rect -62139 -32204 -61511 -31896
rect -61447 -32172 -61203 -31928
rect -61139 -32204 -60511 -31896
rect -60447 -32172 -60203 -31928
rect -60139 -32204 -59511 -31896
rect -59447 -32172 -59203 -31928
rect -59139 -32204 -58511 -31896
rect -58447 -32172 -58203 -31928
rect -58139 -32204 -57511 -31896
rect -57447 -32172 -57203 -31928
rect -57139 -32204 -56511 -31896
rect -56447 -32172 -56203 -31928
rect -56139 -32204 -55511 -31896
rect -55447 -32172 -55203 -31928
rect -55139 -32204 -54511 -31896
rect -54447 -32172 -54203 -31928
rect -54139 -32204 -53511 -31896
rect -53447 -32172 -53203 -31928
rect -53139 -32204 -52511 -31896
rect -52447 -32172 -52203 -31928
rect -52139 -32204 -51511 -31896
rect -51447 -32172 -51203 -31928
rect -51139 -32204 -50511 -31896
rect -50447 -32172 -50203 -31928
rect -50139 -32204 -49511 -31896
rect -49447 -32172 -49203 -31928
rect -49139 -32204 -48831 -31896
rect 8281 -32204 8589 -31896
rect 8653 -32172 8897 -31928
rect 8961 -32204 9589 -31896
rect 9653 -32172 9897 -31928
rect 9961 -32204 10589 -31896
rect 10653 -32172 10897 -31928
rect 10961 -32204 11589 -31896
rect 11653 -32172 11897 -31928
rect 11961 -32204 12589 -31896
rect 12653 -32172 12897 -31928
rect 12961 -32204 13589 -31896
rect 13653 -32172 13897 -31928
rect 13961 -32204 14589 -31896
rect 14653 -32172 14897 -31928
rect 14961 -32204 15589 -31896
rect 15653 -32172 15897 -31928
rect 15961 -32204 16589 -31896
rect 16653 -32172 16897 -31928
rect 16961 -32204 17589 -31896
rect 17653 -32172 17897 -31928
rect 17961 -32204 18589 -31896
rect 18653 -32172 18897 -31928
rect 18961 -32204 19589 -31896
rect 19653 -32172 19897 -31928
rect 19961 -32204 20589 -31896
rect 20653 -32172 20897 -31928
rect 20961 -32204 21589 -31896
rect 21653 -32172 21897 -31928
rect 21961 -32204 22589 -31896
rect 22653 -32172 22897 -31928
rect 22961 -32204 23589 -31896
rect 23653 -32172 23897 -31928
rect 23961 -32204 24589 -31896
rect 24653 -32172 24897 -31928
rect 24961 -32204 25589 -31896
rect 25653 -32172 25897 -31928
rect 25961 -32204 26589 -31896
rect 26653 -32172 26897 -31928
rect 26961 -32204 27589 -31896
rect 27653 -32172 27897 -31928
rect 27961 -32204 28589 -31896
rect 28653 -32172 28897 -31928
rect 28961 -32204 29589 -31896
rect 29653 -32172 29897 -31928
rect 29961 -32204 30589 -31896
rect 30653 -32172 30897 -31928
rect 30961 -32204 31589 -31896
rect 31653 -32172 31897 -31928
rect 31961 -32204 32589 -31896
rect 32653 -32172 32897 -31928
rect 32961 -32204 33589 -31896
rect 33653 -32172 33897 -31928
rect 33961 -32204 34269 -31896
rect -74479 -32864 -74171 -32236
rect -73479 -32864 -73171 -32236
rect -72479 -32864 -72171 -32236
rect -71479 -32864 -71171 -32236
rect -70479 -32864 -70171 -32236
rect -69479 -32864 -69171 -32236
rect -68479 -32864 -68171 -32236
rect -67479 -32864 -67171 -32236
rect -66479 -32864 -66171 -32236
rect -65479 -32864 -65171 -32236
rect -64479 -32864 -64171 -32236
rect -63479 -32864 -63171 -32236
rect -62479 -32864 -62171 -32236
rect -61479 -32864 -61171 -32236
rect -60479 -32864 -60171 -32236
rect -59479 -32864 -59171 -32236
rect -58479 -32864 -58171 -32236
rect -57479 -32864 -57171 -32236
rect -56479 -32864 -56171 -32236
rect -55479 -32864 -55171 -32236
rect -54479 -32864 -54171 -32236
rect -53479 -32864 -53171 -32236
rect -52479 -32864 -52171 -32236
rect -51479 -32864 -51171 -32236
rect -50479 -32864 -50171 -32236
rect -49479 -32864 -49171 -32236
rect -74819 -33204 -74511 -32896
rect -74447 -33172 -74203 -32928
rect -74139 -33204 -73511 -32896
rect -73447 -33172 -73203 -32928
rect -73139 -33204 -72511 -32896
rect -72447 -33172 -72203 -32928
rect -72139 -33204 -71511 -32896
rect -71447 -33172 -71203 -32928
rect -71139 -33204 -70511 -32896
rect -70447 -33172 -70203 -32928
rect -70139 -33204 -69511 -32896
rect -69447 -33172 -69203 -32928
rect -69139 -33204 -68511 -32896
rect -68447 -33172 -68203 -32928
rect -68139 -33204 -67511 -32896
rect -67447 -33172 -67203 -32928
rect -67139 -33204 -66511 -32896
rect -66447 -33172 -66203 -32928
rect -66139 -33204 -65511 -32896
rect -65447 -33172 -65203 -32928
rect -65139 -33204 -64511 -32896
rect -64447 -33172 -64203 -32928
rect -64139 -33204 -63511 -32896
rect -63447 -33172 -63203 -32928
rect -63139 -33204 -62511 -32896
rect -62447 -33172 -62203 -32928
rect -62139 -33204 -61511 -32896
rect -61447 -33172 -61203 -32928
rect -61139 -33204 -60511 -32896
rect -60447 -33172 -60203 -32928
rect -60139 -33204 -59511 -32896
rect -59447 -33172 -59203 -32928
rect -59139 -33204 -58511 -32896
rect -58447 -33172 -58203 -32928
rect -58139 -33204 -57511 -32896
rect -57447 -33172 -57203 -32928
rect -57139 -33204 -56511 -32896
rect -56447 -33172 -56203 -32928
rect -56139 -33204 -55511 -32896
rect -55447 -33172 -55203 -32928
rect -55139 -33204 -54511 -32896
rect -54447 -33172 -54203 -32928
rect -54139 -33204 -53511 -32896
rect -53447 -33172 -53203 -32928
rect -53139 -33204 -52511 -32896
rect -52447 -33172 -52203 -32928
rect -52139 -33204 -51511 -32896
rect -51447 -33172 -51203 -32928
rect -51139 -33204 -50511 -32896
rect -50447 -33172 -50203 -32928
rect -50139 -33204 -49511 -32896
rect -49447 -33172 -49203 -32928
rect -49139 -33204 -48831 -32896
rect -74479 -33864 -74171 -33236
rect -73479 -33864 -73171 -33236
rect -72479 -33864 -72171 -33236
rect -71479 -33864 -71171 -33236
rect -70479 -33864 -70171 -33236
rect -69479 -33864 -69171 -33236
rect -68479 -33864 -68171 -33236
rect -67479 -33864 -67171 -33236
rect -66479 -33864 -66171 -33236
rect -65479 -33864 -65171 -33236
rect -64479 -33864 -64171 -33236
rect -63479 -33864 -63171 -33236
rect -62479 -33864 -62171 -33236
rect -61479 -33864 -61171 -33236
rect -60479 -33864 -60171 -33236
rect -59479 -33864 -59171 -33236
rect -58479 -33864 -58171 -33236
rect -57479 -33864 -57171 -33236
rect -56479 -33864 -56171 -33236
rect -55479 -33864 -55171 -33236
rect -54479 -33864 -54171 -33236
rect -53479 -33864 -53171 -33236
rect -52479 -33864 -52171 -33236
rect -51479 -33864 -51171 -33236
rect -50479 -33864 -50171 -33236
rect -49479 -33864 -49171 -33236
rect -74819 -34204 -74511 -33896
rect -74447 -34172 -74203 -33928
rect -74139 -34204 -73511 -33896
rect -73447 -34172 -73203 -33928
rect -73139 -34204 -72511 -33896
rect -72447 -34172 -72203 -33928
rect -72139 -34204 -71511 -33896
rect -71447 -34172 -71203 -33928
rect -71139 -34204 -70511 -33896
rect -70447 -34172 -70203 -33928
rect -70139 -34204 -69511 -33896
rect -69447 -34172 -69203 -33928
rect -69139 -34204 -68511 -33896
rect -68447 -34172 -68203 -33928
rect -68139 -34204 -67511 -33896
rect -67447 -34172 -67203 -33928
rect -67139 -34204 -66511 -33896
rect -66447 -34172 -66203 -33928
rect -66139 -34204 -65511 -33896
rect -65447 -34172 -65203 -33928
rect -65139 -34204 -64511 -33896
rect -64447 -34172 -64203 -33928
rect -64139 -34204 -63511 -33896
rect -63447 -34172 -63203 -33928
rect -63139 -34204 -62511 -33896
rect -62447 -34172 -62203 -33928
rect -62139 -34204 -61511 -33896
rect -61447 -34172 -61203 -33928
rect -61139 -34204 -60511 -33896
rect -60447 -34172 -60203 -33928
rect -60139 -34204 -59511 -33896
rect -59447 -34172 -59203 -33928
rect -59139 -34204 -58511 -33896
rect -58447 -34172 -58203 -33928
rect -58139 -34204 -57511 -33896
rect -57447 -34172 -57203 -33928
rect -57139 -34204 -56511 -33896
rect -56447 -34172 -56203 -33928
rect -56139 -34204 -55511 -33896
rect -55447 -34172 -55203 -33928
rect -55139 -34204 -54511 -33896
rect -54447 -34172 -54203 -33928
rect -54139 -34204 -53511 -33896
rect -53447 -34172 -53203 -33928
rect -53139 -34204 -52511 -33896
rect -52447 -34172 -52203 -33928
rect -52139 -34204 -51511 -33896
rect -51447 -34172 -51203 -33928
rect -51139 -34204 -50511 -33896
rect -50447 -34172 -50203 -33928
rect -50139 -34204 -49511 -33896
rect -49447 -34172 -49203 -33928
rect -49139 -34204 -48831 -33896
rect -74479 -34864 -74171 -34236
rect -73479 -34864 -73171 -34236
rect -72479 -34864 -72171 -34236
rect -71479 -34864 -71171 -34236
rect -70479 -34864 -70171 -34236
rect -69479 -34864 -69171 -34236
rect -68479 -34864 -68171 -34236
rect -67479 -34864 -67171 -34236
rect -66479 -34864 -66171 -34236
rect -65479 -34864 -65171 -34236
rect -64479 -34864 -64171 -34236
rect -63479 -34864 -63171 -34236
rect -62479 -34864 -62171 -34236
rect -61479 -34864 -61171 -34236
rect -60479 -34864 -60171 -34236
rect -59479 -34864 -59171 -34236
rect -58479 -34864 -58171 -34236
rect -57479 -34864 -57171 -34236
rect -56479 -34864 -56171 -34236
rect -55479 -34864 -55171 -34236
rect -54479 -34864 -54171 -34236
rect -53479 -34864 -53171 -34236
rect -52479 -34864 -52171 -34236
rect -51479 -34864 -51171 -34236
rect -50479 -34864 -50171 -34236
rect -49479 -34864 -49171 -34236
rect -74819 -35204 -74511 -34896
rect -74447 -35172 -74203 -34928
rect -74139 -35204 -73511 -34896
rect -73447 -35172 -73203 -34928
rect -73139 -35204 -72511 -34896
rect -72447 -35172 -72203 -34928
rect -72139 -35204 -71511 -34896
rect -71447 -35172 -71203 -34928
rect -71139 -35204 -70511 -34896
rect -70447 -35172 -70203 -34928
rect -70139 -35204 -69511 -34896
rect -69447 -35172 -69203 -34928
rect -69139 -35204 -68511 -34896
rect -68447 -35172 -68203 -34928
rect -68139 -35204 -67511 -34896
rect -67447 -35172 -67203 -34928
rect -67139 -35204 -66511 -34896
rect -66447 -35172 -66203 -34928
rect -66139 -35204 -65511 -34896
rect -65447 -35172 -65203 -34928
rect -65139 -35204 -64511 -34896
rect -64447 -35172 -64203 -34928
rect -64139 -35204 -63511 -34896
rect -63447 -35172 -63203 -34928
rect -63139 -35204 -62511 -34896
rect -62447 -35172 -62203 -34928
rect -62139 -35204 -61511 -34896
rect -61447 -35172 -61203 -34928
rect -61139 -35204 -60511 -34896
rect -60447 -35172 -60203 -34928
rect -60139 -35204 -59511 -34896
rect -59447 -35172 -59203 -34928
rect -59139 -35204 -58511 -34896
rect -58447 -35172 -58203 -34928
rect -58139 -35204 -57511 -34896
rect -57447 -35172 -57203 -34928
rect -57139 -35204 -56511 -34896
rect -56447 -35172 -56203 -34928
rect -56139 -35204 -55511 -34896
rect -55447 -35172 -55203 -34928
rect -55139 -35204 -54511 -34896
rect -54447 -35172 -54203 -34928
rect -54139 -35204 -53511 -34896
rect -53447 -35172 -53203 -34928
rect -53139 -35204 -52511 -34896
rect -52447 -35172 -52203 -34928
rect -52139 -35204 -51511 -34896
rect -51447 -35172 -51203 -34928
rect -51139 -35204 -50511 -34896
rect -50447 -35172 -50203 -34928
rect -50139 -35204 -49511 -34896
rect -49447 -35172 -49203 -34928
rect -49139 -35204 -48831 -34896
rect -74479 -35864 -74171 -35236
rect -73479 -35864 -73171 -35236
rect -72479 -35864 -72171 -35236
rect -71479 -35864 -71171 -35236
rect -70479 -35864 -70171 -35236
rect -69479 -35864 -69171 -35236
rect -68479 -35864 -68171 -35236
rect -67479 -35864 -67171 -35236
rect -66479 -35864 -66171 -35236
rect -65479 -35864 -65171 -35236
rect -64479 -35864 -64171 -35236
rect -63479 -35864 -63171 -35236
rect -62479 -35864 -62171 -35236
rect -61479 -35864 -61171 -35236
rect -60479 -35864 -60171 -35236
rect -59479 -35864 -59171 -35236
rect -58479 -35864 -58171 -35236
rect -57479 -35864 -57171 -35236
rect -56479 -35864 -56171 -35236
rect -55479 -35864 -55171 -35236
rect -54479 -35864 -54171 -35236
rect -53479 -35864 -53171 -35236
rect -52479 -35864 -52171 -35236
rect -51479 -35864 -51171 -35236
rect -50479 -35864 -50171 -35236
rect -49479 -35864 -49171 -35236
rect -74819 -36204 -74511 -35896
rect -74447 -36172 -74203 -35928
rect -74139 -36204 -73511 -35896
rect -73447 -36172 -73203 -35928
rect -73139 -36204 -72511 -35896
rect -72447 -36172 -72203 -35928
rect -72139 -36204 -71511 -35896
rect -71447 -36172 -71203 -35928
rect -71139 -36204 -70511 -35896
rect -70447 -36172 -70203 -35928
rect -70139 -36204 -69511 -35896
rect -69447 -36172 -69203 -35928
rect -69139 -36204 -68511 -35896
rect -68447 -36172 -68203 -35928
rect -68139 -36204 -67511 -35896
rect -67447 -36172 -67203 -35928
rect -67139 -36204 -66511 -35896
rect -66447 -36172 -66203 -35928
rect -66139 -36204 -65511 -35896
rect -65447 -36172 -65203 -35928
rect -65139 -36204 -64511 -35896
rect -64447 -36172 -64203 -35928
rect -64139 -36204 -63511 -35896
rect -63447 -36172 -63203 -35928
rect -63139 -36204 -62511 -35896
rect -62447 -36172 -62203 -35928
rect -62139 -36204 -61511 -35896
rect -61447 -36172 -61203 -35928
rect -61139 -36204 -60511 -35896
rect -60447 -36172 -60203 -35928
rect -60139 -36204 -59511 -35896
rect -59447 -36172 -59203 -35928
rect -59139 -36204 -58511 -35896
rect -58447 -36172 -58203 -35928
rect -58139 -36204 -57511 -35896
rect -57447 -36172 -57203 -35928
rect -57139 -36204 -56511 -35896
rect -56447 -36172 -56203 -35928
rect -56139 -36204 -55511 -35896
rect -55447 -36172 -55203 -35928
rect -55139 -36204 -54511 -35896
rect -54447 -36172 -54203 -35928
rect -54139 -36204 -53511 -35896
rect -53447 -36172 -53203 -35928
rect -53139 -36204 -52511 -35896
rect -52447 -36172 -52203 -35928
rect -52139 -36204 -51511 -35896
rect -51447 -36172 -51203 -35928
rect -51139 -36204 -50511 -35896
rect -50447 -36172 -50203 -35928
rect -50139 -36204 -49511 -35896
rect -49447 -36172 -49203 -35928
rect -49139 -36204 -48831 -35896
rect -74479 -36864 -74171 -36236
rect -73479 -36864 -73171 -36236
rect -72479 -36864 -72171 -36236
rect -71479 -36864 -71171 -36236
rect -70479 -36864 -70171 -36236
rect -69479 -36864 -69171 -36236
rect -68479 -36864 -68171 -36236
rect -67479 -36864 -67171 -36236
rect -66479 -36864 -66171 -36236
rect -65479 -36864 -65171 -36236
rect -64479 -36864 -64171 -36236
rect -63479 -36864 -63171 -36236
rect -62479 -36864 -62171 -36236
rect -61479 -36864 -61171 -36236
rect -60479 -36864 -60171 -36236
rect -59479 -36864 -59171 -36236
rect -58479 -36864 -58171 -36236
rect -57479 -36864 -57171 -36236
rect -56479 -36864 -56171 -36236
rect -55479 -36864 -55171 -36236
rect -54479 -36864 -54171 -36236
rect -53479 -36864 -53171 -36236
rect -52479 -36864 -52171 -36236
rect -51479 -36864 -51171 -36236
rect -50479 -36864 -50171 -36236
rect -49479 -36864 -49171 -36236
rect -74819 -37204 -74511 -36896
rect -74447 -37172 -74203 -36928
rect -74139 -37204 -73511 -36896
rect -73447 -37172 -73203 -36928
rect -73139 -37204 -72511 -36896
rect -72447 -37172 -72203 -36928
rect -72139 -37204 -71511 -36896
rect -71447 -37172 -71203 -36928
rect -71139 -37204 -70511 -36896
rect -70447 -37172 -70203 -36928
rect -70139 -37204 -69511 -36896
rect -69447 -37172 -69203 -36928
rect -69139 -37204 -68511 -36896
rect -68447 -37172 -68203 -36928
rect -68139 -37204 -67511 -36896
rect -67447 -37172 -67203 -36928
rect -67139 -37204 -66511 -36896
rect -66447 -37172 -66203 -36928
rect -66139 -37204 -65511 -36896
rect -65447 -37172 -65203 -36928
rect -65139 -37204 -64511 -36896
rect -64447 -37172 -64203 -36928
rect -64139 -37204 -63511 -36896
rect -63447 -37172 -63203 -36928
rect -63139 -37204 -62511 -36896
rect -62447 -37172 -62203 -36928
rect -62139 -37204 -61511 -36896
rect -61447 -37172 -61203 -36928
rect -61139 -37204 -60511 -36896
rect -60447 -37172 -60203 -36928
rect -60139 -37204 -59511 -36896
rect -59447 -37172 -59203 -36928
rect -59139 -37204 -58511 -36896
rect -58447 -37172 -58203 -36928
rect -58139 -37204 -57511 -36896
rect -57447 -37172 -57203 -36928
rect -57139 -37204 -56511 -36896
rect -56447 -37172 -56203 -36928
rect -56139 -37204 -55511 -36896
rect -55447 -37172 -55203 -36928
rect -55139 -37204 -54511 -36896
rect -54447 -37172 -54203 -36928
rect -54139 -37204 -53511 -36896
rect -53447 -37172 -53203 -36928
rect -53139 -37204 -52511 -36896
rect -52447 -37172 -52203 -36928
rect -52139 -37204 -51511 -36896
rect -51447 -37172 -51203 -36928
rect -51139 -37204 -50511 -36896
rect -50447 -37172 -50203 -36928
rect -50139 -37204 -49511 -36896
rect -49447 -37172 -49203 -36928
rect -49139 -37204 -48831 -36896
rect -74479 -37864 -74171 -37236
rect -73479 -37864 -73171 -37236
rect -72479 -37864 -72171 -37236
rect -71479 -37864 -71171 -37236
rect -70479 -37864 -70171 -37236
rect -69479 -37864 -69171 -37236
rect -68479 -37864 -68171 -37236
rect -67479 -37864 -67171 -37236
rect -66479 -37864 -66171 -37236
rect -65479 -37864 -65171 -37236
rect -64479 -37864 -64171 -37236
rect -63479 -37864 -63171 -37236
rect -62479 -37864 -62171 -37236
rect -61479 -37864 -61171 -37236
rect -60479 -37864 -60171 -37236
rect -59479 -37864 -59171 -37236
rect -58479 -37864 -58171 -37236
rect -57479 -37864 -57171 -37236
rect -56479 -37864 -56171 -37236
rect -55479 -37864 -55171 -37236
rect -54479 -37864 -54171 -37236
rect -53479 -37864 -53171 -37236
rect -52479 -37864 -52171 -37236
rect -51479 -37864 -51171 -37236
rect -50479 -37864 -50171 -37236
rect -49479 -37864 -49171 -37236
rect -74819 -38204 -74511 -37896
rect -74447 -38172 -74203 -37928
rect -74139 -38204 -73511 -37896
rect -73447 -38172 -73203 -37928
rect -73139 -38204 -72511 -37896
rect -72447 -38172 -72203 -37928
rect -72139 -38204 -71511 -37896
rect -71447 -38172 -71203 -37928
rect -71139 -38204 -70511 -37896
rect -70447 -38172 -70203 -37928
rect -70139 -38204 -69511 -37896
rect -69447 -38172 -69203 -37928
rect -69139 -38204 -68511 -37896
rect -68447 -38172 -68203 -37928
rect -68139 -38204 -67511 -37896
rect -67447 -38172 -67203 -37928
rect -67139 -38204 -66511 -37896
rect -66447 -38172 -66203 -37928
rect -66139 -38204 -65511 -37896
rect -65447 -38172 -65203 -37928
rect -65139 -38204 -64511 -37896
rect -64447 -38172 -64203 -37928
rect -64139 -38204 -63511 -37896
rect -63447 -38172 -63203 -37928
rect -63139 -38204 -62511 -37896
rect -62447 -38172 -62203 -37928
rect -62139 -38204 -61511 -37896
rect -61447 -38172 -61203 -37928
rect -61139 -38204 -60511 -37896
rect -60447 -38172 -60203 -37928
rect -60139 -38204 -59511 -37896
rect -59447 -38172 -59203 -37928
rect -59139 -38204 -58511 -37896
rect -58447 -38172 -58203 -37928
rect -58139 -38204 -57511 -37896
rect -57447 -38172 -57203 -37928
rect -57139 -38204 -56511 -37896
rect -56447 -38172 -56203 -37928
rect -56139 -38204 -55511 -37896
rect -55447 -38172 -55203 -37928
rect -55139 -38204 -54511 -37896
rect -54447 -38172 -54203 -37928
rect -54139 -38204 -53511 -37896
rect -53447 -38172 -53203 -37928
rect -53139 -38204 -52511 -37896
rect -52447 -38172 -52203 -37928
rect -52139 -38204 -51511 -37896
rect -51447 -38172 -51203 -37928
rect -51139 -38204 -50511 -37896
rect -50447 -38172 -50203 -37928
rect -50139 -38204 -49511 -37896
rect -49447 -38172 -49203 -37928
rect -49139 -38204 -48831 -37896
rect -74479 -38864 -74171 -38236
rect -73479 -38864 -73171 -38236
rect -72479 -38864 -72171 -38236
rect -71479 -38864 -71171 -38236
rect -70479 -38864 -70171 -38236
rect -69479 -38864 -69171 -38236
rect -68479 -38864 -68171 -38236
rect -67479 -38864 -67171 -38236
rect -66479 -38864 -66171 -38236
rect -65479 -38864 -65171 -38236
rect -64479 -38864 -64171 -38236
rect -63479 -38864 -63171 -38236
rect -62479 -38864 -62171 -38236
rect -61479 -38864 -61171 -38236
rect -60479 -38864 -60171 -38236
rect -59479 -38864 -59171 -38236
rect -58479 -38864 -58171 -38236
rect -57479 -38864 -57171 -38236
rect -56479 -38864 -56171 -38236
rect -55479 -38864 -55171 -38236
rect -54479 -38864 -54171 -38236
rect -53479 -38864 -53171 -38236
rect -52479 -38864 -52171 -38236
rect -51479 -38864 -51171 -38236
rect -50479 -38864 -50171 -38236
rect -49479 -38864 -49171 -38236
rect -74819 -39204 -74511 -38896
rect -74447 -39172 -74203 -38928
rect -74139 -39204 -73511 -38896
rect -73447 -39172 -73203 -38928
rect -73139 -39204 -72511 -38896
rect -72447 -39172 -72203 -38928
rect -72139 -39204 -71511 -38896
rect -71447 -39172 -71203 -38928
rect -71139 -39204 -70511 -38896
rect -70447 -39172 -70203 -38928
rect -70139 -39204 -69511 -38896
rect -69447 -39172 -69203 -38928
rect -69139 -39204 -68511 -38896
rect -68447 -39172 -68203 -38928
rect -68139 -39204 -67511 -38896
rect -67447 -39172 -67203 -38928
rect -67139 -39204 -66511 -38896
rect -66447 -39172 -66203 -38928
rect -66139 -39204 -65511 -38896
rect -65447 -39172 -65203 -38928
rect -65139 -39204 -64511 -38896
rect -64447 -39172 -64203 -38928
rect -64139 -39204 -63511 -38896
rect -63447 -39172 -63203 -38928
rect -63139 -39204 -62511 -38896
rect -62447 -39172 -62203 -38928
rect -62139 -39204 -61511 -38896
rect -61447 -39172 -61203 -38928
rect -61139 -39204 -60511 -38896
rect -60447 -39172 -60203 -38928
rect -60139 -39204 -59511 -38896
rect -59447 -39172 -59203 -38928
rect -59139 -39204 -58511 -38896
rect -58447 -39172 -58203 -38928
rect -58139 -39204 -57511 -38896
rect -57447 -39172 -57203 -38928
rect -57139 -39204 -56511 -38896
rect -56447 -39172 -56203 -38928
rect -56139 -39204 -55511 -38896
rect -55447 -39172 -55203 -38928
rect -55139 -39204 -54511 -38896
rect -54447 -39172 -54203 -38928
rect -54139 -39204 -53511 -38896
rect -53447 -39172 -53203 -38928
rect -53139 -39204 -52511 -38896
rect -52447 -39172 -52203 -38928
rect -52139 -39204 -51511 -38896
rect -51447 -39172 -51203 -38928
rect -51139 -39204 -50511 -38896
rect -50447 -39172 -50203 -38928
rect -50139 -39204 -49511 -38896
rect -49447 -39172 -49203 -38928
rect -49139 -39204 -48831 -38896
rect -74479 -39864 -74171 -39236
rect -73479 -39864 -73171 -39236
rect -72479 -39864 -72171 -39236
rect -71479 -39864 -71171 -39236
rect -70479 -39864 -70171 -39236
rect -69479 -39864 -69171 -39236
rect -68479 -39864 -68171 -39236
rect -67479 -39864 -67171 -39236
rect -66479 -39864 -66171 -39236
rect -65479 -39864 -65171 -39236
rect -64479 -39864 -64171 -39236
rect -63479 -39864 -63171 -39236
rect -62479 -39864 -62171 -39236
rect -61479 -39864 -61171 -39236
rect -60479 -39864 -60171 -39236
rect -59479 -39864 -59171 -39236
rect -58479 -39864 -58171 -39236
rect -57479 -39864 -57171 -39236
rect -56479 -39864 -56171 -39236
rect -55479 -39864 -55171 -39236
rect -54479 -39864 -54171 -39236
rect -53479 -39864 -53171 -39236
rect -52479 -39864 -52171 -39236
rect -51479 -39864 -51171 -39236
rect -50479 -39864 -50171 -39236
rect -49479 -39864 -49171 -39236
rect -74819 -40204 -74511 -39896
rect -74447 -40172 -74203 -39928
rect -74139 -40204 -73511 -39896
rect -73447 -40172 -73203 -39928
rect -73139 -40204 -72511 -39896
rect -72447 -40172 -72203 -39928
rect -72139 -40204 -71511 -39896
rect -71447 -40172 -71203 -39928
rect -71139 -40204 -70511 -39896
rect -70447 -40172 -70203 -39928
rect -70139 -40204 -69511 -39896
rect -69447 -40172 -69203 -39928
rect -69139 -40204 -68511 -39896
rect -68447 -40172 -68203 -39928
rect -68139 -40204 -67511 -39896
rect -67447 -40172 -67203 -39928
rect -67139 -40204 -66511 -39896
rect -66447 -40172 -66203 -39928
rect -66139 -40204 -65511 -39896
rect -65447 -40172 -65203 -39928
rect -65139 -40204 -64511 -39896
rect -64447 -40172 -64203 -39928
rect -64139 -40204 -63511 -39896
rect -63447 -40172 -63203 -39928
rect -63139 -40204 -62511 -39896
rect -62447 -40172 -62203 -39928
rect -62139 -40204 -61511 -39896
rect -61447 -40172 -61203 -39928
rect -61139 -40204 -60511 -39896
rect -60447 -40172 -60203 -39928
rect -60139 -40204 -59511 -39896
rect -59447 -40172 -59203 -39928
rect -59139 -40204 -58511 -39896
rect -58447 -40172 -58203 -39928
rect -58139 -40204 -57511 -39896
rect -57447 -40172 -57203 -39928
rect -57139 -40204 -56511 -39896
rect -56447 -40172 -56203 -39928
rect -56139 -40204 -55511 -39896
rect -55447 -40172 -55203 -39928
rect -55139 -40204 -54511 -39896
rect -54447 -40172 -54203 -39928
rect -54139 -40204 -53511 -39896
rect -53447 -40172 -53203 -39928
rect -53139 -40204 -52511 -39896
rect -52447 -40172 -52203 -39928
rect -52139 -40204 -51511 -39896
rect -51447 -40172 -51203 -39928
rect -51139 -40204 -50511 -39896
rect -50447 -40172 -50203 -39928
rect -50139 -40204 -49511 -39896
rect -49447 -40172 -49203 -39928
rect -49139 -40204 -48831 -39896
rect -74479 -40864 -74171 -40236
rect -73479 -40864 -73171 -40236
rect -72479 -40864 -72171 -40236
rect -71479 -40864 -71171 -40236
rect -70479 -40864 -70171 -40236
rect -69479 -40864 -69171 -40236
rect -68479 -40864 -68171 -40236
rect -67479 -40864 -67171 -40236
rect -66479 -40864 -66171 -40236
rect -65479 -40864 -65171 -40236
rect -64479 -40864 -64171 -40236
rect -63479 -40864 -63171 -40236
rect -62479 -40864 -62171 -40236
rect -61479 -40864 -61171 -40236
rect -60479 -40864 -60171 -40236
rect -59479 -40864 -59171 -40236
rect -58479 -40864 -58171 -40236
rect -57479 -40864 -57171 -40236
rect -56479 -40864 -56171 -40236
rect -55479 -40864 -55171 -40236
rect -54479 -40864 -54171 -40236
rect -53479 -40864 -53171 -40236
rect -52479 -40864 -52171 -40236
rect -51479 -40864 -51171 -40236
rect -50479 -40864 -50171 -40236
rect -49479 -40864 -49171 -40236
rect -74819 -41204 -74511 -40896
rect -74447 -41172 -74203 -40928
rect -74139 -41204 -73511 -40896
rect -73447 -41172 -73203 -40928
rect -73139 -41204 -72511 -40896
rect -72447 -41172 -72203 -40928
rect -72139 -41204 -71511 -40896
rect -71447 -41172 -71203 -40928
rect -71139 -41204 -70511 -40896
rect -70447 -41172 -70203 -40928
rect -70139 -41204 -69511 -40896
rect -69447 -41172 -69203 -40928
rect -69139 -41204 -68511 -40896
rect -68447 -41172 -68203 -40928
rect -68139 -41204 -67511 -40896
rect -67447 -41172 -67203 -40928
rect -67139 -41204 -66511 -40896
rect -66447 -41172 -66203 -40928
rect -66139 -41204 -65511 -40896
rect -65447 -41172 -65203 -40928
rect -65139 -41204 -64511 -40896
rect -64447 -41172 -64203 -40928
rect -64139 -41204 -63511 -40896
rect -63447 -41172 -63203 -40928
rect -63139 -41204 -62511 -40896
rect -62447 -41172 -62203 -40928
rect -62139 -41204 -61511 -40896
rect -61447 -41172 -61203 -40928
rect -61139 -41204 -60511 -40896
rect -60447 -41172 -60203 -40928
rect -60139 -41204 -59511 -40896
rect -59447 -41172 -59203 -40928
rect -59139 -41204 -58511 -40896
rect -58447 -41172 -58203 -40928
rect -58139 -41204 -57511 -40896
rect -57447 -41172 -57203 -40928
rect -57139 -41204 -56511 -40896
rect -56447 -41172 -56203 -40928
rect -56139 -41204 -55511 -40896
rect -55447 -41172 -55203 -40928
rect -55139 -41204 -54511 -40896
rect -54447 -41172 -54203 -40928
rect -54139 -41204 -53511 -40896
rect -53447 -41172 -53203 -40928
rect -53139 -41204 -52511 -40896
rect -52447 -41172 -52203 -40928
rect -52139 -41204 -51511 -40896
rect -51447 -41172 -51203 -40928
rect -51139 -41204 -50511 -40896
rect -50447 -41172 -50203 -40928
rect -50139 -41204 -49511 -40896
rect -49447 -41172 -49203 -40928
rect -49139 -41204 -48831 -40896
rect -74479 -41864 -74171 -41236
rect -73479 -41864 -73171 -41236
rect -72479 -41864 -72171 -41236
rect -71479 -41864 -71171 -41236
rect -70479 -41864 -70171 -41236
rect -69479 -41864 -69171 -41236
rect -68479 -41864 -68171 -41236
rect -67479 -41864 -67171 -41236
rect -66479 -41864 -66171 -41236
rect -65479 -41864 -65171 -41236
rect -64479 -41864 -64171 -41236
rect -63479 -41864 -63171 -41236
rect -62479 -41864 -62171 -41236
rect -61479 -41864 -61171 -41236
rect -60479 -41864 -60171 -41236
rect -59479 -41864 -59171 -41236
rect -58479 -41864 -58171 -41236
rect -57479 -41864 -57171 -41236
rect -56479 -41864 -56171 -41236
rect -55479 -41864 -55171 -41236
rect -54479 -41864 -54171 -41236
rect -53479 -41864 -53171 -41236
rect -52479 -41864 -52171 -41236
rect -51479 -41864 -51171 -41236
rect -50479 -41864 -50171 -41236
rect -49479 -41864 -49171 -41236
rect -74819 -42204 -74511 -41896
rect -74447 -42172 -74203 -41928
rect -74139 -42204 -73511 -41896
rect -73447 -42172 -73203 -41928
rect -73139 -42204 -72511 -41896
rect -72447 -42172 -72203 -41928
rect -72139 -42204 -71511 -41896
rect -71447 -42172 -71203 -41928
rect -71139 -42204 -70511 -41896
rect -70447 -42172 -70203 -41928
rect -70139 -42204 -69511 -41896
rect -69447 -42172 -69203 -41928
rect -69139 -42204 -68511 -41896
rect -68447 -42172 -68203 -41928
rect -68139 -42204 -67511 -41896
rect -67447 -42172 -67203 -41928
rect -67139 -42204 -66511 -41896
rect -66447 -42172 -66203 -41928
rect -66139 -42204 -65511 -41896
rect -65447 -42172 -65203 -41928
rect -65139 -42204 -64511 -41896
rect -64447 -42172 -64203 -41928
rect -64139 -42204 -63511 -41896
rect -63447 -42172 -63203 -41928
rect -63139 -42204 -62511 -41896
rect -62447 -42172 -62203 -41928
rect -62139 -42204 -61511 -41896
rect -61447 -42172 -61203 -41928
rect -61139 -42204 -60511 -41896
rect -60447 -42172 -60203 -41928
rect -60139 -42204 -59511 -41896
rect -59447 -42172 -59203 -41928
rect -59139 -42204 -58511 -41896
rect -58447 -42172 -58203 -41928
rect -58139 -42204 -57511 -41896
rect -57447 -42172 -57203 -41928
rect -57139 -42204 -56511 -41896
rect -56447 -42172 -56203 -41928
rect -56139 -42204 -55511 -41896
rect -55447 -42172 -55203 -41928
rect -55139 -42204 -54511 -41896
rect -54447 -42172 -54203 -41928
rect -54139 -42204 -53511 -41896
rect -53447 -42172 -53203 -41928
rect -53139 -42204 -52511 -41896
rect -52447 -42172 -52203 -41928
rect -52139 -42204 -51511 -41896
rect -51447 -42172 -51203 -41928
rect -51139 -42204 -50511 -41896
rect -50447 -42172 -50203 -41928
rect -50139 -42204 -49511 -41896
rect -49447 -42172 -49203 -41928
rect -49139 -42204 -48831 -41896
rect -74479 -42864 -74171 -42236
rect -73479 -42864 -73171 -42236
rect -72479 -42864 -72171 -42236
rect -71479 -42864 -71171 -42236
rect -70479 -42864 -70171 -42236
rect -69479 -42864 -69171 -42236
rect -68479 -42864 -68171 -42236
rect -67479 -42864 -67171 -42236
rect -66479 -42864 -66171 -42236
rect -65479 -42864 -65171 -42236
rect -64479 -42864 -64171 -42236
rect -63479 -42864 -63171 -42236
rect -62479 -42864 -62171 -42236
rect -61479 -42864 -61171 -42236
rect -60479 -42864 -60171 -42236
rect -59479 -42864 -59171 -42236
rect -58479 -42864 -58171 -42236
rect -57479 -42864 -57171 -42236
rect -56479 -42864 -56171 -42236
rect -55479 -42864 -55171 -42236
rect -54479 -42864 -54171 -42236
rect -53479 -42864 -53171 -42236
rect -52479 -42864 -52171 -42236
rect -51479 -42864 -51171 -42236
rect -50479 -42864 -50171 -42236
rect -49479 -42864 -49171 -42236
rect -74819 -43204 -74511 -42896
rect -74447 -43172 -74203 -42928
rect -74139 -43204 -73511 -42896
rect -73447 -43172 -73203 -42928
rect -73139 -43204 -72511 -42896
rect -72447 -43172 -72203 -42928
rect -72139 -43204 -71511 -42896
rect -71447 -43172 -71203 -42928
rect -71139 -43204 -70511 -42896
rect -70447 -43172 -70203 -42928
rect -70139 -43204 -69511 -42896
rect -69447 -43172 -69203 -42928
rect -69139 -43204 -68511 -42896
rect -68447 -43172 -68203 -42928
rect -68139 -43204 -67511 -42896
rect -67447 -43172 -67203 -42928
rect -67139 -43204 -66511 -42896
rect -66447 -43172 -66203 -42928
rect -66139 -43204 -65511 -42896
rect -65447 -43172 -65203 -42928
rect -65139 -43204 -64511 -42896
rect -64447 -43172 -64203 -42928
rect -64139 -43204 -63511 -42896
rect -63447 -43172 -63203 -42928
rect -63139 -43204 -62511 -42896
rect -62447 -43172 -62203 -42928
rect -62139 -43204 -61511 -42896
rect -61447 -43172 -61203 -42928
rect -61139 -43204 -60511 -42896
rect -60447 -43172 -60203 -42928
rect -60139 -43204 -59511 -42896
rect -59447 -43172 -59203 -42928
rect -59139 -43204 -58511 -42896
rect -58447 -43172 -58203 -42928
rect -58139 -43204 -57511 -42896
rect -57447 -43172 -57203 -42928
rect -57139 -43204 -56511 -42896
rect -56447 -43172 -56203 -42928
rect -56139 -43204 -55511 -42896
rect -55447 -43172 -55203 -42928
rect -55139 -43204 -54511 -42896
rect -54447 -43172 -54203 -42928
rect -54139 -43204 -53511 -42896
rect -53447 -43172 -53203 -42928
rect -53139 -43204 -52511 -42896
rect -52447 -43172 -52203 -42928
rect -52139 -43204 -51511 -42896
rect -51447 -43172 -51203 -42928
rect -51139 -43204 -50511 -42896
rect -50447 -43172 -50203 -42928
rect -50139 -43204 -49511 -42896
rect -49447 -43172 -49203 -42928
rect -49139 -43204 -48831 -42896
rect -74479 -43864 -74171 -43236
rect -73479 -43864 -73171 -43236
rect -72479 -43864 -72171 -43236
rect -71479 -43864 -71171 -43236
rect -70479 -43864 -70171 -43236
rect -69479 -43864 -69171 -43236
rect -68479 -43864 -68171 -43236
rect -67479 -43864 -67171 -43236
rect -66479 -43864 -66171 -43236
rect -65479 -43864 -65171 -43236
rect -64479 -43864 -64171 -43236
rect -63479 -43864 -63171 -43236
rect -62479 -43864 -62171 -43236
rect -61479 -43864 -61171 -43236
rect -60479 -43864 -60171 -43236
rect -59479 -43864 -59171 -43236
rect -58479 -43864 -58171 -43236
rect -57479 -43864 -57171 -43236
rect -56479 -43864 -56171 -43236
rect -55479 -43864 -55171 -43236
rect -54479 -43864 -54171 -43236
rect -53479 -43864 -53171 -43236
rect -52479 -43864 -52171 -43236
rect -51479 -43864 -51171 -43236
rect -50479 -43864 -50171 -43236
rect -49479 -43864 -49171 -43236
rect -74819 -44204 -74511 -43896
rect -74447 -44172 -74203 -43928
rect -74139 -44204 -73511 -43896
rect -73447 -44172 -73203 -43928
rect -73139 -44204 -72511 -43896
rect -72447 -44172 -72203 -43928
rect -72139 -44204 -71511 -43896
rect -71447 -44172 -71203 -43928
rect -71139 -44204 -70511 -43896
rect -70447 -44172 -70203 -43928
rect -70139 -44204 -69511 -43896
rect -69447 -44172 -69203 -43928
rect -69139 -44204 -68511 -43896
rect -68447 -44172 -68203 -43928
rect -68139 -44204 -67511 -43896
rect -67447 -44172 -67203 -43928
rect -67139 -44204 -66511 -43896
rect -66447 -44172 -66203 -43928
rect -66139 -44204 -65511 -43896
rect -65447 -44172 -65203 -43928
rect -65139 -44204 -64511 -43896
rect -64447 -44172 -64203 -43928
rect -64139 -44204 -63511 -43896
rect -63447 -44172 -63203 -43928
rect -63139 -44204 -62511 -43896
rect -62447 -44172 -62203 -43928
rect -62139 -44204 -61511 -43896
rect -61447 -44172 -61203 -43928
rect -61139 -44204 -60511 -43896
rect -60447 -44172 -60203 -43928
rect -60139 -44204 -59511 -43896
rect -59447 -44172 -59203 -43928
rect -59139 -44204 -58511 -43896
rect -58447 -44172 -58203 -43928
rect -58139 -44204 -57511 -43896
rect -57447 -44172 -57203 -43928
rect -57139 -44204 -56511 -43896
rect -56447 -44172 -56203 -43928
rect -56139 -44204 -55511 -43896
rect -55447 -44172 -55203 -43928
rect -55139 -44204 -54511 -43896
rect -54447 -44172 -54203 -43928
rect -54139 -44204 -53511 -43896
rect -53447 -44172 -53203 -43928
rect -53139 -44204 -52511 -43896
rect -52447 -44172 -52203 -43928
rect -52139 -44204 -51511 -43896
rect -51447 -44172 -51203 -43928
rect -51139 -44204 -50511 -43896
rect -50447 -44172 -50203 -43928
rect -50139 -44204 -49511 -43896
rect -49447 -44172 -49203 -43928
rect -49139 -44204 -48831 -43896
rect -74479 -44864 -74171 -44236
rect -73479 -44864 -73171 -44236
rect -72479 -44864 -72171 -44236
rect -71479 -44864 -71171 -44236
rect -70479 -44864 -70171 -44236
rect -69479 -44864 -69171 -44236
rect -68479 -44864 -68171 -44236
rect -67479 -44864 -67171 -44236
rect -66479 -44864 -66171 -44236
rect -65479 -44864 -65171 -44236
rect -64479 -44864 -64171 -44236
rect -63479 -44864 -63171 -44236
rect -62479 -44864 -62171 -44236
rect -61479 -44864 -61171 -44236
rect -60479 -44864 -60171 -44236
rect -59479 -44864 -59171 -44236
rect -58479 -44864 -58171 -44236
rect -57479 -44864 -57171 -44236
rect -56479 -44864 -56171 -44236
rect -55479 -44864 -55171 -44236
rect -54479 -44864 -54171 -44236
rect -53479 -44864 -53171 -44236
rect -52479 -44864 -52171 -44236
rect -51479 -44864 -51171 -44236
rect -50479 -44864 -50171 -44236
rect -49479 -44864 -49171 -44236
rect -46234 -44496 -36326 -32604
rect -4234 -44496 5674 -32604
rect 8621 -32864 8929 -32236
rect 9621 -32864 9929 -32236
rect 10621 -32864 10929 -32236
rect 11621 -32864 11929 -32236
rect 12621 -32864 12929 -32236
rect 13621 -32864 13929 -32236
rect 14621 -32864 14929 -32236
rect 15621 -32864 15929 -32236
rect 16621 -32864 16929 -32236
rect 17621 -32864 17929 -32236
rect 18621 -32864 18929 -32236
rect 19621 -32864 19929 -32236
rect 20621 -32864 20929 -32236
rect 21621 -32864 21929 -32236
rect 22621 -32864 22929 -32236
rect 23621 -32864 23929 -32236
rect 24621 -32864 24929 -32236
rect 25621 -32864 25929 -32236
rect 26621 -32864 26929 -32236
rect 27621 -32864 27929 -32236
rect 28621 -32864 28929 -32236
rect 29621 -32864 29929 -32236
rect 30621 -32864 30929 -32236
rect 31621 -32864 31929 -32236
rect 32621 -32864 32929 -32236
rect 33621 -32864 33929 -32236
rect 8281 -33204 8589 -32896
rect 8653 -33172 8897 -32928
rect 8961 -33204 9589 -32896
rect 9653 -33172 9897 -32928
rect 9961 -33204 10589 -32896
rect 10653 -33172 10897 -32928
rect 10961 -33204 11589 -32896
rect 11653 -33172 11897 -32928
rect 11961 -33204 12589 -32896
rect 12653 -33172 12897 -32928
rect 12961 -33204 13589 -32896
rect 13653 -33172 13897 -32928
rect 13961 -33204 14589 -32896
rect 14653 -33172 14897 -32928
rect 14961 -33204 15589 -32896
rect 15653 -33172 15897 -32928
rect 15961 -33204 16589 -32896
rect 16653 -33172 16897 -32928
rect 16961 -33204 17589 -32896
rect 17653 -33172 17897 -32928
rect 17961 -33204 18589 -32896
rect 18653 -33172 18897 -32928
rect 18961 -33204 19589 -32896
rect 19653 -33172 19897 -32928
rect 19961 -33204 20589 -32896
rect 20653 -33172 20897 -32928
rect 20961 -33204 21589 -32896
rect 21653 -33172 21897 -32928
rect 21961 -33204 22589 -32896
rect 22653 -33172 22897 -32928
rect 22961 -33204 23589 -32896
rect 23653 -33172 23897 -32928
rect 23961 -33204 24589 -32896
rect 24653 -33172 24897 -32928
rect 24961 -33204 25589 -32896
rect 25653 -33172 25897 -32928
rect 25961 -33204 26589 -32896
rect 26653 -33172 26897 -32928
rect 26961 -33204 27589 -32896
rect 27653 -33172 27897 -32928
rect 27961 -33204 28589 -32896
rect 28653 -33172 28897 -32928
rect 28961 -33204 29589 -32896
rect 29653 -33172 29897 -32928
rect 29961 -33204 30589 -32896
rect 30653 -33172 30897 -32928
rect 30961 -33204 31589 -32896
rect 31653 -33172 31897 -32928
rect 31961 -33204 32589 -32896
rect 32653 -33172 32897 -32928
rect 32961 -33204 33589 -32896
rect 33653 -33172 33897 -32928
rect 33961 -33204 34269 -32896
rect 8621 -33864 8929 -33236
rect 9621 -33864 9929 -33236
rect 10621 -33864 10929 -33236
rect 11621 -33864 11929 -33236
rect 12621 -33864 12929 -33236
rect 13621 -33864 13929 -33236
rect 14621 -33864 14929 -33236
rect 15621 -33864 15929 -33236
rect 16621 -33864 16929 -33236
rect 17621 -33864 17929 -33236
rect 18621 -33864 18929 -33236
rect 19621 -33864 19929 -33236
rect 20621 -33864 20929 -33236
rect 21621 -33864 21929 -33236
rect 22621 -33864 22929 -33236
rect 23621 -33864 23929 -33236
rect 24621 -33864 24929 -33236
rect 25621 -33864 25929 -33236
rect 26621 -33864 26929 -33236
rect 27621 -33864 27929 -33236
rect 28621 -33864 28929 -33236
rect 29621 -33864 29929 -33236
rect 30621 -33864 30929 -33236
rect 31621 -33864 31929 -33236
rect 32621 -33864 32929 -33236
rect 33621 -33864 33929 -33236
rect 8281 -34204 8589 -33896
rect 8653 -34172 8897 -33928
rect 8961 -34204 9589 -33896
rect 9653 -34172 9897 -33928
rect 9961 -34204 10589 -33896
rect 10653 -34172 10897 -33928
rect 10961 -34204 11589 -33896
rect 11653 -34172 11897 -33928
rect 11961 -34204 12589 -33896
rect 12653 -34172 12897 -33928
rect 12961 -34204 13589 -33896
rect 13653 -34172 13897 -33928
rect 13961 -34204 14589 -33896
rect 14653 -34172 14897 -33928
rect 14961 -34204 15589 -33896
rect 15653 -34172 15897 -33928
rect 15961 -34204 16589 -33896
rect 16653 -34172 16897 -33928
rect 16961 -34204 17589 -33896
rect 17653 -34172 17897 -33928
rect 17961 -34204 18589 -33896
rect 18653 -34172 18897 -33928
rect 18961 -34204 19589 -33896
rect 19653 -34172 19897 -33928
rect 19961 -34204 20589 -33896
rect 20653 -34172 20897 -33928
rect 20961 -34204 21589 -33896
rect 21653 -34172 21897 -33928
rect 21961 -34204 22589 -33896
rect 22653 -34172 22897 -33928
rect 22961 -34204 23589 -33896
rect 23653 -34172 23897 -33928
rect 23961 -34204 24589 -33896
rect 24653 -34172 24897 -33928
rect 24961 -34204 25589 -33896
rect 25653 -34172 25897 -33928
rect 25961 -34204 26589 -33896
rect 26653 -34172 26897 -33928
rect 26961 -34204 27589 -33896
rect 27653 -34172 27897 -33928
rect 27961 -34204 28589 -33896
rect 28653 -34172 28897 -33928
rect 28961 -34204 29589 -33896
rect 29653 -34172 29897 -33928
rect 29961 -34204 30589 -33896
rect 30653 -34172 30897 -33928
rect 30961 -34204 31589 -33896
rect 31653 -34172 31897 -33928
rect 31961 -34204 32589 -33896
rect 32653 -34172 32897 -33928
rect 32961 -34204 33589 -33896
rect 33653 -34172 33897 -33928
rect 33961 -34204 34269 -33896
rect 8621 -34864 8929 -34236
rect 9621 -34864 9929 -34236
rect 10621 -34864 10929 -34236
rect 11621 -34864 11929 -34236
rect 12621 -34864 12929 -34236
rect 13621 -34864 13929 -34236
rect 14621 -34864 14929 -34236
rect 15621 -34864 15929 -34236
rect 16621 -34864 16929 -34236
rect 17621 -34864 17929 -34236
rect 18621 -34864 18929 -34236
rect 19621 -34864 19929 -34236
rect 20621 -34864 20929 -34236
rect 21621 -34864 21929 -34236
rect 22621 -34864 22929 -34236
rect 23621 -34864 23929 -34236
rect 24621 -34864 24929 -34236
rect 25621 -34864 25929 -34236
rect 26621 -34864 26929 -34236
rect 27621 -34864 27929 -34236
rect 28621 -34864 28929 -34236
rect 29621 -34864 29929 -34236
rect 30621 -34864 30929 -34236
rect 31621 -34864 31929 -34236
rect 32621 -34864 32929 -34236
rect 33621 -34864 33929 -34236
rect 8281 -35204 8589 -34896
rect 8653 -35172 8897 -34928
rect 8961 -35204 9589 -34896
rect 9653 -35172 9897 -34928
rect 9961 -35204 10589 -34896
rect 10653 -35172 10897 -34928
rect 10961 -35204 11589 -34896
rect 11653 -35172 11897 -34928
rect 11961 -35204 12589 -34896
rect 12653 -35172 12897 -34928
rect 12961 -35204 13589 -34896
rect 13653 -35172 13897 -34928
rect 13961 -35204 14589 -34896
rect 14653 -35172 14897 -34928
rect 14961 -35204 15589 -34896
rect 15653 -35172 15897 -34928
rect 15961 -35204 16589 -34896
rect 16653 -35172 16897 -34928
rect 16961 -35204 17589 -34896
rect 17653 -35172 17897 -34928
rect 17961 -35204 18589 -34896
rect 18653 -35172 18897 -34928
rect 18961 -35204 19589 -34896
rect 19653 -35172 19897 -34928
rect 19961 -35204 20589 -34896
rect 20653 -35172 20897 -34928
rect 20961 -35204 21589 -34896
rect 21653 -35172 21897 -34928
rect 21961 -35204 22589 -34896
rect 22653 -35172 22897 -34928
rect 22961 -35204 23589 -34896
rect 23653 -35172 23897 -34928
rect 23961 -35204 24589 -34896
rect 24653 -35172 24897 -34928
rect 24961 -35204 25589 -34896
rect 25653 -35172 25897 -34928
rect 25961 -35204 26589 -34896
rect 26653 -35172 26897 -34928
rect 26961 -35204 27589 -34896
rect 27653 -35172 27897 -34928
rect 27961 -35204 28589 -34896
rect 28653 -35172 28897 -34928
rect 28961 -35204 29589 -34896
rect 29653 -35172 29897 -34928
rect 29961 -35204 30589 -34896
rect 30653 -35172 30897 -34928
rect 30961 -35204 31589 -34896
rect 31653 -35172 31897 -34928
rect 31961 -35204 32589 -34896
rect 32653 -35172 32897 -34928
rect 32961 -35204 33589 -34896
rect 33653 -35172 33897 -34928
rect 33961 -35204 34269 -34896
rect 8621 -35864 8929 -35236
rect 9621 -35864 9929 -35236
rect 10621 -35864 10929 -35236
rect 11621 -35864 11929 -35236
rect 12621 -35864 12929 -35236
rect 13621 -35864 13929 -35236
rect 14621 -35864 14929 -35236
rect 15621 -35864 15929 -35236
rect 16621 -35864 16929 -35236
rect 17621 -35864 17929 -35236
rect 18621 -35864 18929 -35236
rect 19621 -35864 19929 -35236
rect 20621 -35864 20929 -35236
rect 21621 -35864 21929 -35236
rect 22621 -35864 22929 -35236
rect 23621 -35864 23929 -35236
rect 24621 -35864 24929 -35236
rect 25621 -35864 25929 -35236
rect 26621 -35864 26929 -35236
rect 27621 -35864 27929 -35236
rect 28621 -35864 28929 -35236
rect 29621 -35864 29929 -35236
rect 30621 -35864 30929 -35236
rect 31621 -35864 31929 -35236
rect 32621 -35864 32929 -35236
rect 33621 -35864 33929 -35236
rect 8281 -36204 8589 -35896
rect 8653 -36172 8897 -35928
rect 8961 -36204 9589 -35896
rect 9653 -36172 9897 -35928
rect 9961 -36204 10589 -35896
rect 10653 -36172 10897 -35928
rect 10961 -36204 11589 -35896
rect 11653 -36172 11897 -35928
rect 11961 -36204 12589 -35896
rect 12653 -36172 12897 -35928
rect 12961 -36204 13589 -35896
rect 13653 -36172 13897 -35928
rect 13961 -36204 14589 -35896
rect 14653 -36172 14897 -35928
rect 14961 -36204 15589 -35896
rect 15653 -36172 15897 -35928
rect 15961 -36204 16589 -35896
rect 16653 -36172 16897 -35928
rect 16961 -36204 17589 -35896
rect 17653 -36172 17897 -35928
rect 17961 -36204 18589 -35896
rect 18653 -36172 18897 -35928
rect 18961 -36204 19589 -35896
rect 19653 -36172 19897 -35928
rect 19961 -36204 20589 -35896
rect 20653 -36172 20897 -35928
rect 20961 -36204 21589 -35896
rect 21653 -36172 21897 -35928
rect 21961 -36204 22589 -35896
rect 22653 -36172 22897 -35928
rect 22961 -36204 23589 -35896
rect 23653 -36172 23897 -35928
rect 23961 -36204 24589 -35896
rect 24653 -36172 24897 -35928
rect 24961 -36204 25589 -35896
rect 25653 -36172 25897 -35928
rect 25961 -36204 26589 -35896
rect 26653 -36172 26897 -35928
rect 26961 -36204 27589 -35896
rect 27653 -36172 27897 -35928
rect 27961 -36204 28589 -35896
rect 28653 -36172 28897 -35928
rect 28961 -36204 29589 -35896
rect 29653 -36172 29897 -35928
rect 29961 -36204 30589 -35896
rect 30653 -36172 30897 -35928
rect 30961 -36204 31589 -35896
rect 31653 -36172 31897 -35928
rect 31961 -36204 32589 -35896
rect 32653 -36172 32897 -35928
rect 32961 -36204 33589 -35896
rect 33653 -36172 33897 -35928
rect 33961 -36204 34269 -35896
rect 8621 -36864 8929 -36236
rect 9621 -36864 9929 -36236
rect 10621 -36864 10929 -36236
rect 11621 -36864 11929 -36236
rect 12621 -36864 12929 -36236
rect 13621 -36864 13929 -36236
rect 14621 -36864 14929 -36236
rect 15621 -36864 15929 -36236
rect 16621 -36864 16929 -36236
rect 17621 -36864 17929 -36236
rect 18621 -36864 18929 -36236
rect 19621 -36864 19929 -36236
rect 20621 -36864 20929 -36236
rect 21621 -36864 21929 -36236
rect 22621 -36864 22929 -36236
rect 23621 -36864 23929 -36236
rect 24621 -36864 24929 -36236
rect 25621 -36864 25929 -36236
rect 26621 -36864 26929 -36236
rect 27621 -36864 27929 -36236
rect 28621 -36864 28929 -36236
rect 29621 -36864 29929 -36236
rect 30621 -36864 30929 -36236
rect 31621 -36864 31929 -36236
rect 32621 -36864 32929 -36236
rect 33621 -36864 33929 -36236
rect 8281 -37204 8589 -36896
rect 8653 -37172 8897 -36928
rect 8961 -37204 9589 -36896
rect 9653 -37172 9897 -36928
rect 9961 -37204 10589 -36896
rect 10653 -37172 10897 -36928
rect 10961 -37204 11589 -36896
rect 11653 -37172 11897 -36928
rect 11961 -37204 12589 -36896
rect 12653 -37172 12897 -36928
rect 12961 -37204 13589 -36896
rect 13653 -37172 13897 -36928
rect 13961 -37204 14589 -36896
rect 14653 -37172 14897 -36928
rect 14961 -37204 15589 -36896
rect 15653 -37172 15897 -36928
rect 15961 -37204 16589 -36896
rect 16653 -37172 16897 -36928
rect 16961 -37204 17589 -36896
rect 17653 -37172 17897 -36928
rect 17961 -37204 18589 -36896
rect 18653 -37172 18897 -36928
rect 18961 -37204 19589 -36896
rect 19653 -37172 19897 -36928
rect 19961 -37204 20589 -36896
rect 20653 -37172 20897 -36928
rect 20961 -37204 21589 -36896
rect 21653 -37172 21897 -36928
rect 21961 -37204 22589 -36896
rect 22653 -37172 22897 -36928
rect 22961 -37204 23589 -36896
rect 23653 -37172 23897 -36928
rect 23961 -37204 24589 -36896
rect 24653 -37172 24897 -36928
rect 24961 -37204 25589 -36896
rect 25653 -37172 25897 -36928
rect 25961 -37204 26589 -36896
rect 26653 -37172 26897 -36928
rect 26961 -37204 27589 -36896
rect 27653 -37172 27897 -36928
rect 27961 -37204 28589 -36896
rect 28653 -37172 28897 -36928
rect 28961 -37204 29589 -36896
rect 29653 -37172 29897 -36928
rect 29961 -37204 30589 -36896
rect 30653 -37172 30897 -36928
rect 30961 -37204 31589 -36896
rect 31653 -37172 31897 -36928
rect 31961 -37204 32589 -36896
rect 32653 -37172 32897 -36928
rect 32961 -37204 33589 -36896
rect 33653 -37172 33897 -36928
rect 33961 -37204 34269 -36896
rect 8621 -37864 8929 -37236
rect 9621 -37864 9929 -37236
rect 10621 -37864 10929 -37236
rect 11621 -37864 11929 -37236
rect 12621 -37864 12929 -37236
rect 13621 -37864 13929 -37236
rect 14621 -37864 14929 -37236
rect 15621 -37864 15929 -37236
rect 16621 -37864 16929 -37236
rect 17621 -37864 17929 -37236
rect 18621 -37864 18929 -37236
rect 19621 -37864 19929 -37236
rect 20621 -37864 20929 -37236
rect 21621 -37864 21929 -37236
rect 22621 -37864 22929 -37236
rect 23621 -37864 23929 -37236
rect 24621 -37864 24929 -37236
rect 25621 -37864 25929 -37236
rect 26621 -37864 26929 -37236
rect 27621 -37864 27929 -37236
rect 28621 -37864 28929 -37236
rect 29621 -37864 29929 -37236
rect 30621 -37864 30929 -37236
rect 31621 -37864 31929 -37236
rect 32621 -37864 32929 -37236
rect 33621 -37864 33929 -37236
rect 8281 -38204 8589 -37896
rect 8653 -38172 8897 -37928
rect 8961 -38204 9589 -37896
rect 9653 -38172 9897 -37928
rect 9961 -38204 10589 -37896
rect 10653 -38172 10897 -37928
rect 10961 -38204 11589 -37896
rect 11653 -38172 11897 -37928
rect 11961 -38204 12589 -37896
rect 12653 -38172 12897 -37928
rect 12961 -38204 13589 -37896
rect 13653 -38172 13897 -37928
rect 13961 -38204 14589 -37896
rect 14653 -38172 14897 -37928
rect 14961 -38204 15589 -37896
rect 15653 -38172 15897 -37928
rect 15961 -38204 16589 -37896
rect 16653 -38172 16897 -37928
rect 16961 -38204 17589 -37896
rect 17653 -38172 17897 -37928
rect 17961 -38204 18589 -37896
rect 18653 -38172 18897 -37928
rect 18961 -38204 19589 -37896
rect 19653 -38172 19897 -37928
rect 19961 -38204 20589 -37896
rect 20653 -38172 20897 -37928
rect 20961 -38204 21589 -37896
rect 21653 -38172 21897 -37928
rect 21961 -38204 22589 -37896
rect 22653 -38172 22897 -37928
rect 22961 -38204 23589 -37896
rect 23653 -38172 23897 -37928
rect 23961 -38204 24589 -37896
rect 24653 -38172 24897 -37928
rect 24961 -38204 25589 -37896
rect 25653 -38172 25897 -37928
rect 25961 -38204 26589 -37896
rect 26653 -38172 26897 -37928
rect 26961 -38204 27589 -37896
rect 27653 -38172 27897 -37928
rect 27961 -38204 28589 -37896
rect 28653 -38172 28897 -37928
rect 28961 -38204 29589 -37896
rect 29653 -38172 29897 -37928
rect 29961 -38204 30589 -37896
rect 30653 -38172 30897 -37928
rect 30961 -38204 31589 -37896
rect 31653 -38172 31897 -37928
rect 31961 -38204 32589 -37896
rect 32653 -38172 32897 -37928
rect 32961 -38204 33589 -37896
rect 33653 -38172 33897 -37928
rect 33961 -38204 34269 -37896
rect 8621 -38864 8929 -38236
rect 9621 -38864 9929 -38236
rect 10621 -38864 10929 -38236
rect 11621 -38864 11929 -38236
rect 12621 -38864 12929 -38236
rect 13621 -38864 13929 -38236
rect 14621 -38864 14929 -38236
rect 15621 -38864 15929 -38236
rect 16621 -38864 16929 -38236
rect 17621 -38864 17929 -38236
rect 18621 -38864 18929 -38236
rect 19621 -38864 19929 -38236
rect 20621 -38864 20929 -38236
rect 21621 -38864 21929 -38236
rect 22621 -38864 22929 -38236
rect 23621 -38864 23929 -38236
rect 24621 -38864 24929 -38236
rect 25621 -38864 25929 -38236
rect 26621 -38864 26929 -38236
rect 27621 -38864 27929 -38236
rect 28621 -38864 28929 -38236
rect 29621 -38864 29929 -38236
rect 30621 -38864 30929 -38236
rect 31621 -38864 31929 -38236
rect 32621 -38864 32929 -38236
rect 33621 -38864 33929 -38236
rect 8281 -39204 8589 -38896
rect 8653 -39172 8897 -38928
rect 8961 -39204 9589 -38896
rect 9653 -39172 9897 -38928
rect 9961 -39204 10589 -38896
rect 10653 -39172 10897 -38928
rect 10961 -39204 11589 -38896
rect 11653 -39172 11897 -38928
rect 11961 -39204 12589 -38896
rect 12653 -39172 12897 -38928
rect 12961 -39204 13589 -38896
rect 13653 -39172 13897 -38928
rect 13961 -39204 14589 -38896
rect 14653 -39172 14897 -38928
rect 14961 -39204 15589 -38896
rect 15653 -39172 15897 -38928
rect 15961 -39204 16589 -38896
rect 16653 -39172 16897 -38928
rect 16961 -39204 17589 -38896
rect 17653 -39172 17897 -38928
rect 17961 -39204 18589 -38896
rect 18653 -39172 18897 -38928
rect 18961 -39204 19589 -38896
rect 19653 -39172 19897 -38928
rect 19961 -39204 20589 -38896
rect 20653 -39172 20897 -38928
rect 20961 -39204 21589 -38896
rect 21653 -39172 21897 -38928
rect 21961 -39204 22589 -38896
rect 22653 -39172 22897 -38928
rect 22961 -39204 23589 -38896
rect 23653 -39172 23897 -38928
rect 23961 -39204 24589 -38896
rect 24653 -39172 24897 -38928
rect 24961 -39204 25589 -38896
rect 25653 -39172 25897 -38928
rect 25961 -39204 26589 -38896
rect 26653 -39172 26897 -38928
rect 26961 -39204 27589 -38896
rect 27653 -39172 27897 -38928
rect 27961 -39204 28589 -38896
rect 28653 -39172 28897 -38928
rect 28961 -39204 29589 -38896
rect 29653 -39172 29897 -38928
rect 29961 -39204 30589 -38896
rect 30653 -39172 30897 -38928
rect 30961 -39204 31589 -38896
rect 31653 -39172 31897 -38928
rect 31961 -39204 32589 -38896
rect 32653 -39172 32897 -38928
rect 32961 -39204 33589 -38896
rect 33653 -39172 33897 -38928
rect 33961 -39204 34269 -38896
rect 8621 -39864 8929 -39236
rect 9621 -39864 9929 -39236
rect 10621 -39864 10929 -39236
rect 11621 -39864 11929 -39236
rect 12621 -39864 12929 -39236
rect 13621 -39864 13929 -39236
rect 14621 -39864 14929 -39236
rect 15621 -39864 15929 -39236
rect 16621 -39864 16929 -39236
rect 17621 -39864 17929 -39236
rect 18621 -39864 18929 -39236
rect 19621 -39864 19929 -39236
rect 20621 -39864 20929 -39236
rect 21621 -39864 21929 -39236
rect 22621 -39864 22929 -39236
rect 23621 -39864 23929 -39236
rect 24621 -39864 24929 -39236
rect 25621 -39864 25929 -39236
rect 26621 -39864 26929 -39236
rect 27621 -39864 27929 -39236
rect 28621 -39864 28929 -39236
rect 29621 -39864 29929 -39236
rect 30621 -39864 30929 -39236
rect 31621 -39864 31929 -39236
rect 32621 -39864 32929 -39236
rect 33621 -39864 33929 -39236
rect 8281 -40204 8589 -39896
rect 8653 -40172 8897 -39928
rect 8961 -40204 9589 -39896
rect 9653 -40172 9897 -39928
rect 9961 -40204 10589 -39896
rect 10653 -40172 10897 -39928
rect 10961 -40204 11589 -39896
rect 11653 -40172 11897 -39928
rect 11961 -40204 12589 -39896
rect 12653 -40172 12897 -39928
rect 12961 -40204 13589 -39896
rect 13653 -40172 13897 -39928
rect 13961 -40204 14589 -39896
rect 14653 -40172 14897 -39928
rect 14961 -40204 15589 -39896
rect 15653 -40172 15897 -39928
rect 15961 -40204 16589 -39896
rect 16653 -40172 16897 -39928
rect 16961 -40204 17589 -39896
rect 17653 -40172 17897 -39928
rect 17961 -40204 18589 -39896
rect 18653 -40172 18897 -39928
rect 18961 -40204 19589 -39896
rect 19653 -40172 19897 -39928
rect 19961 -40204 20589 -39896
rect 20653 -40172 20897 -39928
rect 20961 -40204 21589 -39896
rect 21653 -40172 21897 -39928
rect 21961 -40204 22589 -39896
rect 22653 -40172 22897 -39928
rect 22961 -40204 23589 -39896
rect 23653 -40172 23897 -39928
rect 23961 -40204 24589 -39896
rect 24653 -40172 24897 -39928
rect 24961 -40204 25589 -39896
rect 25653 -40172 25897 -39928
rect 25961 -40204 26589 -39896
rect 26653 -40172 26897 -39928
rect 26961 -40204 27589 -39896
rect 27653 -40172 27897 -39928
rect 27961 -40204 28589 -39896
rect 28653 -40172 28897 -39928
rect 28961 -40204 29589 -39896
rect 29653 -40172 29897 -39928
rect 29961 -40204 30589 -39896
rect 30653 -40172 30897 -39928
rect 30961 -40204 31589 -39896
rect 31653 -40172 31897 -39928
rect 31961 -40204 32589 -39896
rect 32653 -40172 32897 -39928
rect 32961 -40204 33589 -39896
rect 33653 -40172 33897 -39928
rect 33961 -40204 34269 -39896
rect 8621 -40864 8929 -40236
rect 9621 -40864 9929 -40236
rect 10621 -40864 10929 -40236
rect 11621 -40864 11929 -40236
rect 12621 -40864 12929 -40236
rect 13621 -40864 13929 -40236
rect 14621 -40864 14929 -40236
rect 15621 -40864 15929 -40236
rect 16621 -40864 16929 -40236
rect 17621 -40864 17929 -40236
rect 18621 -40864 18929 -40236
rect 19621 -40864 19929 -40236
rect 20621 -40864 20929 -40236
rect 21621 -40864 21929 -40236
rect 22621 -40864 22929 -40236
rect 23621 -40864 23929 -40236
rect 24621 -40864 24929 -40236
rect 25621 -40864 25929 -40236
rect 26621 -40864 26929 -40236
rect 27621 -40864 27929 -40236
rect 28621 -40864 28929 -40236
rect 29621 -40864 29929 -40236
rect 30621 -40864 30929 -40236
rect 31621 -40864 31929 -40236
rect 32621 -40864 32929 -40236
rect 33621 -40864 33929 -40236
rect 8281 -41204 8589 -40896
rect 8653 -41172 8897 -40928
rect 8961 -41204 9589 -40896
rect 9653 -41172 9897 -40928
rect 9961 -41204 10589 -40896
rect 10653 -41172 10897 -40928
rect 10961 -41204 11589 -40896
rect 11653 -41172 11897 -40928
rect 11961 -41204 12589 -40896
rect 12653 -41172 12897 -40928
rect 12961 -41204 13589 -40896
rect 13653 -41172 13897 -40928
rect 13961 -41204 14589 -40896
rect 14653 -41172 14897 -40928
rect 14961 -41204 15589 -40896
rect 15653 -41172 15897 -40928
rect 15961 -41204 16589 -40896
rect 16653 -41172 16897 -40928
rect 16961 -41204 17589 -40896
rect 17653 -41172 17897 -40928
rect 17961 -41204 18589 -40896
rect 18653 -41172 18897 -40928
rect 18961 -41204 19589 -40896
rect 19653 -41172 19897 -40928
rect 19961 -41204 20589 -40896
rect 20653 -41172 20897 -40928
rect 20961 -41204 21589 -40896
rect 21653 -41172 21897 -40928
rect 21961 -41204 22589 -40896
rect 22653 -41172 22897 -40928
rect 22961 -41204 23589 -40896
rect 23653 -41172 23897 -40928
rect 23961 -41204 24589 -40896
rect 24653 -41172 24897 -40928
rect 24961 -41204 25589 -40896
rect 25653 -41172 25897 -40928
rect 25961 -41204 26589 -40896
rect 26653 -41172 26897 -40928
rect 26961 -41204 27589 -40896
rect 27653 -41172 27897 -40928
rect 27961 -41204 28589 -40896
rect 28653 -41172 28897 -40928
rect 28961 -41204 29589 -40896
rect 29653 -41172 29897 -40928
rect 29961 -41204 30589 -40896
rect 30653 -41172 30897 -40928
rect 30961 -41204 31589 -40896
rect 31653 -41172 31897 -40928
rect 31961 -41204 32589 -40896
rect 32653 -41172 32897 -40928
rect 32961 -41204 33589 -40896
rect 33653 -41172 33897 -40928
rect 33961 -41204 34269 -40896
rect 8621 -41864 8929 -41236
rect 9621 -41864 9929 -41236
rect 10621 -41864 10929 -41236
rect 11621 -41864 11929 -41236
rect 12621 -41864 12929 -41236
rect 13621 -41864 13929 -41236
rect 14621 -41864 14929 -41236
rect 15621 -41864 15929 -41236
rect 16621 -41864 16929 -41236
rect 17621 -41864 17929 -41236
rect 18621 -41864 18929 -41236
rect 19621 -41864 19929 -41236
rect 20621 -41864 20929 -41236
rect 21621 -41864 21929 -41236
rect 22621 -41864 22929 -41236
rect 23621 -41864 23929 -41236
rect 24621 -41864 24929 -41236
rect 25621 -41864 25929 -41236
rect 26621 -41864 26929 -41236
rect 27621 -41864 27929 -41236
rect 28621 -41864 28929 -41236
rect 29621 -41864 29929 -41236
rect 30621 -41864 30929 -41236
rect 31621 -41864 31929 -41236
rect 32621 -41864 32929 -41236
rect 33621 -41864 33929 -41236
rect 8281 -42204 8589 -41896
rect 8653 -42172 8897 -41928
rect 8961 -42204 9589 -41896
rect 9653 -42172 9897 -41928
rect 9961 -42204 10589 -41896
rect 10653 -42172 10897 -41928
rect 10961 -42204 11589 -41896
rect 11653 -42172 11897 -41928
rect 11961 -42204 12589 -41896
rect 12653 -42172 12897 -41928
rect 12961 -42204 13589 -41896
rect 13653 -42172 13897 -41928
rect 13961 -42204 14589 -41896
rect 14653 -42172 14897 -41928
rect 14961 -42204 15589 -41896
rect 15653 -42172 15897 -41928
rect 15961 -42204 16589 -41896
rect 16653 -42172 16897 -41928
rect 16961 -42204 17589 -41896
rect 17653 -42172 17897 -41928
rect 17961 -42204 18589 -41896
rect 18653 -42172 18897 -41928
rect 18961 -42204 19589 -41896
rect 19653 -42172 19897 -41928
rect 19961 -42204 20589 -41896
rect 20653 -42172 20897 -41928
rect 20961 -42204 21589 -41896
rect 21653 -42172 21897 -41928
rect 21961 -42204 22589 -41896
rect 22653 -42172 22897 -41928
rect 22961 -42204 23589 -41896
rect 23653 -42172 23897 -41928
rect 23961 -42204 24589 -41896
rect 24653 -42172 24897 -41928
rect 24961 -42204 25589 -41896
rect 25653 -42172 25897 -41928
rect 25961 -42204 26589 -41896
rect 26653 -42172 26897 -41928
rect 26961 -42204 27589 -41896
rect 27653 -42172 27897 -41928
rect 27961 -42204 28589 -41896
rect 28653 -42172 28897 -41928
rect 28961 -42204 29589 -41896
rect 29653 -42172 29897 -41928
rect 29961 -42204 30589 -41896
rect 30653 -42172 30897 -41928
rect 30961 -42204 31589 -41896
rect 31653 -42172 31897 -41928
rect 31961 -42204 32589 -41896
rect 32653 -42172 32897 -41928
rect 32961 -42204 33589 -41896
rect 33653 -42172 33897 -41928
rect 33961 -42204 34269 -41896
rect 8621 -42864 8929 -42236
rect 9621 -42864 9929 -42236
rect 10621 -42864 10929 -42236
rect 11621 -42864 11929 -42236
rect 12621 -42864 12929 -42236
rect 13621 -42864 13929 -42236
rect 14621 -42864 14929 -42236
rect 15621 -42864 15929 -42236
rect 16621 -42864 16929 -42236
rect 17621 -42864 17929 -42236
rect 18621 -42864 18929 -42236
rect 19621 -42864 19929 -42236
rect 20621 -42864 20929 -42236
rect 21621 -42864 21929 -42236
rect 22621 -42864 22929 -42236
rect 23621 -42864 23929 -42236
rect 24621 -42864 24929 -42236
rect 25621 -42864 25929 -42236
rect 26621 -42864 26929 -42236
rect 27621 -42864 27929 -42236
rect 28621 -42864 28929 -42236
rect 29621 -42864 29929 -42236
rect 30621 -42864 30929 -42236
rect 31621 -42864 31929 -42236
rect 32621 -42864 32929 -42236
rect 33621 -42864 33929 -42236
rect 8281 -43204 8589 -42896
rect 8653 -43172 8897 -42928
rect 8961 -43204 9589 -42896
rect 9653 -43172 9897 -42928
rect 9961 -43204 10589 -42896
rect 10653 -43172 10897 -42928
rect 10961 -43204 11589 -42896
rect 11653 -43172 11897 -42928
rect 11961 -43204 12589 -42896
rect 12653 -43172 12897 -42928
rect 12961 -43204 13589 -42896
rect 13653 -43172 13897 -42928
rect 13961 -43204 14589 -42896
rect 14653 -43172 14897 -42928
rect 14961 -43204 15589 -42896
rect 15653 -43172 15897 -42928
rect 15961 -43204 16589 -42896
rect 16653 -43172 16897 -42928
rect 16961 -43204 17589 -42896
rect 17653 -43172 17897 -42928
rect 17961 -43204 18589 -42896
rect 18653 -43172 18897 -42928
rect 18961 -43204 19589 -42896
rect 19653 -43172 19897 -42928
rect 19961 -43204 20589 -42896
rect 20653 -43172 20897 -42928
rect 20961 -43204 21589 -42896
rect 21653 -43172 21897 -42928
rect 21961 -43204 22589 -42896
rect 22653 -43172 22897 -42928
rect 22961 -43204 23589 -42896
rect 23653 -43172 23897 -42928
rect 23961 -43204 24589 -42896
rect 24653 -43172 24897 -42928
rect 24961 -43204 25589 -42896
rect 25653 -43172 25897 -42928
rect 25961 -43204 26589 -42896
rect 26653 -43172 26897 -42928
rect 26961 -43204 27589 -42896
rect 27653 -43172 27897 -42928
rect 27961 -43204 28589 -42896
rect 28653 -43172 28897 -42928
rect 28961 -43204 29589 -42896
rect 29653 -43172 29897 -42928
rect 29961 -43204 30589 -42896
rect 30653 -43172 30897 -42928
rect 30961 -43204 31589 -42896
rect 31653 -43172 31897 -42928
rect 31961 -43204 32589 -42896
rect 32653 -43172 32897 -42928
rect 32961 -43204 33589 -42896
rect 33653 -43172 33897 -42928
rect 33961 -43204 34269 -42896
rect 8621 -43864 8929 -43236
rect 9621 -43864 9929 -43236
rect 10621 -43864 10929 -43236
rect 11621 -43864 11929 -43236
rect 12621 -43864 12929 -43236
rect 13621 -43864 13929 -43236
rect 14621 -43864 14929 -43236
rect 15621 -43864 15929 -43236
rect 16621 -43864 16929 -43236
rect 17621 -43864 17929 -43236
rect 18621 -43864 18929 -43236
rect 19621 -43864 19929 -43236
rect 20621 -43864 20929 -43236
rect 21621 -43864 21929 -43236
rect 22621 -43864 22929 -43236
rect 23621 -43864 23929 -43236
rect 24621 -43864 24929 -43236
rect 25621 -43864 25929 -43236
rect 26621 -43864 26929 -43236
rect 27621 -43864 27929 -43236
rect 28621 -43864 28929 -43236
rect 29621 -43864 29929 -43236
rect 30621 -43864 30929 -43236
rect 31621 -43864 31929 -43236
rect 32621 -43864 32929 -43236
rect 33621 -43864 33929 -43236
rect 8281 -44204 8589 -43896
rect 8653 -44172 8897 -43928
rect 8961 -44204 9589 -43896
rect 9653 -44172 9897 -43928
rect 9961 -44204 10589 -43896
rect 10653 -44172 10897 -43928
rect 10961 -44204 11589 -43896
rect 11653 -44172 11897 -43928
rect 11961 -44204 12589 -43896
rect 12653 -44172 12897 -43928
rect 12961 -44204 13589 -43896
rect 13653 -44172 13897 -43928
rect 13961 -44204 14589 -43896
rect 14653 -44172 14897 -43928
rect 14961 -44204 15589 -43896
rect 15653 -44172 15897 -43928
rect 15961 -44204 16589 -43896
rect 16653 -44172 16897 -43928
rect 16961 -44204 17589 -43896
rect 17653 -44172 17897 -43928
rect 17961 -44204 18589 -43896
rect 18653 -44172 18897 -43928
rect 18961 -44204 19589 -43896
rect 19653 -44172 19897 -43928
rect 19961 -44204 20589 -43896
rect 20653 -44172 20897 -43928
rect 20961 -44204 21589 -43896
rect 21653 -44172 21897 -43928
rect 21961 -44204 22589 -43896
rect 22653 -44172 22897 -43928
rect 22961 -44204 23589 -43896
rect 23653 -44172 23897 -43928
rect 23961 -44204 24589 -43896
rect 24653 -44172 24897 -43928
rect 24961 -44204 25589 -43896
rect 25653 -44172 25897 -43928
rect 25961 -44204 26589 -43896
rect 26653 -44172 26897 -43928
rect 26961 -44204 27589 -43896
rect 27653 -44172 27897 -43928
rect 27961 -44204 28589 -43896
rect 28653 -44172 28897 -43928
rect 28961 -44204 29589 -43896
rect 29653 -44172 29897 -43928
rect 29961 -44204 30589 -43896
rect 30653 -44172 30897 -43928
rect 30961 -44204 31589 -43896
rect 31653 -44172 31897 -43928
rect 31961 -44204 32589 -43896
rect 32653 -44172 32897 -43928
rect 32961 -44204 33589 -43896
rect 33653 -44172 33897 -43928
rect 33961 -44204 34269 -43896
rect 8621 -44864 8929 -44236
rect 9621 -44864 9929 -44236
rect 10621 -44864 10929 -44236
rect 11621 -44864 11929 -44236
rect 12621 -44864 12929 -44236
rect 13621 -44864 13929 -44236
rect 14621 -44864 14929 -44236
rect 15621 -44864 15929 -44236
rect 16621 -44864 16929 -44236
rect 17621 -44864 17929 -44236
rect 18621 -44864 18929 -44236
rect 19621 -44864 19929 -44236
rect 20621 -44864 20929 -44236
rect 21621 -44864 21929 -44236
rect 22621 -44864 22929 -44236
rect 23621 -44864 23929 -44236
rect 24621 -44864 24929 -44236
rect 25621 -44864 25929 -44236
rect 26621 -44864 26929 -44236
rect 27621 -44864 27929 -44236
rect 28621 -44864 28929 -44236
rect 29621 -44864 29929 -44236
rect 30621 -44864 30929 -44236
rect 31621 -44864 31929 -44236
rect 32621 -44864 32929 -44236
rect 33621 -44864 33929 -44236
rect -74819 -45204 -74511 -44896
rect -74447 -45172 -74203 -44928
rect -74139 -45204 -73511 -44896
rect -73447 -45172 -73203 -44928
rect -73139 -45204 -72511 -44896
rect -72447 -45172 -72203 -44928
rect -72139 -45204 -71511 -44896
rect -71447 -45172 -71203 -44928
rect -71139 -45204 -70511 -44896
rect -70447 -45172 -70203 -44928
rect -70139 -45204 -69511 -44896
rect -69447 -45172 -69203 -44928
rect -69139 -45204 -68511 -44896
rect -68447 -45172 -68203 -44928
rect -68139 -45204 -67511 -44896
rect -67447 -45172 -67203 -44928
rect -67139 -45204 -66511 -44896
rect -66447 -45172 -66203 -44928
rect -66139 -45204 -65511 -44896
rect -65447 -45172 -65203 -44928
rect -65139 -45204 -64511 -44896
rect -64447 -45172 -64203 -44928
rect -64139 -45204 -63511 -44896
rect -63447 -45172 -63203 -44928
rect -63139 -45204 -62511 -44896
rect -62447 -45172 -62203 -44928
rect -62139 -45204 -61511 -44896
rect -61447 -45172 -61203 -44928
rect -61139 -45204 -60511 -44896
rect -60447 -45172 -60203 -44928
rect -60139 -45204 -59511 -44896
rect -59447 -45172 -59203 -44928
rect -59139 -45204 -58511 -44896
rect -58447 -45172 -58203 -44928
rect -58139 -45204 -57511 -44896
rect -57447 -45172 -57203 -44928
rect -57139 -45204 -56511 -44896
rect -56447 -45172 -56203 -44928
rect -56139 -45204 -55511 -44896
rect -55447 -45172 -55203 -44928
rect -55139 -45204 -54511 -44896
rect -54447 -45172 -54203 -44928
rect -54139 -45204 -53511 -44896
rect -53447 -45172 -53203 -44928
rect -53139 -45204 -52511 -44896
rect -52447 -45172 -52203 -44928
rect -52139 -45204 -51511 -44896
rect -51447 -45172 -51203 -44928
rect -51139 -45204 -50511 -44896
rect -50447 -45172 -50203 -44928
rect -50139 -45204 -49511 -44896
rect -49447 -45172 -49203 -44928
rect -49139 -45204 -48831 -44896
rect 8281 -45204 8589 -44896
rect 8653 -45172 8897 -44928
rect 8961 -45204 9589 -44896
rect 9653 -45172 9897 -44928
rect 9961 -45204 10589 -44896
rect 10653 -45172 10897 -44928
rect 10961 -45204 11589 -44896
rect 11653 -45172 11897 -44928
rect 11961 -45204 12589 -44896
rect 12653 -45172 12897 -44928
rect 12961 -45204 13589 -44896
rect 13653 -45172 13897 -44928
rect 13961 -45204 14589 -44896
rect 14653 -45172 14897 -44928
rect 14961 -45204 15589 -44896
rect 15653 -45172 15897 -44928
rect 15961 -45204 16589 -44896
rect 16653 -45172 16897 -44928
rect 16961 -45204 17589 -44896
rect 17653 -45172 17897 -44928
rect 17961 -45204 18589 -44896
rect 18653 -45172 18897 -44928
rect 18961 -45204 19589 -44896
rect 19653 -45172 19897 -44928
rect 19961 -45204 20589 -44896
rect 20653 -45172 20897 -44928
rect 20961 -45204 21589 -44896
rect 21653 -45172 21897 -44928
rect 21961 -45204 22589 -44896
rect 22653 -45172 22897 -44928
rect 22961 -45204 23589 -44896
rect 23653 -45172 23897 -44928
rect 23961 -45204 24589 -44896
rect 24653 -45172 24897 -44928
rect 24961 -45204 25589 -44896
rect 25653 -45172 25897 -44928
rect 25961 -45204 26589 -44896
rect 26653 -45172 26897 -44928
rect 26961 -45204 27589 -44896
rect 27653 -45172 27897 -44928
rect 27961 -45204 28589 -44896
rect 28653 -45172 28897 -44928
rect 28961 -45204 29589 -44896
rect 29653 -45172 29897 -44928
rect 29961 -45204 30589 -44896
rect 30653 -45172 30897 -44928
rect 30961 -45204 31589 -44896
rect 31653 -45172 31897 -44928
rect 31961 -45204 32589 -44896
rect 32653 -45172 32897 -44928
rect 32961 -45204 33589 -44896
rect 33653 -45172 33897 -44928
rect 33961 -45204 34269 -44896
rect -74479 -45864 -74171 -45236
rect -73479 -45864 -73171 -45236
rect -72479 -45864 -72171 -45236
rect -71479 -45864 -71171 -45236
rect -70479 -45864 -70171 -45236
rect -69479 -45864 -69171 -45236
rect -68479 -45864 -68171 -45236
rect -67479 -45864 -67171 -45236
rect -66479 -45864 -66171 -45236
rect -65479 -45864 -65171 -45236
rect -64479 -45864 -64171 -45236
rect -63479 -45864 -63171 -45236
rect -62479 -45864 -62171 -45236
rect -61479 -45864 -61171 -45236
rect -60479 -45864 -60171 -45236
rect -59479 -45864 -59171 -45236
rect -58479 -45864 -58171 -45236
rect -57479 -45864 -57171 -45236
rect -56479 -45864 -56171 -45236
rect -55479 -45864 -55171 -45236
rect -54479 -45864 -54171 -45236
rect -53479 -45864 -53171 -45236
rect -52479 -45864 -52171 -45236
rect -51479 -45864 -51171 -45236
rect -50479 -45864 -50171 -45236
rect -49479 -45864 -49171 -45236
rect 8621 -45864 8929 -45236
rect 9621 -45864 9929 -45236
rect 10621 -45864 10929 -45236
rect 11621 -45864 11929 -45236
rect 12621 -45864 12929 -45236
rect 13621 -45864 13929 -45236
rect 14621 -45864 14929 -45236
rect 15621 -45864 15929 -45236
rect 16621 -45864 16929 -45236
rect 17621 -45864 17929 -45236
rect 18621 -45864 18929 -45236
rect 19621 -45864 19929 -45236
rect 20621 -45864 20929 -45236
rect 21621 -45864 21929 -45236
rect 22621 -45864 22929 -45236
rect 23621 -45864 23929 -45236
rect 24621 -45864 24929 -45236
rect 25621 -45864 25929 -45236
rect 26621 -45864 26929 -45236
rect 27621 -45864 27929 -45236
rect 28621 -45864 28929 -45236
rect 29621 -45864 29929 -45236
rect 30621 -45864 30929 -45236
rect 31621 -45864 31929 -45236
rect 32621 -45864 32929 -45236
rect 33621 -45864 33929 -45236
rect -74819 -46204 -74511 -45896
rect -74447 -46172 -74203 -45928
rect -74139 -46204 -73511 -45896
rect -73447 -46172 -73203 -45928
rect -73139 -46204 -72511 -45896
rect -72447 -46172 -72203 -45928
rect -72139 -46204 -71511 -45896
rect -71447 -46172 -71203 -45928
rect -71139 -46204 -70511 -45896
rect -70447 -46172 -70203 -45928
rect -70139 -46204 -69511 -45896
rect -69447 -46172 -69203 -45928
rect -69139 -46204 -68511 -45896
rect -68447 -46172 -68203 -45928
rect -68139 -46204 -67511 -45896
rect -67447 -46172 -67203 -45928
rect -67139 -46204 -66511 -45896
rect -66447 -46172 -66203 -45928
rect -66139 -46204 -65511 -45896
rect -65447 -46172 -65203 -45928
rect -65139 -46204 -64511 -45896
rect -64447 -46172 -64203 -45928
rect -64139 -46204 -63511 -45896
rect -63447 -46172 -63203 -45928
rect -63139 -46204 -62511 -45896
rect -62447 -46172 -62203 -45928
rect -62139 -46204 -61511 -45896
rect -61447 -46172 -61203 -45928
rect -61139 -46204 -60511 -45896
rect -60447 -46172 -60203 -45928
rect -60139 -46204 -59511 -45896
rect -59447 -46172 -59203 -45928
rect -59139 -46204 -58511 -45896
rect -58447 -46172 -58203 -45928
rect -58139 -46204 -57511 -45896
rect -57447 -46172 -57203 -45928
rect -57139 -46204 -56511 -45896
rect -56447 -46172 -56203 -45928
rect -56139 -46204 -55511 -45896
rect -55447 -46172 -55203 -45928
rect -55139 -46204 -54511 -45896
rect -54447 -46172 -54203 -45928
rect -54139 -46204 -53511 -45896
rect -53447 -46172 -53203 -45928
rect -53139 -46204 -52511 -45896
rect -52447 -46172 -52203 -45928
rect -52139 -46204 -51511 -45896
rect -51447 -46172 -51203 -45928
rect -51139 -46204 -50511 -45896
rect -50447 -46172 -50203 -45928
rect -50139 -46204 -49511 -45896
rect -49447 -46172 -49203 -45928
rect -49139 -46204 -48831 -45896
rect 8281 -46204 8589 -45896
rect 8653 -46172 8897 -45928
rect 8961 -46204 9589 -45896
rect 9653 -46172 9897 -45928
rect 9961 -46204 10589 -45896
rect 10653 -46172 10897 -45928
rect 10961 -46204 11589 -45896
rect 11653 -46172 11897 -45928
rect 11961 -46204 12589 -45896
rect 12653 -46172 12897 -45928
rect 12961 -46204 13589 -45896
rect 13653 -46172 13897 -45928
rect 13961 -46204 14589 -45896
rect 14653 -46172 14897 -45928
rect 14961 -46204 15589 -45896
rect 15653 -46172 15897 -45928
rect 15961 -46204 16589 -45896
rect 16653 -46172 16897 -45928
rect 16961 -46204 17589 -45896
rect 17653 -46172 17897 -45928
rect 17961 -46204 18589 -45896
rect 18653 -46172 18897 -45928
rect 18961 -46204 19589 -45896
rect 19653 -46172 19897 -45928
rect 19961 -46204 20589 -45896
rect 20653 -46172 20897 -45928
rect 20961 -46204 21589 -45896
rect 21653 -46172 21897 -45928
rect 21961 -46204 22589 -45896
rect 22653 -46172 22897 -45928
rect 22961 -46204 23589 -45896
rect 23653 -46172 23897 -45928
rect 23961 -46204 24589 -45896
rect 24653 -46172 24897 -45928
rect 24961 -46204 25589 -45896
rect 25653 -46172 25897 -45928
rect 25961 -46204 26589 -45896
rect 26653 -46172 26897 -45928
rect 26961 -46204 27589 -45896
rect 27653 -46172 27897 -45928
rect 27961 -46204 28589 -45896
rect 28653 -46172 28897 -45928
rect 28961 -46204 29589 -45896
rect 29653 -46172 29897 -45928
rect 29961 -46204 30589 -45896
rect 30653 -46172 30897 -45928
rect 30961 -46204 31589 -45896
rect 31653 -46172 31897 -45928
rect 31961 -46204 32589 -45896
rect 32653 -46172 32897 -45928
rect 32961 -46204 33589 -45896
rect 33653 -46172 33897 -45928
rect 33961 -46204 34269 -45896
rect -74479 -46544 -74171 -46236
rect -73479 -46544 -73171 -46236
rect -72479 -46544 -72171 -46236
rect -71479 -46544 -71171 -46236
rect -70479 -46544 -70171 -46236
rect -69479 -46544 -69171 -46236
rect -68479 -46544 -68171 -46236
rect -67479 -46544 -67171 -46236
rect -66479 -46544 -66171 -46236
rect -65479 -46544 -65171 -46236
rect -64479 -46544 -64171 -46236
rect -63479 -46544 -63171 -46236
rect -62479 -46544 -62171 -46236
rect -61479 -46544 -61171 -46236
rect -60479 -46544 -60171 -46236
rect -59479 -46544 -59171 -46236
rect -58479 -46544 -58171 -46236
rect -57479 -46544 -57171 -46236
rect -56479 -46544 -56171 -46236
rect -55479 -46544 -55171 -46236
rect -54479 -46544 -54171 -46236
rect -53479 -46544 -53171 -46236
rect -52479 -46544 -52171 -46236
rect -51479 -46544 -51171 -46236
rect -50479 -46544 -50171 -46236
rect -49479 -46544 -49171 -46236
rect 8621 -46544 8929 -46236
rect 9621 -46544 9929 -46236
rect 10621 -46544 10929 -46236
rect 11621 -46544 11929 -46236
rect 12621 -46544 12929 -46236
rect 13621 -46544 13929 -46236
rect 14621 -46544 14929 -46236
rect 15621 -46544 15929 -46236
rect 16621 -46544 16929 -46236
rect 17621 -46544 17929 -46236
rect 18621 -46544 18929 -46236
rect 19621 -46544 19929 -46236
rect 20621 -46544 20929 -46236
rect 21621 -46544 21929 -46236
rect 22621 -46544 22929 -46236
rect 23621 -46544 23929 -46236
rect 24621 -46544 24929 -46236
rect 25621 -46544 25929 -46236
rect 26621 -46544 26929 -46236
rect 27621 -46544 27929 -46236
rect 28621 -46544 28929 -46236
rect 29621 -46544 29929 -46236
rect 30621 -46544 30929 -46236
rect 31621 -46544 31929 -46236
rect 32621 -46544 32929 -46236
rect 33621 -46544 33929 -46236
<< metal2 >>
rect -74485 38544 -74165 38550
rect -74485 38236 -74479 38544
rect -74171 38236 -74165 38544
rect -74485 38210 -74165 38236
rect -73485 38544 -73165 38550
rect -73485 38236 -73479 38544
rect -73171 38236 -73165 38544
rect -73485 38210 -73165 38236
rect -72485 38544 -72165 38550
rect -72485 38236 -72479 38544
rect -72171 38236 -72165 38544
rect -72485 38210 -72165 38236
rect -71485 38544 -71165 38550
rect -71485 38236 -71479 38544
rect -71171 38236 -71165 38544
rect -71485 38210 -71165 38236
rect -70485 38544 -70165 38550
rect -70485 38236 -70479 38544
rect -70171 38236 -70165 38544
rect -70485 38210 -70165 38236
rect -69485 38544 -69165 38550
rect -69485 38236 -69479 38544
rect -69171 38236 -69165 38544
rect -69485 38210 -69165 38236
rect -68485 38544 -68165 38550
rect -68485 38236 -68479 38544
rect -68171 38236 -68165 38544
rect -68485 38210 -68165 38236
rect -67485 38544 -67165 38550
rect -67485 38236 -67479 38544
rect -67171 38236 -67165 38544
rect -67485 38210 -67165 38236
rect -66485 38544 -66165 38550
rect -66485 38236 -66479 38544
rect -66171 38236 -66165 38544
rect -66485 38210 -66165 38236
rect -65485 38544 -65165 38550
rect -65485 38236 -65479 38544
rect -65171 38236 -65165 38544
rect -65485 38210 -65165 38236
rect -64485 38544 -64165 38550
rect -64485 38236 -64479 38544
rect -64171 38236 -64165 38544
rect -64485 38210 -64165 38236
rect -63485 38544 -63165 38550
rect -63485 38236 -63479 38544
rect -63171 38236 -63165 38544
rect -63485 38210 -63165 38236
rect -62485 38544 -62165 38550
rect -62485 38236 -62479 38544
rect -62171 38236 -62165 38544
rect -62485 38210 -62165 38236
rect -61485 38544 -61165 38550
rect -61485 38236 -61479 38544
rect -61171 38236 -61165 38544
rect -61485 38210 -61165 38236
rect -60485 38544 -60165 38550
rect -60485 38236 -60479 38544
rect -60171 38236 -60165 38544
rect -60485 38210 -60165 38236
rect -59485 38544 -59165 38550
rect -59485 38236 -59479 38544
rect -59171 38236 -59165 38544
rect -59485 38210 -59165 38236
rect 9994 38544 10314 38550
rect 9994 38236 10000 38544
rect 10308 38236 10314 38544
rect 9994 38210 10314 38236
rect 10994 38544 11314 38550
rect 10994 38236 11000 38544
rect 11308 38236 11314 38544
rect 10994 38210 11314 38236
rect 11994 38544 12314 38550
rect 11994 38236 12000 38544
rect 12308 38236 12314 38544
rect 11994 38210 12314 38236
rect 12994 38544 13314 38550
rect 12994 38236 13000 38544
rect 13308 38236 13314 38544
rect 12994 38210 13314 38236
rect 13994 38544 14314 38550
rect 13994 38236 14000 38544
rect 14308 38236 14314 38544
rect 13994 38210 14314 38236
rect 14994 38544 15314 38550
rect 14994 38236 15000 38544
rect 15308 38236 15314 38544
rect 14994 38210 15314 38236
rect 15994 38544 16314 38550
rect 15994 38236 16000 38544
rect 16308 38236 16314 38544
rect 15994 38210 16314 38236
rect 16994 38544 17314 38550
rect 16994 38236 17000 38544
rect 17308 38236 17314 38544
rect 16994 38210 17314 38236
rect 17994 38544 18314 38550
rect 17994 38236 18000 38544
rect 18308 38236 18314 38544
rect 17994 38210 18314 38236
rect 18994 38544 19314 38550
rect 18994 38236 19000 38544
rect 19308 38236 19314 38544
rect 18994 38210 19314 38236
rect 19994 38544 20314 38550
rect 19994 38236 20000 38544
rect 20308 38236 20314 38544
rect 19994 38210 20314 38236
rect 20994 38544 21314 38550
rect 20994 38236 21000 38544
rect 21308 38236 21314 38544
rect 20994 38210 21314 38236
rect 21994 38544 22314 38550
rect 21994 38236 22000 38544
rect 22308 38236 22314 38544
rect 21994 38210 22314 38236
rect 22994 38544 23314 38550
rect 22994 38236 23000 38544
rect 23308 38236 23314 38544
rect 22994 38210 23314 38236
rect 23994 38544 24314 38550
rect 23994 38236 24000 38544
rect 24308 38236 24314 38544
rect 23994 38210 24314 38236
rect 24994 38544 25314 38550
rect 24994 38236 25000 38544
rect 25308 38236 25314 38544
rect 24994 38210 25314 38236
rect 25994 38544 26314 38550
rect 25994 38236 26000 38544
rect 26308 38236 26314 38544
rect 25994 38210 26314 38236
rect 26994 38544 27314 38550
rect 26994 38236 27000 38544
rect 27308 38236 27314 38544
rect 26994 38210 27314 38236
rect 27994 38544 28314 38550
rect 27994 38236 28000 38544
rect 28308 38236 28314 38544
rect 27994 38210 28314 38236
rect 28994 38544 29314 38550
rect 28994 38236 29000 38544
rect 29308 38236 29314 38544
rect 28994 38210 29314 38236
rect 29994 38544 30314 38550
rect 29994 38236 30000 38544
rect 30308 38236 30314 38544
rect 29994 38210 30314 38236
rect 30994 38544 31314 38550
rect 30994 38236 31000 38544
rect 31308 38236 31314 38544
rect 30994 38210 31314 38236
rect 31994 38544 32314 38550
rect 31994 38236 32000 38544
rect 32308 38236 32314 38544
rect 31994 38210 32314 38236
rect 32994 38544 33314 38550
rect 32994 38236 33000 38544
rect 33308 38236 33314 38544
rect 32994 38210 33314 38236
rect 33994 38544 34314 38550
rect 33994 38236 34000 38544
rect 34308 38236 34314 38544
rect 33994 38210 34314 38236
rect -74825 38204 -58825 38210
rect -74825 37896 -74819 38204
rect -74511 38198 -74139 38204
rect -73511 38198 -73139 38204
rect -72511 38198 -72139 38204
rect -71511 38198 -71139 38204
rect -70511 38198 -70139 38204
rect -69511 38198 -69139 38204
rect -68511 38198 -68139 38204
rect -67511 38198 -67139 38204
rect -66511 38198 -66139 38204
rect -65511 38198 -65139 38204
rect -64511 38198 -64139 38204
rect -63511 38198 -63139 38204
rect -62511 38198 -62139 38204
rect -61511 38198 -61139 38204
rect -60511 38198 -60139 38204
rect -59511 38198 -59139 38204
rect -74511 37902 -74473 38198
rect -74177 37902 -74139 38198
rect -73511 37902 -73473 38198
rect -73177 37902 -73139 38198
rect -72511 37902 -72473 38198
rect -72177 37902 -72139 38198
rect -71511 37902 -71473 38198
rect -71177 37902 -71139 38198
rect -70511 37902 -70473 38198
rect -70177 37902 -70139 38198
rect -69511 37902 -69473 38198
rect -69177 37902 -69139 38198
rect -68511 37902 -68473 38198
rect -68177 37902 -68139 38198
rect -67511 37902 -67473 38198
rect -67177 37902 -67139 38198
rect -66511 37902 -66473 38198
rect -66177 37902 -66139 38198
rect -65511 37902 -65473 38198
rect -65177 37902 -65139 38198
rect -64511 37902 -64473 38198
rect -64177 37902 -64139 38198
rect -63511 37902 -63473 38198
rect -63177 37902 -63139 38198
rect -62511 37902 -62473 38198
rect -62177 37902 -62139 38198
rect -61511 37902 -61473 38198
rect -61177 37902 -61139 38198
rect -60511 37902 -60473 38198
rect -60177 37902 -60139 38198
rect -59511 37902 -59473 38198
rect -59177 37902 -59139 38198
rect -74511 37896 -74139 37902
rect -73511 37896 -73139 37902
rect -72511 37896 -72139 37902
rect -71511 37896 -71139 37902
rect -70511 37896 -70139 37902
rect -69511 37896 -69139 37902
rect -68511 37896 -68139 37902
rect -67511 37896 -67139 37902
rect -66511 37896 -66139 37902
rect -65511 37896 -65139 37902
rect -64511 37896 -64139 37902
rect -63511 37896 -63139 37902
rect -62511 37896 -62139 37902
rect -61511 37896 -61139 37902
rect -60511 37896 -60139 37902
rect -59511 37896 -59139 37902
rect -58831 37896 -58825 38204
rect -74825 37890 -58825 37896
rect 9654 38204 34654 38210
rect 9654 37896 9660 38204
rect 9968 38198 10340 38204
rect 10968 38198 11340 38204
rect 11968 38198 12340 38204
rect 12968 38198 13340 38204
rect 13968 38198 14340 38204
rect 14968 38198 15340 38204
rect 15968 38198 16340 38204
rect 16968 38198 17340 38204
rect 17968 38198 18340 38204
rect 18968 38198 19340 38204
rect 19968 38198 20340 38204
rect 20968 38198 21340 38204
rect 21968 38198 22340 38204
rect 22968 38198 23340 38204
rect 23968 38198 24340 38204
rect 24968 38198 25340 38204
rect 25968 38198 26340 38204
rect 26968 38198 27340 38204
rect 27968 38198 28340 38204
rect 28968 38198 29340 38204
rect 29968 38198 30340 38204
rect 30968 38198 31340 38204
rect 31968 38198 32340 38204
rect 32968 38198 33340 38204
rect 33968 38198 34340 38204
rect 9968 37902 10006 38198
rect 10302 37902 10340 38198
rect 10968 37902 11006 38198
rect 11302 37902 11340 38198
rect 11968 37902 12006 38198
rect 12302 37902 12340 38198
rect 12968 37902 13006 38198
rect 13302 37902 13340 38198
rect 13968 37902 14006 38198
rect 14302 37902 14340 38198
rect 14968 37902 15006 38198
rect 15302 37902 15340 38198
rect 15968 37902 16006 38198
rect 16302 37902 16340 38198
rect 16968 37902 17006 38198
rect 17302 37902 17340 38198
rect 17968 37902 18006 38198
rect 18302 37902 18340 38198
rect 18968 37902 19006 38198
rect 19302 37902 19340 38198
rect 19968 37902 20006 38198
rect 20302 37902 20340 38198
rect 20968 37902 21006 38198
rect 21302 37902 21340 38198
rect 21968 37902 22006 38198
rect 22302 37902 22340 38198
rect 22968 37902 23006 38198
rect 23302 37902 23340 38198
rect 23968 37902 24006 38198
rect 24302 37902 24340 38198
rect 24968 37902 25006 38198
rect 25302 37902 25340 38198
rect 25968 37902 26006 38198
rect 26302 37902 26340 38198
rect 26968 37902 27006 38198
rect 27302 37902 27340 38198
rect 27968 37902 28006 38198
rect 28302 37902 28340 38198
rect 28968 37902 29006 38198
rect 29302 37902 29340 38198
rect 29968 37902 30006 38198
rect 30302 37902 30340 38198
rect 30968 37902 31006 38198
rect 31302 37902 31340 38198
rect 31968 37902 32006 38198
rect 32302 37902 32340 38198
rect 32968 37902 33006 38198
rect 33302 37902 33340 38198
rect 33968 37902 34006 38198
rect 34302 37902 34340 38198
rect 9968 37896 10340 37902
rect 10968 37896 11340 37902
rect 11968 37896 12340 37902
rect 12968 37896 13340 37902
rect 13968 37896 14340 37902
rect 14968 37896 15340 37902
rect 15968 37896 16340 37902
rect 16968 37896 17340 37902
rect 17968 37896 18340 37902
rect 18968 37896 19340 37902
rect 19968 37896 20340 37902
rect 20968 37896 21340 37902
rect 21968 37896 22340 37902
rect 22968 37896 23340 37902
rect 23968 37896 24340 37902
rect 24968 37896 25340 37902
rect 25968 37896 26340 37902
rect 26968 37896 27340 37902
rect 27968 37896 28340 37902
rect 28968 37896 29340 37902
rect 29968 37896 30340 37902
rect 30968 37896 31340 37902
rect 31968 37896 32340 37902
rect 32968 37896 33340 37902
rect 33968 37896 34340 37902
rect 34648 37896 34654 38204
rect 9654 37890 34654 37896
rect -74485 37864 -74165 37890
rect -74485 37236 -74479 37864
rect -74171 37236 -74165 37864
rect -74485 37210 -74165 37236
rect -73485 37864 -73165 37890
rect -73485 37236 -73479 37864
rect -73171 37236 -73165 37864
rect -73485 37210 -73165 37236
rect -72485 37864 -72165 37890
rect -72485 37236 -72479 37864
rect -72171 37236 -72165 37864
rect -72485 37210 -72165 37236
rect -71485 37864 -71165 37890
rect -71485 37236 -71479 37864
rect -71171 37236 -71165 37864
rect -71485 37210 -71165 37236
rect -70485 37864 -70165 37890
rect -70485 37236 -70479 37864
rect -70171 37236 -70165 37864
rect -70485 37210 -70165 37236
rect -69485 37864 -69165 37890
rect -69485 37236 -69479 37864
rect -69171 37236 -69165 37864
rect -69485 37210 -69165 37236
rect -68485 37864 -68165 37890
rect -68485 37236 -68479 37864
rect -68171 37236 -68165 37864
rect -68485 37210 -68165 37236
rect -67485 37864 -67165 37890
rect -67485 37236 -67479 37864
rect -67171 37236 -67165 37864
rect -67485 37210 -67165 37236
rect -66485 37864 -66165 37890
rect -66485 37236 -66479 37864
rect -66171 37236 -66165 37864
rect -66485 37210 -66165 37236
rect -65485 37864 -65165 37890
rect -65485 37236 -65479 37864
rect -65171 37236 -65165 37864
rect -65485 37210 -65165 37236
rect -64485 37864 -64165 37890
rect -64485 37236 -64479 37864
rect -64171 37236 -64165 37864
rect -64485 37210 -64165 37236
rect -63485 37864 -63165 37890
rect -63485 37236 -63479 37864
rect -63171 37236 -63165 37864
rect -63485 37210 -63165 37236
rect -62485 37864 -62165 37890
rect -62485 37236 -62479 37864
rect -62171 37236 -62165 37864
rect -62485 37210 -62165 37236
rect -61485 37864 -61165 37890
rect -61485 37236 -61479 37864
rect -61171 37236 -61165 37864
rect -61485 37210 -61165 37236
rect -60485 37864 -60165 37890
rect -60485 37236 -60479 37864
rect -60171 37236 -60165 37864
rect -60485 37210 -60165 37236
rect -59485 37864 -59165 37890
rect -59485 37236 -59479 37864
rect -59171 37236 -59165 37864
rect -59485 37210 -59165 37236
rect 9994 37864 10314 37890
rect 9994 37236 10000 37864
rect 10308 37236 10314 37864
rect 9994 37210 10314 37236
rect 10994 37864 11314 37890
rect 10994 37236 11000 37864
rect 11308 37236 11314 37864
rect 10994 37210 11314 37236
rect 11994 37864 12314 37890
rect 11994 37236 12000 37864
rect 12308 37236 12314 37864
rect 11994 37210 12314 37236
rect 12994 37864 13314 37890
rect 12994 37236 13000 37864
rect 13308 37236 13314 37864
rect 12994 37210 13314 37236
rect 13994 37864 14314 37890
rect 13994 37236 14000 37864
rect 14308 37236 14314 37864
rect 13994 37210 14314 37236
rect 14994 37864 15314 37890
rect 14994 37236 15000 37864
rect 15308 37236 15314 37864
rect 14994 37210 15314 37236
rect 15994 37864 16314 37890
rect 15994 37236 16000 37864
rect 16308 37236 16314 37864
rect 15994 37210 16314 37236
rect 16994 37864 17314 37890
rect 16994 37236 17000 37864
rect 17308 37236 17314 37864
rect 16994 37210 17314 37236
rect 17994 37864 18314 37890
rect 17994 37236 18000 37864
rect 18308 37236 18314 37864
rect 17994 37210 18314 37236
rect 18994 37864 19314 37890
rect 18994 37236 19000 37864
rect 19308 37236 19314 37864
rect 18994 37210 19314 37236
rect 19994 37864 20314 37890
rect 19994 37236 20000 37864
rect 20308 37236 20314 37864
rect 19994 37210 20314 37236
rect 20994 37864 21314 37890
rect 20994 37236 21000 37864
rect 21308 37236 21314 37864
rect 20994 37210 21314 37236
rect 21994 37864 22314 37890
rect 21994 37236 22000 37864
rect 22308 37236 22314 37864
rect 21994 37210 22314 37236
rect 22994 37864 23314 37890
rect 22994 37236 23000 37864
rect 23308 37236 23314 37864
rect 22994 37210 23314 37236
rect 23994 37864 24314 37890
rect 23994 37236 24000 37864
rect 24308 37236 24314 37864
rect 23994 37210 24314 37236
rect 24994 37864 25314 37890
rect 24994 37236 25000 37864
rect 25308 37236 25314 37864
rect 24994 37210 25314 37236
rect 25994 37864 26314 37890
rect 25994 37236 26000 37864
rect 26308 37236 26314 37864
rect 25994 37210 26314 37236
rect 26994 37864 27314 37890
rect 26994 37236 27000 37864
rect 27308 37236 27314 37864
rect 26994 37210 27314 37236
rect 27994 37864 28314 37890
rect 27994 37236 28000 37864
rect 28308 37236 28314 37864
rect 27994 37210 28314 37236
rect 28994 37864 29314 37890
rect 28994 37236 29000 37864
rect 29308 37236 29314 37864
rect 28994 37210 29314 37236
rect 29994 37864 30314 37890
rect 29994 37236 30000 37864
rect 30308 37236 30314 37864
rect 29994 37210 30314 37236
rect 30994 37864 31314 37890
rect 30994 37236 31000 37864
rect 31308 37236 31314 37864
rect 30994 37210 31314 37236
rect 31994 37864 32314 37890
rect 31994 37236 32000 37864
rect 32308 37236 32314 37864
rect 31994 37210 32314 37236
rect 32994 37864 33314 37890
rect 32994 37236 33000 37864
rect 33308 37236 33314 37864
rect 32994 37210 33314 37236
rect 33994 37864 34314 37890
rect 33994 37236 34000 37864
rect 34308 37236 34314 37864
rect 33994 37210 34314 37236
rect -74825 37204 -58825 37210
rect -74825 36896 -74819 37204
rect -74511 37198 -74139 37204
rect -73511 37198 -73139 37204
rect -72511 37198 -72139 37204
rect -71511 37198 -71139 37204
rect -70511 37198 -70139 37204
rect -69511 37198 -69139 37204
rect -68511 37198 -68139 37204
rect -67511 37198 -67139 37204
rect -66511 37198 -66139 37204
rect -65511 37198 -65139 37204
rect -64511 37198 -64139 37204
rect -63511 37198 -63139 37204
rect -62511 37198 -62139 37204
rect -61511 37198 -61139 37204
rect -60511 37198 -60139 37204
rect -59511 37198 -59139 37204
rect -74511 36902 -74473 37198
rect -74177 36902 -74139 37198
rect -73511 36902 -73473 37198
rect -73177 36902 -73139 37198
rect -72511 36902 -72473 37198
rect -72177 36902 -72139 37198
rect -71511 36902 -71473 37198
rect -71177 36902 -71139 37198
rect -70511 36902 -70473 37198
rect -70177 36902 -70139 37198
rect -69511 36902 -69473 37198
rect -69177 36902 -69139 37198
rect -68511 36902 -68473 37198
rect -68177 36902 -68139 37198
rect -67511 36902 -67473 37198
rect -67177 36902 -67139 37198
rect -66511 36902 -66473 37198
rect -66177 36902 -66139 37198
rect -65511 36902 -65473 37198
rect -65177 36902 -65139 37198
rect -64511 36902 -64473 37198
rect -64177 36902 -64139 37198
rect -63511 36902 -63473 37198
rect -63177 36902 -63139 37198
rect -62511 36902 -62473 37198
rect -62177 36902 -62139 37198
rect -61511 36902 -61473 37198
rect -61177 36902 -61139 37198
rect -60511 36902 -60473 37198
rect -60177 36902 -60139 37198
rect -59511 36902 -59473 37198
rect -59177 36902 -59139 37198
rect -74511 36896 -74139 36902
rect -73511 36896 -73139 36902
rect -72511 36896 -72139 36902
rect -71511 36896 -71139 36902
rect -70511 36896 -70139 36902
rect -69511 36896 -69139 36902
rect -68511 36896 -68139 36902
rect -67511 36896 -67139 36902
rect -66511 36896 -66139 36902
rect -65511 36896 -65139 36902
rect -64511 36896 -64139 36902
rect -63511 36896 -63139 36902
rect -62511 36896 -62139 36902
rect -61511 36896 -61139 36902
rect -60511 36896 -60139 36902
rect -59511 36896 -59139 36902
rect -58831 36896 -58825 37204
rect -74825 36890 -58825 36896
rect 9654 37204 34654 37210
rect 9654 36896 9660 37204
rect 9968 37198 10340 37204
rect 10968 37198 11340 37204
rect 11968 37198 12340 37204
rect 12968 37198 13340 37204
rect 13968 37198 14340 37204
rect 14968 37198 15340 37204
rect 15968 37198 16340 37204
rect 16968 37198 17340 37204
rect 17968 37198 18340 37204
rect 18968 37198 19340 37204
rect 19968 37198 20340 37204
rect 20968 37198 21340 37204
rect 21968 37198 22340 37204
rect 22968 37198 23340 37204
rect 23968 37198 24340 37204
rect 24968 37198 25340 37204
rect 25968 37198 26340 37204
rect 26968 37198 27340 37204
rect 27968 37198 28340 37204
rect 28968 37198 29340 37204
rect 29968 37198 30340 37204
rect 30968 37198 31340 37204
rect 31968 37198 32340 37204
rect 32968 37198 33340 37204
rect 33968 37198 34340 37204
rect 9968 36902 10006 37198
rect 10302 36902 10340 37198
rect 10968 36902 11006 37198
rect 11302 36902 11340 37198
rect 11968 36902 12006 37198
rect 12302 36902 12340 37198
rect 12968 36902 13006 37198
rect 13302 36902 13340 37198
rect 13968 36902 14006 37198
rect 14302 36902 14340 37198
rect 14968 36902 15006 37198
rect 15302 36902 15340 37198
rect 15968 36902 16006 37198
rect 16302 36902 16340 37198
rect 16968 36902 17006 37198
rect 17302 36902 17340 37198
rect 17968 36902 18006 37198
rect 18302 36902 18340 37198
rect 18968 36902 19006 37198
rect 19302 36902 19340 37198
rect 19968 36902 20006 37198
rect 20302 36902 20340 37198
rect 20968 36902 21006 37198
rect 21302 36902 21340 37198
rect 21968 36902 22006 37198
rect 22302 36902 22340 37198
rect 22968 36902 23006 37198
rect 23302 36902 23340 37198
rect 23968 36902 24006 37198
rect 24302 36902 24340 37198
rect 24968 36902 25006 37198
rect 25302 36902 25340 37198
rect 25968 36902 26006 37198
rect 26302 36902 26340 37198
rect 26968 36902 27006 37198
rect 27302 36902 27340 37198
rect 27968 36902 28006 37198
rect 28302 36902 28340 37198
rect 28968 36902 29006 37198
rect 29302 36902 29340 37198
rect 29968 36902 30006 37198
rect 30302 36902 30340 37198
rect 30968 36902 31006 37198
rect 31302 36902 31340 37198
rect 31968 36902 32006 37198
rect 32302 36902 32340 37198
rect 32968 36902 33006 37198
rect 33302 36902 33340 37198
rect 33968 36902 34006 37198
rect 34302 36902 34340 37198
rect 9968 36896 10340 36902
rect 10968 36896 11340 36902
rect 11968 36896 12340 36902
rect 12968 36896 13340 36902
rect 13968 36896 14340 36902
rect 14968 36896 15340 36902
rect 15968 36896 16340 36902
rect 16968 36896 17340 36902
rect 17968 36896 18340 36902
rect 18968 36896 19340 36902
rect 19968 36896 20340 36902
rect 20968 36896 21340 36902
rect 21968 36896 22340 36902
rect 22968 36896 23340 36902
rect 23968 36896 24340 36902
rect 24968 36896 25340 36902
rect 25968 36896 26340 36902
rect 26968 36896 27340 36902
rect 27968 36896 28340 36902
rect 28968 36896 29340 36902
rect 29968 36896 30340 36902
rect 30968 36896 31340 36902
rect 31968 36896 32340 36902
rect 32968 36896 33340 36902
rect 33968 36896 34340 36902
rect 34648 36896 34654 37204
rect 9654 36890 34654 36896
rect -74485 36864 -74165 36890
rect -74485 36236 -74479 36864
rect -74171 36236 -74165 36864
rect -74485 36210 -74165 36236
rect -73485 36864 -73165 36890
rect -73485 36236 -73479 36864
rect -73171 36236 -73165 36864
rect -73485 36210 -73165 36236
rect -72485 36864 -72165 36890
rect -72485 36236 -72479 36864
rect -72171 36236 -72165 36864
rect -72485 36210 -72165 36236
rect -71485 36864 -71165 36890
rect -71485 36236 -71479 36864
rect -71171 36236 -71165 36864
rect -71485 36210 -71165 36236
rect -70485 36864 -70165 36890
rect -70485 36236 -70479 36864
rect -70171 36236 -70165 36864
rect -70485 36210 -70165 36236
rect -69485 36864 -69165 36890
rect -69485 36236 -69479 36864
rect -69171 36236 -69165 36864
rect -69485 36210 -69165 36236
rect -68485 36864 -68165 36890
rect -68485 36236 -68479 36864
rect -68171 36236 -68165 36864
rect -68485 36210 -68165 36236
rect -67485 36864 -67165 36890
rect -67485 36236 -67479 36864
rect -67171 36236 -67165 36864
rect -67485 36210 -67165 36236
rect -66485 36864 -66165 36890
rect -66485 36236 -66479 36864
rect -66171 36236 -66165 36864
rect -66485 36210 -66165 36236
rect -65485 36864 -65165 36890
rect -65485 36236 -65479 36864
rect -65171 36236 -65165 36864
rect -65485 36210 -65165 36236
rect -64485 36864 -64165 36890
rect -64485 36236 -64479 36864
rect -64171 36236 -64165 36864
rect -64485 36210 -64165 36236
rect -63485 36864 -63165 36890
rect -63485 36236 -63479 36864
rect -63171 36236 -63165 36864
rect -63485 36210 -63165 36236
rect -62485 36864 -62165 36890
rect -62485 36236 -62479 36864
rect -62171 36236 -62165 36864
rect -62485 36210 -62165 36236
rect -61485 36864 -61165 36890
rect -61485 36236 -61479 36864
rect -61171 36236 -61165 36864
rect -61485 36210 -61165 36236
rect -60485 36864 -60165 36890
rect -60485 36236 -60479 36864
rect -60171 36236 -60165 36864
rect -60485 36210 -60165 36236
rect -59485 36864 -59165 36890
rect -59485 36236 -59479 36864
rect -59171 36236 -59165 36864
rect -59485 36210 -59165 36236
rect 9994 36864 10314 36890
rect 9994 36236 10000 36864
rect 10308 36236 10314 36864
rect 9994 36210 10314 36236
rect 10994 36864 11314 36890
rect 10994 36236 11000 36864
rect 11308 36236 11314 36864
rect 10994 36210 11314 36236
rect 11994 36864 12314 36890
rect 11994 36236 12000 36864
rect 12308 36236 12314 36864
rect 11994 36210 12314 36236
rect 12994 36864 13314 36890
rect 12994 36236 13000 36864
rect 13308 36236 13314 36864
rect 12994 36210 13314 36236
rect 13994 36864 14314 36890
rect 13994 36236 14000 36864
rect 14308 36236 14314 36864
rect 13994 36210 14314 36236
rect 14994 36864 15314 36890
rect 14994 36236 15000 36864
rect 15308 36236 15314 36864
rect 14994 36210 15314 36236
rect 15994 36864 16314 36890
rect 15994 36236 16000 36864
rect 16308 36236 16314 36864
rect 15994 36210 16314 36236
rect 16994 36864 17314 36890
rect 16994 36236 17000 36864
rect 17308 36236 17314 36864
rect 16994 36210 17314 36236
rect 17994 36864 18314 36890
rect 17994 36236 18000 36864
rect 18308 36236 18314 36864
rect 17994 36210 18314 36236
rect 18994 36864 19314 36890
rect 18994 36236 19000 36864
rect 19308 36236 19314 36864
rect 18994 36210 19314 36236
rect 19994 36864 20314 36890
rect 19994 36236 20000 36864
rect 20308 36236 20314 36864
rect 19994 36210 20314 36236
rect 20994 36864 21314 36890
rect 20994 36236 21000 36864
rect 21308 36236 21314 36864
rect 20994 36210 21314 36236
rect 21994 36864 22314 36890
rect 21994 36236 22000 36864
rect 22308 36236 22314 36864
rect 21994 36210 22314 36236
rect 22994 36864 23314 36890
rect 22994 36236 23000 36864
rect 23308 36236 23314 36864
rect 22994 36210 23314 36236
rect 23994 36864 24314 36890
rect 23994 36236 24000 36864
rect 24308 36236 24314 36864
rect 23994 36210 24314 36236
rect 24994 36864 25314 36890
rect 24994 36236 25000 36864
rect 25308 36236 25314 36864
rect 24994 36210 25314 36236
rect 25994 36864 26314 36890
rect 25994 36236 26000 36864
rect 26308 36236 26314 36864
rect 25994 36210 26314 36236
rect 26994 36864 27314 36890
rect 26994 36236 27000 36864
rect 27308 36236 27314 36864
rect 26994 36210 27314 36236
rect 27994 36864 28314 36890
rect 27994 36236 28000 36864
rect 28308 36236 28314 36864
rect 27994 36210 28314 36236
rect 28994 36864 29314 36890
rect 28994 36236 29000 36864
rect 29308 36236 29314 36864
rect 28994 36210 29314 36236
rect 29994 36864 30314 36890
rect 29994 36236 30000 36864
rect 30308 36236 30314 36864
rect 29994 36210 30314 36236
rect 30994 36864 31314 36890
rect 30994 36236 31000 36864
rect 31308 36236 31314 36864
rect 30994 36210 31314 36236
rect 31994 36864 32314 36890
rect 31994 36236 32000 36864
rect 32308 36236 32314 36864
rect 31994 36210 32314 36236
rect 32994 36864 33314 36890
rect 32994 36236 33000 36864
rect 33308 36236 33314 36864
rect 32994 36210 33314 36236
rect 33994 36864 34314 36890
rect 33994 36236 34000 36864
rect 34308 36236 34314 36864
rect 33994 36210 34314 36236
rect -74825 36204 -58825 36210
rect -74825 35896 -74819 36204
rect -74511 36198 -74139 36204
rect -73511 36198 -73139 36204
rect -72511 36198 -72139 36204
rect -71511 36198 -71139 36204
rect -70511 36198 -70139 36204
rect -69511 36198 -69139 36204
rect -68511 36198 -68139 36204
rect -67511 36198 -67139 36204
rect -66511 36198 -66139 36204
rect -65511 36198 -65139 36204
rect -64511 36198 -64139 36204
rect -63511 36198 -63139 36204
rect -62511 36198 -62139 36204
rect -61511 36198 -61139 36204
rect -60511 36198 -60139 36204
rect -59511 36198 -59139 36204
rect -74511 35902 -74473 36198
rect -74177 35902 -74139 36198
rect -73511 35902 -73473 36198
rect -73177 35902 -73139 36198
rect -72511 35902 -72473 36198
rect -72177 35902 -72139 36198
rect -71511 35902 -71473 36198
rect -71177 35902 -71139 36198
rect -70511 35902 -70473 36198
rect -70177 35902 -70139 36198
rect -69511 35902 -69473 36198
rect -69177 35902 -69139 36198
rect -68511 35902 -68473 36198
rect -68177 35902 -68139 36198
rect -67511 35902 -67473 36198
rect -67177 35902 -67139 36198
rect -66511 35902 -66473 36198
rect -66177 35902 -66139 36198
rect -65511 35902 -65473 36198
rect -65177 35902 -65139 36198
rect -64511 35902 -64473 36198
rect -64177 35902 -64139 36198
rect -63511 35902 -63473 36198
rect -63177 35902 -63139 36198
rect -62511 35902 -62473 36198
rect -62177 35902 -62139 36198
rect -61511 35902 -61473 36198
rect -61177 35902 -61139 36198
rect -60511 35902 -60473 36198
rect -60177 35902 -60139 36198
rect -59511 35902 -59473 36198
rect -59177 35902 -59139 36198
rect -74511 35896 -74139 35902
rect -73511 35896 -73139 35902
rect -72511 35896 -72139 35902
rect -71511 35896 -71139 35902
rect -70511 35896 -70139 35902
rect -69511 35896 -69139 35902
rect -68511 35896 -68139 35902
rect -67511 35896 -67139 35902
rect -66511 35896 -66139 35902
rect -65511 35896 -65139 35902
rect -64511 35896 -64139 35902
rect -63511 35896 -63139 35902
rect -62511 35896 -62139 35902
rect -61511 35896 -61139 35902
rect -60511 35896 -60139 35902
rect -59511 35896 -59139 35902
rect -58831 35896 -58825 36204
rect -74825 35890 -58825 35896
rect 9654 36204 34654 36210
rect 9654 35896 9660 36204
rect 9968 36198 10340 36204
rect 10968 36198 11340 36204
rect 11968 36198 12340 36204
rect 12968 36198 13340 36204
rect 13968 36198 14340 36204
rect 14968 36198 15340 36204
rect 15968 36198 16340 36204
rect 16968 36198 17340 36204
rect 17968 36198 18340 36204
rect 18968 36198 19340 36204
rect 19968 36198 20340 36204
rect 20968 36198 21340 36204
rect 21968 36198 22340 36204
rect 22968 36198 23340 36204
rect 23968 36198 24340 36204
rect 24968 36198 25340 36204
rect 25968 36198 26340 36204
rect 26968 36198 27340 36204
rect 27968 36198 28340 36204
rect 28968 36198 29340 36204
rect 29968 36198 30340 36204
rect 30968 36198 31340 36204
rect 31968 36198 32340 36204
rect 32968 36198 33340 36204
rect 33968 36198 34340 36204
rect 9968 35902 10006 36198
rect 10302 35902 10340 36198
rect 10968 35902 11006 36198
rect 11302 35902 11340 36198
rect 11968 35902 12006 36198
rect 12302 35902 12340 36198
rect 12968 35902 13006 36198
rect 13302 35902 13340 36198
rect 13968 35902 14006 36198
rect 14302 35902 14340 36198
rect 14968 35902 15006 36198
rect 15302 35902 15340 36198
rect 15968 35902 16006 36198
rect 16302 35902 16340 36198
rect 16968 35902 17006 36198
rect 17302 35902 17340 36198
rect 17968 35902 18006 36198
rect 18302 35902 18340 36198
rect 18968 35902 19006 36198
rect 19302 35902 19340 36198
rect 19968 35902 20006 36198
rect 20302 35902 20340 36198
rect 20968 35902 21006 36198
rect 21302 35902 21340 36198
rect 21968 35902 22006 36198
rect 22302 35902 22340 36198
rect 22968 35902 23006 36198
rect 23302 35902 23340 36198
rect 23968 35902 24006 36198
rect 24302 35902 24340 36198
rect 24968 35902 25006 36198
rect 25302 35902 25340 36198
rect 25968 35902 26006 36198
rect 26302 35902 26340 36198
rect 26968 35902 27006 36198
rect 27302 35902 27340 36198
rect 27968 35902 28006 36198
rect 28302 35902 28340 36198
rect 28968 35902 29006 36198
rect 29302 35902 29340 36198
rect 29968 35902 30006 36198
rect 30302 35902 30340 36198
rect 30968 35902 31006 36198
rect 31302 35902 31340 36198
rect 31968 35902 32006 36198
rect 32302 35902 32340 36198
rect 32968 35902 33006 36198
rect 33302 35902 33340 36198
rect 33968 35902 34006 36198
rect 34302 35902 34340 36198
rect 9968 35896 10340 35902
rect 10968 35896 11340 35902
rect 11968 35896 12340 35902
rect 12968 35896 13340 35902
rect 13968 35896 14340 35902
rect 14968 35896 15340 35902
rect 15968 35896 16340 35902
rect 16968 35896 17340 35902
rect 17968 35896 18340 35902
rect 18968 35896 19340 35902
rect 19968 35896 20340 35902
rect 20968 35896 21340 35902
rect 21968 35896 22340 35902
rect 22968 35896 23340 35902
rect 23968 35896 24340 35902
rect 24968 35896 25340 35902
rect 25968 35896 26340 35902
rect 26968 35896 27340 35902
rect 27968 35896 28340 35902
rect 28968 35896 29340 35902
rect 29968 35896 30340 35902
rect 30968 35896 31340 35902
rect 31968 35896 32340 35902
rect 32968 35896 33340 35902
rect 33968 35896 34340 35902
rect 34648 35896 34654 36204
rect 9654 35890 34654 35896
rect -74485 35864 -74165 35890
rect -74485 35236 -74479 35864
rect -74171 35236 -74165 35864
rect -74485 35210 -74165 35236
rect -73485 35864 -73165 35890
rect -73485 35236 -73479 35864
rect -73171 35236 -73165 35864
rect -73485 35210 -73165 35236
rect -72485 35864 -72165 35890
rect -72485 35236 -72479 35864
rect -72171 35236 -72165 35864
rect -72485 35210 -72165 35236
rect -71485 35864 -71165 35890
rect -71485 35236 -71479 35864
rect -71171 35236 -71165 35864
rect -71485 35210 -71165 35236
rect -70485 35864 -70165 35890
rect -70485 35236 -70479 35864
rect -70171 35236 -70165 35864
rect -70485 35210 -70165 35236
rect -69485 35864 -69165 35890
rect -69485 35236 -69479 35864
rect -69171 35236 -69165 35864
rect -69485 35210 -69165 35236
rect -68485 35864 -68165 35890
rect -68485 35236 -68479 35864
rect -68171 35236 -68165 35864
rect -68485 35210 -68165 35236
rect -67485 35864 -67165 35890
rect -67485 35236 -67479 35864
rect -67171 35236 -67165 35864
rect -67485 35210 -67165 35236
rect -66485 35864 -66165 35890
rect -66485 35236 -66479 35864
rect -66171 35236 -66165 35864
rect -66485 35210 -66165 35236
rect -65485 35864 -65165 35890
rect -65485 35236 -65479 35864
rect -65171 35236 -65165 35864
rect -65485 35210 -65165 35236
rect -64485 35864 -64165 35890
rect -64485 35236 -64479 35864
rect -64171 35236 -64165 35864
rect -64485 35210 -64165 35236
rect -63485 35864 -63165 35890
rect -63485 35236 -63479 35864
rect -63171 35236 -63165 35864
rect -63485 35210 -63165 35236
rect -62485 35864 -62165 35890
rect -62485 35236 -62479 35864
rect -62171 35236 -62165 35864
rect -62485 35210 -62165 35236
rect -61485 35864 -61165 35890
rect -61485 35236 -61479 35864
rect -61171 35236 -61165 35864
rect -61485 35210 -61165 35236
rect -60485 35864 -60165 35890
rect -60485 35236 -60479 35864
rect -60171 35236 -60165 35864
rect -60485 35210 -60165 35236
rect -59485 35864 -59165 35890
rect -59485 35236 -59479 35864
rect -59171 35236 -59165 35864
rect -59485 35210 -59165 35236
rect 9994 35864 10314 35890
rect 9994 35236 10000 35864
rect 10308 35236 10314 35864
rect 9994 35210 10314 35236
rect 10994 35864 11314 35890
rect 10994 35236 11000 35864
rect 11308 35236 11314 35864
rect 10994 35210 11314 35236
rect 11994 35864 12314 35890
rect 11994 35236 12000 35864
rect 12308 35236 12314 35864
rect 11994 35210 12314 35236
rect 12994 35864 13314 35890
rect 12994 35236 13000 35864
rect 13308 35236 13314 35864
rect 12994 35210 13314 35236
rect 13994 35864 14314 35890
rect 13994 35236 14000 35864
rect 14308 35236 14314 35864
rect 13994 35210 14314 35236
rect 14994 35864 15314 35890
rect 14994 35236 15000 35864
rect 15308 35236 15314 35864
rect 14994 35210 15314 35236
rect 15994 35864 16314 35890
rect 15994 35236 16000 35864
rect 16308 35236 16314 35864
rect 15994 35210 16314 35236
rect 16994 35864 17314 35890
rect 16994 35236 17000 35864
rect 17308 35236 17314 35864
rect 16994 35210 17314 35236
rect 17994 35864 18314 35890
rect 17994 35236 18000 35864
rect 18308 35236 18314 35864
rect 17994 35210 18314 35236
rect 18994 35864 19314 35890
rect 18994 35236 19000 35864
rect 19308 35236 19314 35864
rect 18994 35210 19314 35236
rect 19994 35864 20314 35890
rect 19994 35236 20000 35864
rect 20308 35236 20314 35864
rect 19994 35210 20314 35236
rect 20994 35864 21314 35890
rect 20994 35236 21000 35864
rect 21308 35236 21314 35864
rect 20994 35210 21314 35236
rect 21994 35864 22314 35890
rect 21994 35236 22000 35864
rect 22308 35236 22314 35864
rect 21994 35210 22314 35236
rect 22994 35864 23314 35890
rect 22994 35236 23000 35864
rect 23308 35236 23314 35864
rect 22994 35210 23314 35236
rect 23994 35864 24314 35890
rect 23994 35236 24000 35864
rect 24308 35236 24314 35864
rect 23994 35210 24314 35236
rect 24994 35864 25314 35890
rect 24994 35236 25000 35864
rect 25308 35236 25314 35864
rect 24994 35210 25314 35236
rect 25994 35864 26314 35890
rect 25994 35236 26000 35864
rect 26308 35236 26314 35864
rect 25994 35210 26314 35236
rect 26994 35864 27314 35890
rect 26994 35236 27000 35864
rect 27308 35236 27314 35864
rect 26994 35210 27314 35236
rect 27994 35864 28314 35890
rect 27994 35236 28000 35864
rect 28308 35236 28314 35864
rect 27994 35210 28314 35236
rect 28994 35864 29314 35890
rect 28994 35236 29000 35864
rect 29308 35236 29314 35864
rect 28994 35210 29314 35236
rect 29994 35864 30314 35890
rect 29994 35236 30000 35864
rect 30308 35236 30314 35864
rect 29994 35210 30314 35236
rect 30994 35864 31314 35890
rect 30994 35236 31000 35864
rect 31308 35236 31314 35864
rect 30994 35210 31314 35236
rect 31994 35864 32314 35890
rect 31994 35236 32000 35864
rect 32308 35236 32314 35864
rect 31994 35210 32314 35236
rect 32994 35864 33314 35890
rect 32994 35236 33000 35864
rect 33308 35236 33314 35864
rect 32994 35210 33314 35236
rect 33994 35864 34314 35890
rect 33994 35236 34000 35864
rect 34308 35236 34314 35864
rect 33994 35210 34314 35236
rect -74825 35204 -58825 35210
rect -74825 34896 -74819 35204
rect -74511 35198 -74139 35204
rect -73511 35198 -73139 35204
rect -72511 35198 -72139 35204
rect -71511 35198 -71139 35204
rect -70511 35198 -70139 35204
rect -69511 35198 -69139 35204
rect -68511 35198 -68139 35204
rect -67511 35198 -67139 35204
rect -66511 35198 -66139 35204
rect -65511 35198 -65139 35204
rect -64511 35198 -64139 35204
rect -63511 35198 -63139 35204
rect -62511 35198 -62139 35204
rect -61511 35198 -61139 35204
rect -60511 35198 -60139 35204
rect -59511 35198 -59139 35204
rect -74511 34902 -74473 35198
rect -74177 34902 -74139 35198
rect -73511 34902 -73473 35198
rect -73177 34902 -73139 35198
rect -72511 34902 -72473 35198
rect -72177 34902 -72139 35198
rect -71511 34902 -71473 35198
rect -71177 34902 -71139 35198
rect -70511 34902 -70473 35198
rect -70177 34902 -70139 35198
rect -69511 34902 -69473 35198
rect -69177 34902 -69139 35198
rect -68511 34902 -68473 35198
rect -68177 34902 -68139 35198
rect -67511 34902 -67473 35198
rect -67177 34902 -67139 35198
rect -66511 34902 -66473 35198
rect -66177 34902 -66139 35198
rect -65511 34902 -65473 35198
rect -65177 34902 -65139 35198
rect -64511 34902 -64473 35198
rect -64177 34902 -64139 35198
rect -63511 34902 -63473 35198
rect -63177 34902 -63139 35198
rect -62511 34902 -62473 35198
rect -62177 34902 -62139 35198
rect -61511 34902 -61473 35198
rect -61177 34902 -61139 35198
rect -60511 34902 -60473 35198
rect -60177 34902 -60139 35198
rect -59511 34902 -59473 35198
rect -59177 34902 -59139 35198
rect -74511 34896 -74139 34902
rect -73511 34896 -73139 34902
rect -72511 34896 -72139 34902
rect -71511 34896 -71139 34902
rect -70511 34896 -70139 34902
rect -69511 34896 -69139 34902
rect -68511 34896 -68139 34902
rect -67511 34896 -67139 34902
rect -66511 34896 -66139 34902
rect -65511 34896 -65139 34902
rect -64511 34896 -64139 34902
rect -63511 34896 -63139 34902
rect -62511 34896 -62139 34902
rect -61511 34896 -61139 34902
rect -60511 34896 -60139 34902
rect -59511 34896 -59139 34902
rect -58831 34896 -58825 35204
rect -74825 34890 -58825 34896
rect 9654 35204 34654 35210
rect 9654 34896 9660 35204
rect 9968 35198 10340 35204
rect 10968 35198 11340 35204
rect 11968 35198 12340 35204
rect 12968 35198 13340 35204
rect 13968 35198 14340 35204
rect 14968 35198 15340 35204
rect 15968 35198 16340 35204
rect 16968 35198 17340 35204
rect 17968 35198 18340 35204
rect 18968 35198 19340 35204
rect 19968 35198 20340 35204
rect 20968 35198 21340 35204
rect 21968 35198 22340 35204
rect 22968 35198 23340 35204
rect 23968 35198 24340 35204
rect 24968 35198 25340 35204
rect 25968 35198 26340 35204
rect 26968 35198 27340 35204
rect 27968 35198 28340 35204
rect 28968 35198 29340 35204
rect 29968 35198 30340 35204
rect 30968 35198 31340 35204
rect 31968 35198 32340 35204
rect 32968 35198 33340 35204
rect 33968 35198 34340 35204
rect 9968 34902 10006 35198
rect 10302 34902 10340 35198
rect 10968 34902 11006 35198
rect 11302 34902 11340 35198
rect 11968 34902 12006 35198
rect 12302 34902 12340 35198
rect 12968 34902 13006 35198
rect 13302 34902 13340 35198
rect 13968 34902 14006 35198
rect 14302 34902 14340 35198
rect 14968 34902 15006 35198
rect 15302 34902 15340 35198
rect 15968 34902 16006 35198
rect 16302 34902 16340 35198
rect 16968 34902 17006 35198
rect 17302 34902 17340 35198
rect 17968 34902 18006 35198
rect 18302 34902 18340 35198
rect 18968 34902 19006 35198
rect 19302 34902 19340 35198
rect 19968 34902 20006 35198
rect 20302 34902 20340 35198
rect 20968 34902 21006 35198
rect 21302 34902 21340 35198
rect 21968 34902 22006 35198
rect 22302 34902 22340 35198
rect 22968 34902 23006 35198
rect 23302 34902 23340 35198
rect 23968 34902 24006 35198
rect 24302 34902 24340 35198
rect 24968 34902 25006 35198
rect 25302 34902 25340 35198
rect 25968 34902 26006 35198
rect 26302 34902 26340 35198
rect 26968 34902 27006 35198
rect 27302 34902 27340 35198
rect 27968 34902 28006 35198
rect 28302 34902 28340 35198
rect 28968 34902 29006 35198
rect 29302 34902 29340 35198
rect 29968 34902 30006 35198
rect 30302 34902 30340 35198
rect 30968 34902 31006 35198
rect 31302 34902 31340 35198
rect 31968 34902 32006 35198
rect 32302 34902 32340 35198
rect 32968 34902 33006 35198
rect 33302 34902 33340 35198
rect 33968 34902 34006 35198
rect 34302 34902 34340 35198
rect 9968 34896 10340 34902
rect 10968 34896 11340 34902
rect 11968 34896 12340 34902
rect 12968 34896 13340 34902
rect 13968 34896 14340 34902
rect 14968 34896 15340 34902
rect 15968 34896 16340 34902
rect 16968 34896 17340 34902
rect 17968 34896 18340 34902
rect 18968 34896 19340 34902
rect 19968 34896 20340 34902
rect 20968 34896 21340 34902
rect 21968 34896 22340 34902
rect 22968 34896 23340 34902
rect 23968 34896 24340 34902
rect 24968 34896 25340 34902
rect 25968 34896 26340 34902
rect 26968 34896 27340 34902
rect 27968 34896 28340 34902
rect 28968 34896 29340 34902
rect 29968 34896 30340 34902
rect 30968 34896 31340 34902
rect 31968 34896 32340 34902
rect 32968 34896 33340 34902
rect 33968 34896 34340 34902
rect 34648 34896 34654 35204
rect 9654 34890 34654 34896
rect -74485 34864 -74165 34890
rect -74485 34236 -74479 34864
rect -74171 34236 -74165 34864
rect -74485 34210 -74165 34236
rect -73485 34864 -73165 34890
rect -73485 34236 -73479 34864
rect -73171 34236 -73165 34864
rect -73485 34210 -73165 34236
rect -72485 34864 -72165 34890
rect -72485 34236 -72479 34864
rect -72171 34236 -72165 34864
rect -72485 34210 -72165 34236
rect -71485 34864 -71165 34890
rect -71485 34236 -71479 34864
rect -71171 34236 -71165 34864
rect -71485 34210 -71165 34236
rect -70485 34864 -70165 34890
rect -70485 34236 -70479 34864
rect -70171 34236 -70165 34864
rect -70485 34210 -70165 34236
rect -69485 34864 -69165 34890
rect -69485 34236 -69479 34864
rect -69171 34236 -69165 34864
rect -69485 34210 -69165 34236
rect -68485 34864 -68165 34890
rect -68485 34236 -68479 34864
rect -68171 34236 -68165 34864
rect -68485 34210 -68165 34236
rect -67485 34864 -67165 34890
rect -67485 34236 -67479 34864
rect -67171 34236 -67165 34864
rect -67485 34210 -67165 34236
rect -66485 34864 -66165 34890
rect -66485 34236 -66479 34864
rect -66171 34236 -66165 34864
rect -66485 34210 -66165 34236
rect -65485 34864 -65165 34890
rect -65485 34236 -65479 34864
rect -65171 34236 -65165 34864
rect -65485 34210 -65165 34236
rect -64485 34864 -64165 34890
rect -64485 34236 -64479 34864
rect -64171 34236 -64165 34864
rect -64485 34210 -64165 34236
rect -63485 34864 -63165 34890
rect -63485 34236 -63479 34864
rect -63171 34236 -63165 34864
rect -63485 34210 -63165 34236
rect -62485 34864 -62165 34890
rect -62485 34236 -62479 34864
rect -62171 34236 -62165 34864
rect -62485 34210 -62165 34236
rect -61485 34864 -61165 34890
rect -61485 34236 -61479 34864
rect -61171 34236 -61165 34864
rect -61485 34210 -61165 34236
rect -60485 34864 -60165 34890
rect -60485 34236 -60479 34864
rect -60171 34236 -60165 34864
rect -60485 34210 -60165 34236
rect -59485 34864 -59165 34890
rect -59485 34236 -59479 34864
rect -59171 34236 -59165 34864
rect -59485 34210 -59165 34236
rect 9994 34864 10314 34890
rect 9994 34236 10000 34864
rect 10308 34236 10314 34864
rect 9994 34210 10314 34236
rect 10994 34864 11314 34890
rect 10994 34236 11000 34864
rect 11308 34236 11314 34864
rect 10994 34210 11314 34236
rect 11994 34864 12314 34890
rect 11994 34236 12000 34864
rect 12308 34236 12314 34864
rect 11994 34210 12314 34236
rect 12994 34864 13314 34890
rect 12994 34236 13000 34864
rect 13308 34236 13314 34864
rect 12994 34210 13314 34236
rect 13994 34864 14314 34890
rect 13994 34236 14000 34864
rect 14308 34236 14314 34864
rect 13994 34210 14314 34236
rect 14994 34864 15314 34890
rect 14994 34236 15000 34864
rect 15308 34236 15314 34864
rect 14994 34210 15314 34236
rect 15994 34864 16314 34890
rect 15994 34236 16000 34864
rect 16308 34236 16314 34864
rect 15994 34210 16314 34236
rect 16994 34864 17314 34890
rect 16994 34236 17000 34864
rect 17308 34236 17314 34864
rect 16994 34210 17314 34236
rect 17994 34864 18314 34890
rect 17994 34236 18000 34864
rect 18308 34236 18314 34864
rect 17994 34210 18314 34236
rect 18994 34864 19314 34890
rect 18994 34236 19000 34864
rect 19308 34236 19314 34864
rect 18994 34210 19314 34236
rect 19994 34864 20314 34890
rect 19994 34236 20000 34864
rect 20308 34236 20314 34864
rect 19994 34210 20314 34236
rect 20994 34864 21314 34890
rect 20994 34236 21000 34864
rect 21308 34236 21314 34864
rect 20994 34210 21314 34236
rect 21994 34864 22314 34890
rect 21994 34236 22000 34864
rect 22308 34236 22314 34864
rect 21994 34210 22314 34236
rect 22994 34864 23314 34890
rect 22994 34236 23000 34864
rect 23308 34236 23314 34864
rect 22994 34210 23314 34236
rect 23994 34864 24314 34890
rect 23994 34236 24000 34864
rect 24308 34236 24314 34864
rect 23994 34210 24314 34236
rect 24994 34864 25314 34890
rect 24994 34236 25000 34864
rect 25308 34236 25314 34864
rect 24994 34210 25314 34236
rect 25994 34864 26314 34890
rect 25994 34236 26000 34864
rect 26308 34236 26314 34864
rect 25994 34210 26314 34236
rect 26994 34864 27314 34890
rect 26994 34236 27000 34864
rect 27308 34236 27314 34864
rect 26994 34210 27314 34236
rect 27994 34864 28314 34890
rect 27994 34236 28000 34864
rect 28308 34236 28314 34864
rect 27994 34210 28314 34236
rect 28994 34864 29314 34890
rect 28994 34236 29000 34864
rect 29308 34236 29314 34864
rect 28994 34210 29314 34236
rect 29994 34864 30314 34890
rect 29994 34236 30000 34864
rect 30308 34236 30314 34864
rect 29994 34210 30314 34236
rect 30994 34864 31314 34890
rect 30994 34236 31000 34864
rect 31308 34236 31314 34864
rect 30994 34210 31314 34236
rect 31994 34864 32314 34890
rect 31994 34236 32000 34864
rect 32308 34236 32314 34864
rect 31994 34210 32314 34236
rect 32994 34864 33314 34890
rect 32994 34236 33000 34864
rect 33308 34236 33314 34864
rect 32994 34210 33314 34236
rect 33994 34864 34314 34890
rect 33994 34236 34000 34864
rect 34308 34236 34314 34864
rect 33994 34210 34314 34236
rect -74825 34204 -58825 34210
rect -74825 33896 -74819 34204
rect -74511 34198 -74139 34204
rect -73511 34198 -73139 34204
rect -72511 34198 -72139 34204
rect -71511 34198 -71139 34204
rect -70511 34198 -70139 34204
rect -69511 34198 -69139 34204
rect -68511 34198 -68139 34204
rect -67511 34198 -67139 34204
rect -66511 34198 -66139 34204
rect -65511 34198 -65139 34204
rect -64511 34198 -64139 34204
rect -63511 34198 -63139 34204
rect -62511 34198 -62139 34204
rect -61511 34198 -61139 34204
rect -60511 34198 -60139 34204
rect -59511 34198 -59139 34204
rect -74511 33902 -74473 34198
rect -74177 33902 -74139 34198
rect -73511 33902 -73473 34198
rect -73177 33902 -73139 34198
rect -72511 33902 -72473 34198
rect -72177 33902 -72139 34198
rect -71511 33902 -71473 34198
rect -71177 33902 -71139 34198
rect -70511 33902 -70473 34198
rect -70177 33902 -70139 34198
rect -69511 33902 -69473 34198
rect -69177 33902 -69139 34198
rect -68511 33902 -68473 34198
rect -68177 33902 -68139 34198
rect -67511 33902 -67473 34198
rect -67177 33902 -67139 34198
rect -66511 33902 -66473 34198
rect -66177 33902 -66139 34198
rect -65511 33902 -65473 34198
rect -65177 33902 -65139 34198
rect -64511 33902 -64473 34198
rect -64177 33902 -64139 34198
rect -63511 33902 -63473 34198
rect -63177 33902 -63139 34198
rect -62511 33902 -62473 34198
rect -62177 33902 -62139 34198
rect -61511 33902 -61473 34198
rect -61177 33902 -61139 34198
rect -60511 33902 -60473 34198
rect -60177 33902 -60139 34198
rect -59511 33902 -59473 34198
rect -59177 33902 -59139 34198
rect -74511 33896 -74139 33902
rect -73511 33896 -73139 33902
rect -72511 33896 -72139 33902
rect -71511 33896 -71139 33902
rect -70511 33896 -70139 33902
rect -69511 33896 -69139 33902
rect -68511 33896 -68139 33902
rect -67511 33896 -67139 33902
rect -66511 33896 -66139 33902
rect -65511 33896 -65139 33902
rect -64511 33896 -64139 33902
rect -63511 33896 -63139 33902
rect -62511 33896 -62139 33902
rect -61511 33896 -61139 33902
rect -60511 33896 -60139 33902
rect -59511 33896 -59139 33902
rect -58831 33896 -58825 34204
rect 9654 34204 34654 34210
rect -74825 33890 -58825 33896
rect -50472 34170 -48808 34176
rect -74485 33864 -74165 33890
rect -74485 33236 -74479 33864
rect -74171 33236 -74165 33864
rect -74485 33210 -74165 33236
rect -73485 33864 -73165 33890
rect -73485 33236 -73479 33864
rect -73171 33236 -73165 33864
rect -73485 33210 -73165 33236
rect -72485 33864 -72165 33890
rect -72485 33236 -72479 33864
rect -72171 33236 -72165 33864
rect -72485 33210 -72165 33236
rect -71485 33864 -71165 33890
rect -71485 33236 -71479 33864
rect -71171 33236 -71165 33864
rect -71485 33210 -71165 33236
rect -70485 33864 -70165 33890
rect -70485 33236 -70479 33864
rect -70171 33236 -70165 33864
rect -70485 33210 -70165 33236
rect -69485 33864 -69165 33890
rect -69485 33236 -69479 33864
rect -69171 33236 -69165 33864
rect -69485 33210 -69165 33236
rect -68485 33864 -68165 33890
rect -68485 33236 -68479 33864
rect -68171 33236 -68165 33864
rect -68485 33210 -68165 33236
rect -67485 33864 -67165 33890
rect -67485 33236 -67479 33864
rect -67171 33236 -67165 33864
rect -67485 33210 -67165 33236
rect -66485 33864 -66165 33890
rect -66485 33236 -66479 33864
rect -66171 33236 -66165 33864
rect -66485 33210 -66165 33236
rect -65485 33864 -65165 33890
rect -65485 33236 -65479 33864
rect -65171 33236 -65165 33864
rect -65485 33210 -65165 33236
rect -64485 33864 -64165 33890
rect -64485 33236 -64479 33864
rect -64171 33236 -64165 33864
rect -64485 33210 -64165 33236
rect -63485 33864 -63165 33890
rect -63485 33236 -63479 33864
rect -63171 33236 -63165 33864
rect -63485 33210 -63165 33236
rect -62485 33864 -62165 33890
rect -62485 33236 -62479 33864
rect -62171 33236 -62165 33864
rect -62485 33210 -62165 33236
rect -61485 33864 -61165 33890
rect -61485 33236 -61479 33864
rect -61171 33236 -61165 33864
rect -61485 33210 -61165 33236
rect -60485 33864 -60165 33890
rect -60485 33236 -60479 33864
rect -60171 33236 -60165 33864
rect -60485 33210 -60165 33236
rect -59485 33864 -59165 33890
rect -59485 33236 -59479 33864
rect -59171 33236 -59165 33864
rect -50472 33542 -50466 34170
rect -48814 33542 -48808 34170
rect -50472 33536 -48808 33542
rect 2875 34170 4539 34176
rect 2875 33542 2881 34170
rect 4533 33542 4539 34170
rect 9654 33896 9660 34204
rect 9968 34198 10340 34204
rect 10968 34198 11340 34204
rect 11968 34198 12340 34204
rect 12968 34198 13340 34204
rect 13968 34198 14340 34204
rect 14968 34198 15340 34204
rect 15968 34198 16340 34204
rect 16968 34198 17340 34204
rect 17968 34198 18340 34204
rect 18968 34198 19340 34204
rect 19968 34198 20340 34204
rect 20968 34198 21340 34204
rect 21968 34198 22340 34204
rect 22968 34198 23340 34204
rect 23968 34198 24340 34204
rect 24968 34198 25340 34204
rect 25968 34198 26340 34204
rect 26968 34198 27340 34204
rect 27968 34198 28340 34204
rect 28968 34198 29340 34204
rect 29968 34198 30340 34204
rect 30968 34198 31340 34204
rect 31968 34198 32340 34204
rect 32968 34198 33340 34204
rect 33968 34198 34340 34204
rect 9968 33902 10006 34198
rect 10302 33902 10340 34198
rect 10968 33902 11006 34198
rect 11302 33902 11340 34198
rect 11968 33902 12006 34198
rect 12302 33902 12340 34198
rect 12968 33902 13006 34198
rect 13302 33902 13340 34198
rect 13968 33902 14006 34198
rect 14302 33902 14340 34198
rect 14968 33902 15006 34198
rect 15302 33902 15340 34198
rect 15968 33902 16006 34198
rect 16302 33902 16340 34198
rect 16968 33902 17006 34198
rect 17302 33902 17340 34198
rect 17968 33902 18006 34198
rect 18302 33902 18340 34198
rect 18968 33902 19006 34198
rect 19302 33902 19340 34198
rect 19968 33902 20006 34198
rect 20302 33902 20340 34198
rect 20968 33902 21006 34198
rect 21302 33902 21340 34198
rect 21968 33902 22006 34198
rect 22302 33902 22340 34198
rect 22968 33902 23006 34198
rect 23302 33902 23340 34198
rect 23968 33902 24006 34198
rect 24302 33902 24340 34198
rect 24968 33902 25006 34198
rect 25302 33902 25340 34198
rect 25968 33902 26006 34198
rect 26302 33902 26340 34198
rect 26968 33902 27006 34198
rect 27302 33902 27340 34198
rect 27968 33902 28006 34198
rect 28302 33902 28340 34198
rect 28968 33902 29006 34198
rect 29302 33902 29340 34198
rect 29968 33902 30006 34198
rect 30302 33902 30340 34198
rect 30968 33902 31006 34198
rect 31302 33902 31340 34198
rect 31968 33902 32006 34198
rect 32302 33902 32340 34198
rect 32968 33902 33006 34198
rect 33302 33902 33340 34198
rect 33968 33902 34006 34198
rect 34302 33902 34340 34198
rect 9968 33896 10340 33902
rect 10968 33896 11340 33902
rect 11968 33896 12340 33902
rect 12968 33896 13340 33902
rect 13968 33896 14340 33902
rect 14968 33896 15340 33902
rect 15968 33896 16340 33902
rect 16968 33896 17340 33902
rect 17968 33896 18340 33902
rect 18968 33896 19340 33902
rect 19968 33896 20340 33902
rect 20968 33896 21340 33902
rect 21968 33896 22340 33902
rect 22968 33896 23340 33902
rect 23968 33896 24340 33902
rect 24968 33896 25340 33902
rect 25968 33896 26340 33902
rect 26968 33896 27340 33902
rect 27968 33896 28340 33902
rect 28968 33896 29340 33902
rect 29968 33896 30340 33902
rect 30968 33896 31340 33902
rect 31968 33896 32340 33902
rect 32968 33896 33340 33902
rect 33968 33896 34340 33902
rect 34648 33896 34654 34204
rect 9654 33890 34654 33896
rect 2875 33536 4539 33542
rect 9994 33864 10314 33890
rect -59485 33210 -59165 33236
rect -50304 33298 -48430 33304
rect -50304 33246 -50298 33298
rect -50246 33246 -49982 33298
rect -49930 33246 -49666 33298
rect -49614 33246 -49350 33298
rect -49298 33246 -49034 33298
rect -48982 33246 -48430 33298
rect -50304 33234 -48430 33246
rect -74825 33204 -58825 33210
rect -74825 32896 -74819 33204
rect -74511 33198 -74139 33204
rect -73511 33198 -73139 33204
rect -72511 33198 -72139 33204
rect -71511 33198 -71139 33204
rect -70511 33198 -70139 33204
rect -69511 33198 -69139 33204
rect -68511 33198 -68139 33204
rect -67511 33198 -67139 33204
rect -66511 33198 -66139 33204
rect -65511 33198 -65139 33204
rect -64511 33198 -64139 33204
rect -63511 33198 -63139 33204
rect -62511 33198 -62139 33204
rect -61511 33198 -61139 33204
rect -60511 33198 -60139 33204
rect -59511 33198 -59139 33204
rect -74511 32902 -74473 33198
rect -74177 32902 -74139 33198
rect -73511 32902 -73473 33198
rect -73177 32902 -73139 33198
rect -72511 32902 -72473 33198
rect -72177 32902 -72139 33198
rect -71511 32902 -71473 33198
rect -71177 32902 -71139 33198
rect -70511 32902 -70473 33198
rect -70177 32902 -70139 33198
rect -69511 32902 -69473 33198
rect -69177 32902 -69139 33198
rect -68511 32902 -68473 33198
rect -68177 32902 -68139 33198
rect -67511 32902 -67473 33198
rect -67177 32902 -67139 33198
rect -66511 32902 -66473 33198
rect -66177 32902 -66139 33198
rect -65511 32902 -65473 33198
rect -65177 32902 -65139 33198
rect -64511 32902 -64473 33198
rect -64177 32902 -64139 33198
rect -63511 32902 -63473 33198
rect -63177 32902 -63139 33198
rect -62511 32902 -62473 33198
rect -62177 32902 -62139 33198
rect -61511 32902 -61473 33198
rect -61177 32902 -61139 33198
rect -60511 32902 -60473 33198
rect -60177 32902 -60139 33198
rect -59511 32902 -59473 33198
rect -59177 32902 -59139 33198
rect -74511 32896 -74139 32902
rect -73511 32896 -73139 32902
rect -72511 32896 -72139 32902
rect -71511 32896 -71139 32902
rect -70511 32896 -70139 32902
rect -69511 32896 -69139 32902
rect -68511 32896 -68139 32902
rect -67511 32896 -67139 32902
rect -66511 32896 -66139 32902
rect -65511 32896 -65139 32902
rect -64511 32896 -64139 32902
rect -63511 32896 -63139 32902
rect -62511 32896 -62139 32902
rect -61511 32896 -61139 32902
rect -60511 32896 -60139 32902
rect -59511 32896 -59139 32902
rect -58831 32896 -58825 33204
rect -50304 33182 -50298 33234
rect -50246 33182 -49982 33234
rect -49930 33182 -49666 33234
rect -49614 33182 -49350 33234
rect -49298 33182 -49034 33234
rect -48982 33184 -48430 33234
rect 3043 33298 7220 33304
rect 3043 33246 3049 33298
rect 3101 33246 3365 33298
rect 3417 33246 3681 33298
rect 3733 33246 3997 33298
rect 4049 33246 4313 33298
rect 4365 33246 7220 33298
rect 3043 33234 7220 33246
rect -48982 33182 2774 33184
rect -50304 33170 2774 33182
rect -50304 33118 -50298 33170
rect -50246 33118 -49982 33170
rect -49930 33118 -49666 33170
rect -49614 33118 -49350 33170
rect -49298 33118 -49034 33170
rect -48982 33118 2774 33170
rect -50304 33106 2774 33118
rect -50304 33054 -50298 33106
rect -50246 33054 -49982 33106
rect -49930 33054 -49666 33106
rect -49614 33054 -49350 33106
rect -49298 33054 -49034 33106
rect -48982 33054 2774 33106
rect -50304 33042 2774 33054
rect -50304 32990 -50298 33042
rect -50246 32990 -49982 33042
rect -49930 32990 -49666 33042
rect -49614 32990 -49350 33042
rect -49298 32990 -49034 33042
rect -48982 32990 2774 33042
rect -50304 32978 2774 32990
rect -74825 32890 -58825 32896
rect -50964 32967 -50570 32976
rect -74485 32864 -74165 32890
rect -74485 32236 -74479 32864
rect -74171 32236 -74165 32864
rect -74485 32210 -74165 32236
rect -73485 32864 -73165 32890
rect -73485 32236 -73479 32864
rect -73171 32236 -73165 32864
rect -73485 32210 -73165 32236
rect -72485 32864 -72165 32890
rect -72485 32236 -72479 32864
rect -72171 32236 -72165 32864
rect -72485 32210 -72165 32236
rect -71485 32864 -71165 32890
rect -71485 32236 -71479 32864
rect -71171 32236 -71165 32864
rect -71485 32210 -71165 32236
rect -70485 32864 -70165 32890
rect -70485 32236 -70479 32864
rect -70171 32236 -70165 32864
rect -70485 32210 -70165 32236
rect -69485 32864 -69165 32890
rect -69485 32236 -69479 32864
rect -69171 32236 -69165 32864
rect -69485 32210 -69165 32236
rect -68485 32864 -68165 32890
rect -68485 32236 -68479 32864
rect -68171 32236 -68165 32864
rect -68485 32210 -68165 32236
rect -67485 32864 -67165 32890
rect -67485 32236 -67479 32864
rect -67171 32236 -67165 32864
rect -67485 32210 -67165 32236
rect -66485 32864 -66165 32890
rect -66485 32236 -66479 32864
rect -66171 32236 -66165 32864
rect -66485 32210 -66165 32236
rect -65485 32864 -65165 32890
rect -65485 32236 -65479 32864
rect -65171 32236 -65165 32864
rect -65485 32210 -65165 32236
rect -64485 32864 -64165 32890
rect -64485 32236 -64479 32864
rect -64171 32236 -64165 32864
rect -64485 32210 -64165 32236
rect -63485 32864 -63165 32890
rect -63485 32236 -63479 32864
rect -63171 32236 -63165 32864
rect -63485 32210 -63165 32236
rect -62485 32864 -62165 32890
rect -62485 32236 -62479 32864
rect -62171 32236 -62165 32864
rect -62485 32210 -62165 32236
rect -61485 32864 -61165 32890
rect -61485 32236 -61479 32864
rect -61171 32236 -61165 32864
rect -61485 32210 -61165 32236
rect -60485 32864 -60165 32890
rect -60485 32236 -60479 32864
rect -60171 32236 -60165 32864
rect -60485 32210 -60165 32236
rect -59485 32864 -59165 32890
rect -59485 32236 -59479 32864
rect -59171 32236 -59165 32864
rect -50964 32591 -50955 32967
rect -50579 32591 -50570 32967
rect -50304 32926 -50298 32978
rect -50246 32926 -49982 32978
rect -49930 32926 -49666 32978
rect -49614 32926 -49350 32978
rect -49298 32926 -49034 32978
rect -48982 32965 2774 32978
rect -48982 32926 2396 32965
rect -50304 32920 2396 32926
rect -48721 32651 2396 32920
rect -50964 32582 -50570 32591
rect -50304 32645 2396 32651
rect -50304 32593 -50298 32645
rect -50246 32593 -49982 32645
rect -49930 32593 -49666 32645
rect -49614 32593 -49350 32645
rect -49298 32593 -49034 32645
rect -48982 32593 2396 32645
rect 2768 32593 2774 32965
rect 3043 33182 3049 33234
rect 3101 33182 3365 33234
rect 3417 33182 3681 33234
rect 3733 33182 3997 33234
rect 4049 33182 4313 33234
rect 4365 33182 7220 33234
rect 9994 33236 10000 33864
rect 10308 33236 10314 33864
rect 9994 33210 10314 33236
rect 10994 33864 11314 33890
rect 10994 33236 11000 33864
rect 11308 33236 11314 33864
rect 10994 33210 11314 33236
rect 11994 33864 12314 33890
rect 11994 33236 12000 33864
rect 12308 33236 12314 33864
rect 11994 33210 12314 33236
rect 12994 33864 13314 33890
rect 12994 33236 13000 33864
rect 13308 33236 13314 33864
rect 12994 33210 13314 33236
rect 13994 33864 14314 33890
rect 13994 33236 14000 33864
rect 14308 33236 14314 33864
rect 13994 33210 14314 33236
rect 14994 33864 15314 33890
rect 14994 33236 15000 33864
rect 15308 33236 15314 33864
rect 14994 33210 15314 33236
rect 15994 33864 16314 33890
rect 15994 33236 16000 33864
rect 16308 33236 16314 33864
rect 15994 33210 16314 33236
rect 16994 33864 17314 33890
rect 16994 33236 17000 33864
rect 17308 33236 17314 33864
rect 16994 33210 17314 33236
rect 17994 33864 18314 33890
rect 17994 33236 18000 33864
rect 18308 33236 18314 33864
rect 17994 33210 18314 33236
rect 18994 33864 19314 33890
rect 18994 33236 19000 33864
rect 19308 33236 19314 33864
rect 18994 33210 19314 33236
rect 19994 33864 20314 33890
rect 19994 33236 20000 33864
rect 20308 33236 20314 33864
rect 19994 33210 20314 33236
rect 20994 33864 21314 33890
rect 20994 33236 21000 33864
rect 21308 33236 21314 33864
rect 20994 33210 21314 33236
rect 21994 33864 22314 33890
rect 21994 33236 22000 33864
rect 22308 33236 22314 33864
rect 21994 33210 22314 33236
rect 22994 33864 23314 33890
rect 22994 33236 23000 33864
rect 23308 33236 23314 33864
rect 22994 33210 23314 33236
rect 23994 33864 24314 33890
rect 23994 33236 24000 33864
rect 24308 33236 24314 33864
rect 23994 33210 24314 33236
rect 24994 33864 25314 33890
rect 24994 33236 25000 33864
rect 25308 33236 25314 33864
rect 24994 33210 25314 33236
rect 25994 33864 26314 33890
rect 25994 33236 26000 33864
rect 26308 33236 26314 33864
rect 25994 33210 26314 33236
rect 26994 33864 27314 33890
rect 26994 33236 27000 33864
rect 27308 33236 27314 33864
rect 26994 33210 27314 33236
rect 27994 33864 28314 33890
rect 27994 33236 28000 33864
rect 28308 33236 28314 33864
rect 27994 33210 28314 33236
rect 28994 33864 29314 33890
rect 28994 33236 29000 33864
rect 29308 33236 29314 33864
rect 28994 33210 29314 33236
rect 29994 33864 30314 33890
rect 29994 33236 30000 33864
rect 30308 33236 30314 33864
rect 29994 33210 30314 33236
rect 30994 33864 31314 33890
rect 30994 33236 31000 33864
rect 31308 33236 31314 33864
rect 30994 33210 31314 33236
rect 31994 33864 32314 33890
rect 31994 33236 32000 33864
rect 32308 33236 32314 33864
rect 31994 33210 32314 33236
rect 32994 33864 33314 33890
rect 32994 33236 33000 33864
rect 33308 33236 33314 33864
rect 32994 33210 33314 33236
rect 33994 33864 34314 33890
rect 33994 33236 34000 33864
rect 34308 33236 34314 33864
rect 33994 33210 34314 33236
rect 3043 33170 7220 33182
rect 3043 33118 3049 33170
rect 3101 33118 3365 33170
rect 3417 33118 3681 33170
rect 3733 33118 3997 33170
rect 4049 33118 4313 33170
rect 4365 33118 7220 33170
rect 3043 33106 7220 33118
rect 3043 33054 3049 33106
rect 3101 33054 3365 33106
rect 3417 33054 3681 33106
rect 3733 33054 3997 33106
rect 4049 33054 4313 33106
rect 4365 33054 7220 33106
rect 3043 33042 7220 33054
rect 3043 32990 3049 33042
rect 3101 32990 3365 33042
rect 3417 32990 3681 33042
rect 3733 32990 3997 33042
rect 4049 32990 4313 33042
rect 4365 32990 7220 33042
rect 3043 32978 7220 32990
rect 3043 32926 3049 32978
rect 3101 32926 3365 32978
rect 3417 32926 3681 32978
rect 3733 32926 3997 32978
rect 4049 32926 4313 32978
rect 4365 32926 7220 32978
rect 3043 32920 7220 32926
rect 4626 32704 7220 32920
rect 9654 33204 34654 33210
rect 9654 32896 9660 33204
rect 9968 33198 10340 33204
rect 10968 33198 11340 33204
rect 11968 33198 12340 33204
rect 12968 33198 13340 33204
rect 13968 33198 14340 33204
rect 14968 33198 15340 33204
rect 15968 33198 16340 33204
rect 16968 33198 17340 33204
rect 17968 33198 18340 33204
rect 18968 33198 19340 33204
rect 19968 33198 20340 33204
rect 20968 33198 21340 33204
rect 21968 33198 22340 33204
rect 22968 33198 23340 33204
rect 23968 33198 24340 33204
rect 24968 33198 25340 33204
rect 25968 33198 26340 33204
rect 26968 33198 27340 33204
rect 27968 33198 28340 33204
rect 28968 33198 29340 33204
rect 29968 33198 30340 33204
rect 30968 33198 31340 33204
rect 31968 33198 32340 33204
rect 32968 33198 33340 33204
rect 33968 33198 34340 33204
rect 9968 32902 10006 33198
rect 10302 32902 10340 33198
rect 10968 32902 11006 33198
rect 11302 32902 11340 33198
rect 11968 32902 12006 33198
rect 12302 32902 12340 33198
rect 12968 32902 13006 33198
rect 13302 32902 13340 33198
rect 13968 32902 14006 33198
rect 14302 32902 14340 33198
rect 14968 32902 15006 33198
rect 15302 32902 15340 33198
rect 15968 32902 16006 33198
rect 16302 32902 16340 33198
rect 16968 32902 17006 33198
rect 17302 32902 17340 33198
rect 17968 32902 18006 33198
rect 18302 32902 18340 33198
rect 18968 32902 19006 33198
rect 19302 32902 19340 33198
rect 19968 32902 20006 33198
rect 20302 32902 20340 33198
rect 20968 32902 21006 33198
rect 21302 32902 21340 33198
rect 21968 32902 22006 33198
rect 22302 32902 22340 33198
rect 22968 32902 23006 33198
rect 23302 32902 23340 33198
rect 23968 32902 24006 33198
rect 24302 32902 24340 33198
rect 24968 32902 25006 33198
rect 25302 32902 25340 33198
rect 25968 32902 26006 33198
rect 26302 32902 26340 33198
rect 26968 32902 27006 33198
rect 27302 32902 27340 33198
rect 27968 32902 28006 33198
rect 28302 32902 28340 33198
rect 28968 32902 29006 33198
rect 29302 32902 29340 33198
rect 29968 32902 30006 33198
rect 30302 32902 30340 33198
rect 30968 32902 31006 33198
rect 31302 32902 31340 33198
rect 31968 32902 32006 33198
rect 32302 32902 32340 33198
rect 32968 32902 33006 33198
rect 33302 32902 33340 33198
rect 33968 32902 34006 33198
rect 34302 32902 34340 33198
rect 9968 32896 10340 32902
rect 10968 32896 11340 32902
rect 11968 32896 12340 32902
rect 12968 32896 13340 32902
rect 13968 32896 14340 32902
rect 14968 32896 15340 32902
rect 15968 32896 16340 32902
rect 16968 32896 17340 32902
rect 17968 32896 18340 32902
rect 18968 32896 19340 32902
rect 19968 32896 20340 32902
rect 20968 32896 21340 32902
rect 21968 32896 22340 32902
rect 22968 32896 23340 32902
rect 23968 32896 24340 32902
rect 24968 32896 25340 32902
rect 25968 32896 26340 32902
rect 26968 32896 27340 32902
rect 27968 32896 28340 32902
rect 28968 32896 29340 32902
rect 29968 32896 30340 32902
rect 30968 32896 31340 32902
rect 31968 32896 32340 32902
rect 32968 32896 33340 32902
rect 33968 32896 34340 32902
rect 34648 32896 34654 33204
rect 9654 32890 34654 32896
rect 4626 32651 4917 32704
rect -50304 32584 2774 32593
rect 3043 32645 4917 32651
rect 3043 32593 3049 32645
rect 3101 32593 3365 32645
rect 3417 32593 3681 32645
rect 3733 32593 3997 32645
rect 4049 32593 4313 32645
rect 4365 32593 4917 32645
rect -50304 32581 -48430 32584
rect -50304 32529 -50298 32581
rect -50246 32529 -49982 32581
rect -49930 32529 -49666 32581
rect -49614 32529 -49350 32581
rect -49298 32529 -49034 32581
rect -48982 32529 -48430 32581
rect -50304 32517 -48430 32529
rect -50304 32465 -50298 32517
rect -50246 32465 -49982 32517
rect -49930 32465 -49666 32517
rect -49614 32465 -49350 32517
rect -49298 32465 -49034 32517
rect -48982 32465 -48430 32517
rect -50304 32459 -48430 32465
rect -59485 32210 -59165 32236
rect -74825 32204 -58825 32210
rect -74825 31896 -74819 32204
rect -74511 32198 -74139 32204
rect -73511 32198 -73139 32204
rect -72511 32198 -72139 32204
rect -71511 32198 -71139 32204
rect -70511 32198 -70139 32204
rect -69511 32198 -69139 32204
rect -68511 32198 -68139 32204
rect -67511 32198 -67139 32204
rect -66511 32198 -66139 32204
rect -65511 32198 -65139 32204
rect -64511 32198 -64139 32204
rect -63511 32198 -63139 32204
rect -62511 32198 -62139 32204
rect -61511 32198 -61139 32204
rect -60511 32198 -60139 32204
rect -59511 32198 -59139 32204
rect -74511 31902 -74473 32198
rect -74177 31902 -74139 32198
rect -73511 31902 -73473 32198
rect -73177 31902 -73139 32198
rect -72511 31902 -72473 32198
rect -72177 31902 -72139 32198
rect -71511 31902 -71473 32198
rect -71177 31902 -71139 32198
rect -70511 31902 -70473 32198
rect -70177 31902 -70139 32198
rect -69511 31902 -69473 32198
rect -69177 31902 -69139 32198
rect -68511 31902 -68473 32198
rect -68177 31902 -68139 32198
rect -67511 31902 -67473 32198
rect -67177 31902 -67139 32198
rect -66511 31902 -66473 32198
rect -66177 31902 -66139 32198
rect -65511 31902 -65473 32198
rect -65177 31902 -65139 32198
rect -64511 31902 -64473 32198
rect -64177 31902 -64139 32198
rect -63511 31902 -63473 32198
rect -63177 31902 -63139 32198
rect -62511 31902 -62473 32198
rect -62177 31902 -62139 32198
rect -61511 31902 -61473 32198
rect -61177 31902 -61139 32198
rect -60511 31902 -60473 32198
rect -60177 31902 -60139 32198
rect -59511 31902 -59473 32198
rect -59177 31902 -59139 32198
rect -74511 31896 -74139 31902
rect -73511 31896 -73139 31902
rect -72511 31896 -72139 31902
rect -71511 31896 -71139 31902
rect -70511 31896 -70139 31902
rect -69511 31896 -69139 31902
rect -68511 31896 -68139 31902
rect -67511 31896 -67139 31902
rect -66511 31896 -66139 31902
rect -65511 31896 -65139 31902
rect -64511 31896 -64139 31902
rect -63511 31896 -63139 31902
rect -62511 31896 -62139 31902
rect -61511 31896 -61139 31902
rect -60511 31896 -60139 31902
rect -59511 31896 -59139 31902
rect -58831 31896 -58825 32204
rect -74825 31890 -58825 31896
rect -74485 31864 -74165 31890
rect -74485 31236 -74479 31864
rect -74171 31236 -74165 31864
rect -74485 31210 -74165 31236
rect -73485 31864 -73165 31890
rect -73485 31236 -73479 31864
rect -73171 31236 -73165 31864
rect -73485 31210 -73165 31236
rect -72485 31864 -72165 31890
rect -72485 31236 -72479 31864
rect -72171 31236 -72165 31864
rect -72485 31210 -72165 31236
rect -71485 31864 -71165 31890
rect -71485 31236 -71479 31864
rect -71171 31236 -71165 31864
rect -71485 31210 -71165 31236
rect -70485 31864 -70165 31890
rect -70485 31236 -70479 31864
rect -70171 31236 -70165 31864
rect -70485 31210 -70165 31236
rect -69485 31864 -69165 31890
rect -69485 31236 -69479 31864
rect -69171 31236 -69165 31864
rect -69485 31210 -69165 31236
rect -68485 31864 -68165 31890
rect -68485 31236 -68479 31864
rect -68171 31236 -68165 31864
rect -68485 31210 -68165 31236
rect -67485 31864 -67165 31890
rect -67485 31236 -67479 31864
rect -67171 31236 -67165 31864
rect -67485 31210 -67165 31236
rect -66485 31864 -66165 31890
rect -66485 31236 -66479 31864
rect -66171 31236 -66165 31864
rect -66485 31210 -66165 31236
rect -65485 31864 -65165 31890
rect -65485 31236 -65479 31864
rect -65171 31236 -65165 31864
rect -65485 31210 -65165 31236
rect -64485 31864 -64165 31890
rect -64485 31236 -64479 31864
rect -64171 31236 -64165 31864
rect -64485 31210 -64165 31236
rect -63485 31864 -63165 31890
rect -63485 31236 -63479 31864
rect -63171 31236 -63165 31864
rect -63485 31210 -63165 31236
rect -62485 31864 -62165 31890
rect -62485 31236 -62479 31864
rect -62171 31236 -62165 31864
rect -62485 31210 -62165 31236
rect -61485 31864 -61165 31890
rect -61485 31236 -61479 31864
rect -61171 31236 -61165 31864
rect -61485 31210 -61165 31236
rect -60485 31864 -60165 31890
rect -60485 31236 -60479 31864
rect -60171 31236 -60165 31864
rect -60485 31210 -60165 31236
rect -59485 31864 -59165 31890
rect -59485 31236 -59479 31864
rect -59171 31236 -59165 31864
rect -59485 31210 -59165 31236
rect -74825 31204 -58825 31210
rect -74825 30896 -74819 31204
rect -74511 31198 -74139 31204
rect -73511 31198 -73139 31204
rect -72511 31198 -72139 31204
rect -71511 31198 -71139 31204
rect -70511 31198 -70139 31204
rect -69511 31198 -69139 31204
rect -68511 31198 -68139 31204
rect -67511 31198 -67139 31204
rect -66511 31198 -66139 31204
rect -65511 31198 -65139 31204
rect -64511 31198 -64139 31204
rect -63511 31198 -63139 31204
rect -62511 31198 -62139 31204
rect -61511 31198 -61139 31204
rect -60511 31198 -60139 31204
rect -59511 31198 -59139 31204
rect -74511 30902 -74473 31198
rect -74177 30902 -74139 31198
rect -73511 30902 -73473 31198
rect -73177 30902 -73139 31198
rect -72511 30902 -72473 31198
rect -72177 30902 -72139 31198
rect -71511 30902 -71473 31198
rect -71177 30902 -71139 31198
rect -70511 30902 -70473 31198
rect -70177 30902 -70139 31198
rect -69511 30902 -69473 31198
rect -69177 30902 -69139 31198
rect -68511 30902 -68473 31198
rect -68177 30902 -68139 31198
rect -67511 30902 -67473 31198
rect -67177 30902 -67139 31198
rect -66511 30902 -66473 31198
rect -66177 30902 -66139 31198
rect -65511 30902 -65473 31198
rect -65177 30902 -65139 31198
rect -64511 30902 -64473 31198
rect -64177 30902 -64139 31198
rect -63511 30902 -63473 31198
rect -63177 30902 -63139 31198
rect -62511 30902 -62473 31198
rect -62177 30902 -62139 31198
rect -61511 30902 -61473 31198
rect -61177 30902 -61139 31198
rect -60511 30902 -60473 31198
rect -60177 30902 -60139 31198
rect -59511 30902 -59473 31198
rect -59177 30902 -59139 31198
rect -74511 30896 -74139 30902
rect -73511 30896 -73139 30902
rect -72511 30896 -72139 30902
rect -71511 30896 -71139 30902
rect -70511 30896 -70139 30902
rect -69511 30896 -69139 30902
rect -68511 30896 -68139 30902
rect -67511 30896 -67139 30902
rect -66511 30896 -66139 30902
rect -65511 30896 -65139 30902
rect -64511 30896 -64139 30902
rect -63511 30896 -63139 30902
rect -62511 30896 -62139 30902
rect -61511 30896 -61139 30902
rect -60511 30896 -60139 30902
rect -59511 30896 -59139 30902
rect -58831 30896 -58825 31204
rect -74825 30890 -58825 30896
rect -74485 30864 -74165 30890
rect -74485 30236 -74479 30864
rect -74171 30236 -74165 30864
rect -74485 30210 -74165 30236
rect -73485 30864 -73165 30890
rect -73485 30236 -73479 30864
rect -73171 30236 -73165 30864
rect -73485 30210 -73165 30236
rect -72485 30864 -72165 30890
rect -72485 30236 -72479 30864
rect -72171 30236 -72165 30864
rect -72485 30210 -72165 30236
rect -71485 30864 -71165 30890
rect -71485 30236 -71479 30864
rect -71171 30236 -71165 30864
rect -71485 30210 -71165 30236
rect -70485 30864 -70165 30890
rect -70485 30236 -70479 30864
rect -70171 30236 -70165 30864
rect -70485 30210 -70165 30236
rect -69485 30864 -69165 30890
rect -69485 30236 -69479 30864
rect -69171 30236 -69165 30864
rect -69485 30210 -69165 30236
rect -68485 30864 -68165 30890
rect -68485 30236 -68479 30864
rect -68171 30236 -68165 30864
rect -68485 30210 -68165 30236
rect -67485 30864 -67165 30890
rect -67485 30236 -67479 30864
rect -67171 30236 -67165 30864
rect -67485 30210 -67165 30236
rect -66485 30864 -66165 30890
rect -66485 30236 -66479 30864
rect -66171 30236 -66165 30864
rect -66485 30210 -66165 30236
rect -65485 30864 -65165 30890
rect -65485 30236 -65479 30864
rect -65171 30236 -65165 30864
rect -65485 30210 -65165 30236
rect -64485 30864 -64165 30890
rect -64485 30236 -64479 30864
rect -64171 30236 -64165 30864
rect -64485 30210 -64165 30236
rect -63485 30864 -63165 30890
rect -63485 30236 -63479 30864
rect -63171 30236 -63165 30864
rect -63485 30210 -63165 30236
rect -62485 30864 -62165 30890
rect -62485 30236 -62479 30864
rect -62171 30236 -62165 30864
rect -62485 30210 -62165 30236
rect -61485 30864 -61165 30890
rect -61485 30236 -61479 30864
rect -61171 30236 -61165 30864
rect -61485 30210 -61165 30236
rect -60485 30864 -60165 30890
rect -60485 30236 -60479 30864
rect -60171 30236 -60165 30864
rect -60485 30210 -60165 30236
rect -59485 30864 -59165 30890
rect -59485 30236 -59479 30864
rect -59171 30236 -59165 30864
rect -59485 30210 -59165 30236
rect -74825 30204 -58825 30210
rect -74825 29896 -74819 30204
rect -74511 30198 -74139 30204
rect -73511 30198 -73139 30204
rect -72511 30198 -72139 30204
rect -71511 30198 -71139 30204
rect -70511 30198 -70139 30204
rect -69511 30198 -69139 30204
rect -68511 30198 -68139 30204
rect -67511 30198 -67139 30204
rect -66511 30198 -66139 30204
rect -65511 30198 -65139 30204
rect -64511 30198 -64139 30204
rect -63511 30198 -63139 30204
rect -62511 30198 -62139 30204
rect -61511 30198 -61139 30204
rect -60511 30198 -60139 30204
rect -59511 30198 -59139 30204
rect -74511 29902 -74473 30198
rect -74177 29902 -74139 30198
rect -73511 29902 -73473 30198
rect -73177 29902 -73139 30198
rect -72511 29902 -72473 30198
rect -72177 29902 -72139 30198
rect -71511 29902 -71473 30198
rect -71177 29902 -71139 30198
rect -70511 29902 -70473 30198
rect -70177 29902 -70139 30198
rect -69511 29902 -69473 30198
rect -69177 29902 -69139 30198
rect -68511 29902 -68473 30198
rect -68177 29902 -68139 30198
rect -67511 29902 -67473 30198
rect -67177 29902 -67139 30198
rect -66511 29902 -66473 30198
rect -66177 29902 -66139 30198
rect -65511 29902 -65473 30198
rect -65177 29902 -65139 30198
rect -64511 29902 -64473 30198
rect -64177 29902 -64139 30198
rect -63511 29902 -63473 30198
rect -63177 29902 -63139 30198
rect -62511 29902 -62473 30198
rect -62177 29902 -62139 30198
rect -61511 29902 -61473 30198
rect -61177 29902 -61139 30198
rect -60511 29902 -60473 30198
rect -60177 29902 -60139 30198
rect -59511 29902 -59473 30198
rect -59177 29902 -59139 30198
rect -74511 29896 -74139 29902
rect -73511 29896 -73139 29902
rect -72511 29896 -72139 29902
rect -71511 29896 -71139 29902
rect -70511 29896 -70139 29902
rect -69511 29896 -69139 29902
rect -68511 29896 -68139 29902
rect -67511 29896 -67139 29902
rect -66511 29896 -66139 29902
rect -65511 29896 -65139 29902
rect -64511 29896 -64139 29902
rect -63511 29896 -63139 29902
rect -62511 29896 -62139 29902
rect -61511 29896 -61139 29902
rect -60511 29896 -60139 29902
rect -59511 29896 -59139 29902
rect -58831 29896 -58825 30204
rect -74825 29890 -58825 29896
rect -74485 29864 -74165 29890
rect -74485 29236 -74479 29864
rect -74171 29236 -74165 29864
rect -74485 29210 -74165 29236
rect -73485 29864 -73165 29890
rect -73485 29236 -73479 29864
rect -73171 29236 -73165 29864
rect -73485 29210 -73165 29236
rect -72485 29864 -72165 29890
rect -72485 29236 -72479 29864
rect -72171 29236 -72165 29864
rect -72485 29210 -72165 29236
rect -71485 29864 -71165 29890
rect -71485 29236 -71479 29864
rect -71171 29236 -71165 29864
rect -71485 29210 -71165 29236
rect -70485 29864 -70165 29890
rect -70485 29236 -70479 29864
rect -70171 29236 -70165 29864
rect -70485 29210 -70165 29236
rect -69485 29864 -69165 29890
rect -69485 29236 -69479 29864
rect -69171 29236 -69165 29864
rect -69485 29210 -69165 29236
rect -68485 29864 -68165 29890
rect -68485 29236 -68479 29864
rect -68171 29236 -68165 29864
rect -68485 29210 -68165 29236
rect -67485 29864 -67165 29890
rect -67485 29236 -67479 29864
rect -67171 29236 -67165 29864
rect -67485 29210 -67165 29236
rect -66485 29864 -66165 29890
rect -66485 29236 -66479 29864
rect -66171 29236 -66165 29864
rect -66485 29210 -66165 29236
rect -65485 29864 -65165 29890
rect -65485 29236 -65479 29864
rect -65171 29236 -65165 29864
rect -65485 29210 -65165 29236
rect -64485 29864 -64165 29890
rect -64485 29236 -64479 29864
rect -64171 29236 -64165 29864
rect -64485 29210 -64165 29236
rect -63485 29864 -63165 29890
rect -63485 29236 -63479 29864
rect -63171 29236 -63165 29864
rect -63485 29210 -63165 29236
rect -62485 29864 -62165 29890
rect -62485 29236 -62479 29864
rect -62171 29236 -62165 29864
rect -62485 29210 -62165 29236
rect -61485 29864 -61165 29890
rect -61485 29236 -61479 29864
rect -61171 29236 -61165 29864
rect -61485 29210 -61165 29236
rect -60485 29864 -60165 29890
rect -60485 29236 -60479 29864
rect -60171 29236 -60165 29864
rect -60485 29210 -60165 29236
rect -59485 29864 -59165 29890
rect -59485 29236 -59479 29864
rect -59171 29236 -59165 29864
rect -59485 29210 -59165 29236
rect -74825 29204 -58825 29210
rect -74825 28896 -74819 29204
rect -74511 29198 -74139 29204
rect -73511 29198 -73139 29204
rect -72511 29198 -72139 29204
rect -71511 29198 -71139 29204
rect -70511 29198 -70139 29204
rect -69511 29198 -69139 29204
rect -68511 29198 -68139 29204
rect -67511 29198 -67139 29204
rect -66511 29198 -66139 29204
rect -65511 29198 -65139 29204
rect -64511 29198 -64139 29204
rect -63511 29198 -63139 29204
rect -62511 29198 -62139 29204
rect -61511 29198 -61139 29204
rect -60511 29198 -60139 29204
rect -59511 29198 -59139 29204
rect -74511 28902 -74473 29198
rect -74177 28902 -74139 29198
rect -73511 28902 -73473 29198
rect -73177 28902 -73139 29198
rect -72511 28902 -72473 29198
rect -72177 28902 -72139 29198
rect -71511 28902 -71473 29198
rect -71177 28902 -71139 29198
rect -70511 28902 -70473 29198
rect -70177 28902 -70139 29198
rect -69511 28902 -69473 29198
rect -69177 28902 -69139 29198
rect -68511 28902 -68473 29198
rect -68177 28902 -68139 29198
rect -67511 28902 -67473 29198
rect -67177 28902 -67139 29198
rect -66511 28902 -66473 29198
rect -66177 28902 -66139 29198
rect -65511 28902 -65473 29198
rect -65177 28902 -65139 29198
rect -64511 28902 -64473 29198
rect -64177 28902 -64139 29198
rect -63511 28902 -63473 29198
rect -63177 28902 -63139 29198
rect -62511 28902 -62473 29198
rect -62177 28902 -62139 29198
rect -61511 28902 -61473 29198
rect -61177 28902 -61139 29198
rect -60511 28902 -60473 29198
rect -60177 28902 -60139 29198
rect -59511 28902 -59473 29198
rect -59177 28902 -59139 29198
rect -74511 28896 -74139 28902
rect -73511 28896 -73139 28902
rect -72511 28896 -72139 28902
rect -71511 28896 -71139 28902
rect -70511 28896 -70139 28902
rect -69511 28896 -69139 28902
rect -68511 28896 -68139 28902
rect -67511 28896 -67139 28902
rect -66511 28896 -66139 28902
rect -65511 28896 -65139 28902
rect -64511 28896 -64139 28902
rect -63511 28896 -63139 28902
rect -62511 28896 -62139 28902
rect -61511 28896 -61139 28902
rect -60511 28896 -60139 28902
rect -59511 28896 -59139 28902
rect -58831 28896 -58825 29204
rect -74825 28890 -58825 28896
rect -74485 28864 -74165 28890
rect -74485 28556 -74479 28864
rect -74171 28556 -74165 28864
rect -74485 28550 -74165 28556
rect -73485 28864 -73165 28890
rect -73485 28556 -73479 28864
rect -73171 28556 -73165 28864
rect -73485 28550 -73165 28556
rect -72485 28864 -72165 28890
rect -72485 28556 -72479 28864
rect -72171 28556 -72165 28864
rect -72485 28550 -72165 28556
rect -71485 28864 -71165 28890
rect -71485 28556 -71479 28864
rect -71171 28556 -71165 28864
rect -71485 28550 -71165 28556
rect -70485 28864 -70165 28890
rect -70485 28556 -70479 28864
rect -70171 28556 -70165 28864
rect -70485 28550 -70165 28556
rect -69485 28864 -69165 28890
rect -69485 28556 -69479 28864
rect -69171 28556 -69165 28864
rect -69485 28550 -69165 28556
rect -68485 28864 -68165 28890
rect -68485 28556 -68479 28864
rect -68171 28556 -68165 28864
rect -68485 28550 -68165 28556
rect -67485 28864 -67165 28890
rect -67485 28556 -67479 28864
rect -67171 28556 -67165 28864
rect -67485 28550 -67165 28556
rect -66485 28864 -66165 28890
rect -66485 28556 -66479 28864
rect -66171 28556 -66165 28864
rect -66485 28550 -66165 28556
rect -65485 28864 -65165 28890
rect -65485 28556 -65479 28864
rect -65171 28556 -65165 28864
rect -65485 28550 -65165 28556
rect -64485 28864 -64165 28890
rect -64485 28556 -64479 28864
rect -64171 28556 -64165 28864
rect -64485 28550 -64165 28556
rect -63485 28864 -63165 28890
rect -63485 28556 -63479 28864
rect -63171 28556 -63165 28864
rect -63485 28550 -63165 28556
rect -62485 28864 -62165 28890
rect -62485 28556 -62479 28864
rect -62171 28556 -62165 28864
rect -62485 28550 -62165 28556
rect -61485 28864 -61165 28890
rect -61485 28556 -61479 28864
rect -61171 28556 -61165 28864
rect -61485 28550 -61165 28556
rect -60485 28864 -60165 28890
rect -60485 28556 -60479 28864
rect -60171 28556 -60165 28864
rect -60485 28550 -60165 28556
rect -59485 28864 -59165 28890
rect -59485 28556 -59479 28864
rect -59171 28556 -59165 28864
rect -59485 28550 -59165 28556
rect -47625 26087 -47025 32584
rect 3043 32581 4917 32593
rect 3043 32529 3049 32581
rect 3101 32529 3365 32581
rect 3417 32529 3681 32581
rect 3733 32529 3997 32581
rect 4049 32529 4313 32581
rect 4365 32529 4917 32581
rect 3043 32517 4917 32529
rect 3043 32465 3049 32517
rect 3101 32465 3365 32517
rect 3417 32465 3681 32517
rect 3733 32465 3997 32517
rect 4049 32465 4313 32517
rect 4365 32465 4917 32517
rect 3043 32459 4917 32465
rect -72825 25949 -60825 26000
rect -72825 25943 -72776 25949
rect -60884 25943 -60825 25949
rect -72825 16047 -72778 25943
rect -60882 16047 -60825 25943
rect -47625 25523 -47607 26087
rect -47043 25523 -47025 26087
rect 6620 26131 7220 32704
rect 9994 32864 10314 32890
rect 9994 32236 10000 32864
rect 10308 32236 10314 32864
rect 9994 32210 10314 32236
rect 10994 32864 11314 32890
rect 10994 32236 11000 32864
rect 11308 32236 11314 32864
rect 10994 32210 11314 32236
rect 11994 32864 12314 32890
rect 11994 32236 12000 32864
rect 12308 32236 12314 32864
rect 11994 32210 12314 32236
rect 12994 32864 13314 32890
rect 12994 32236 13000 32864
rect 13308 32236 13314 32864
rect 12994 32210 13314 32236
rect 13994 32864 14314 32890
rect 13994 32236 14000 32864
rect 14308 32236 14314 32864
rect 13994 32210 14314 32236
rect 14994 32864 15314 32890
rect 14994 32236 15000 32864
rect 15308 32236 15314 32864
rect 14994 32210 15314 32236
rect 15994 32864 16314 32890
rect 15994 32236 16000 32864
rect 16308 32236 16314 32864
rect 15994 32210 16314 32236
rect 16994 32864 17314 32890
rect 16994 32236 17000 32864
rect 17308 32236 17314 32864
rect 16994 32210 17314 32236
rect 17994 32864 18314 32890
rect 17994 32236 18000 32864
rect 18308 32236 18314 32864
rect 17994 32210 18314 32236
rect 18994 32864 19314 32890
rect 18994 32236 19000 32864
rect 19308 32236 19314 32864
rect 18994 32210 19314 32236
rect 19994 32864 20314 32890
rect 19994 32236 20000 32864
rect 20308 32236 20314 32864
rect 19994 32210 20314 32236
rect 20994 32864 21314 32890
rect 20994 32236 21000 32864
rect 21308 32236 21314 32864
rect 20994 32210 21314 32236
rect 21994 32864 22314 32890
rect 21994 32236 22000 32864
rect 22308 32236 22314 32864
rect 21994 32210 22314 32236
rect 22994 32864 23314 32890
rect 22994 32236 23000 32864
rect 23308 32236 23314 32864
rect 22994 32210 23314 32236
rect 23994 32864 24314 32890
rect 23994 32236 24000 32864
rect 24308 32236 24314 32864
rect 23994 32210 24314 32236
rect 24994 32864 25314 32890
rect 24994 32236 25000 32864
rect 25308 32236 25314 32864
rect 24994 32210 25314 32236
rect 25994 32864 26314 32890
rect 25994 32236 26000 32864
rect 26308 32236 26314 32864
rect 25994 32210 26314 32236
rect 26994 32864 27314 32890
rect 26994 32236 27000 32864
rect 27308 32236 27314 32864
rect 26994 32210 27314 32236
rect 27994 32864 28314 32890
rect 27994 32236 28000 32864
rect 28308 32236 28314 32864
rect 27994 32210 28314 32236
rect 28994 32864 29314 32890
rect 28994 32236 29000 32864
rect 29308 32236 29314 32864
rect 28994 32210 29314 32236
rect 29994 32864 30314 32890
rect 29994 32236 30000 32864
rect 30308 32236 30314 32864
rect 29994 32210 30314 32236
rect 30994 32864 31314 32890
rect 30994 32236 31000 32864
rect 31308 32236 31314 32864
rect 30994 32210 31314 32236
rect 31994 32864 32314 32890
rect 31994 32236 32000 32864
rect 32308 32236 32314 32864
rect 31994 32210 32314 32236
rect 32994 32864 33314 32890
rect 32994 32236 33000 32864
rect 33308 32236 33314 32864
rect 32994 32210 33314 32236
rect 33994 32864 34314 32890
rect 33994 32236 34000 32864
rect 34308 32236 34314 32864
rect 33994 32210 34314 32236
rect 9654 32204 34654 32210
rect 9654 31896 9660 32204
rect 9968 32198 10340 32204
rect 10968 32198 11340 32204
rect 11968 32198 12340 32204
rect 12968 32198 13340 32204
rect 13968 32198 14340 32204
rect 14968 32198 15340 32204
rect 15968 32198 16340 32204
rect 16968 32198 17340 32204
rect 17968 32198 18340 32204
rect 18968 32198 19340 32204
rect 19968 32198 20340 32204
rect 20968 32198 21340 32204
rect 21968 32198 22340 32204
rect 22968 32198 23340 32204
rect 23968 32198 24340 32204
rect 24968 32198 25340 32204
rect 25968 32198 26340 32204
rect 26968 32198 27340 32204
rect 27968 32198 28340 32204
rect 28968 32198 29340 32204
rect 29968 32198 30340 32204
rect 30968 32198 31340 32204
rect 31968 32198 32340 32204
rect 32968 32198 33340 32204
rect 33968 32198 34340 32204
rect 9968 31902 10006 32198
rect 10302 31902 10340 32198
rect 10968 31902 11006 32198
rect 11302 31902 11340 32198
rect 11968 31902 12006 32198
rect 12302 31902 12340 32198
rect 12968 31902 13006 32198
rect 13302 31902 13340 32198
rect 13968 31902 14006 32198
rect 14302 31902 14340 32198
rect 14968 31902 15006 32198
rect 15302 31902 15340 32198
rect 15968 31902 16006 32198
rect 16302 31902 16340 32198
rect 16968 31902 17006 32198
rect 17302 31902 17340 32198
rect 17968 31902 18006 32198
rect 18302 31902 18340 32198
rect 18968 31902 19006 32198
rect 19302 31902 19340 32198
rect 19968 31902 20006 32198
rect 20302 31902 20340 32198
rect 20968 31902 21006 32198
rect 21302 31902 21340 32198
rect 21968 31902 22006 32198
rect 22302 31902 22340 32198
rect 22968 31902 23006 32198
rect 23302 31902 23340 32198
rect 23968 31902 24006 32198
rect 24302 31902 24340 32198
rect 24968 31902 25006 32198
rect 25302 31902 25340 32198
rect 25968 31902 26006 32198
rect 26302 31902 26340 32198
rect 26968 31902 27006 32198
rect 27302 31902 27340 32198
rect 27968 31902 28006 32198
rect 28302 31902 28340 32198
rect 28968 31902 29006 32198
rect 29302 31902 29340 32198
rect 29968 31902 30006 32198
rect 30302 31902 30340 32198
rect 30968 31902 31006 32198
rect 31302 31902 31340 32198
rect 31968 31902 32006 32198
rect 32302 31902 32340 32198
rect 32968 31902 33006 32198
rect 33302 31902 33340 32198
rect 33968 31902 34006 32198
rect 34302 31902 34340 32198
rect 9968 31896 10340 31902
rect 10968 31896 11340 31902
rect 11968 31896 12340 31902
rect 12968 31896 13340 31902
rect 13968 31896 14340 31902
rect 14968 31896 15340 31902
rect 15968 31896 16340 31902
rect 16968 31896 17340 31902
rect 17968 31896 18340 31902
rect 18968 31896 19340 31902
rect 19968 31896 20340 31902
rect 20968 31896 21340 31902
rect 21968 31896 22340 31902
rect 22968 31896 23340 31902
rect 23968 31896 24340 31902
rect 24968 31896 25340 31902
rect 25968 31896 26340 31902
rect 26968 31896 27340 31902
rect 27968 31896 28340 31902
rect 28968 31896 29340 31902
rect 29968 31896 30340 31902
rect 30968 31896 31340 31902
rect 31968 31896 32340 31902
rect 32968 31896 33340 31902
rect 33968 31896 34340 31902
rect 34648 31896 34654 32204
rect 9654 31890 34654 31896
rect 9994 31864 10314 31890
rect 9994 31236 10000 31864
rect 10308 31236 10314 31864
rect 9994 31210 10314 31236
rect 10994 31864 11314 31890
rect 10994 31236 11000 31864
rect 11308 31236 11314 31864
rect 10994 31210 11314 31236
rect 11994 31864 12314 31890
rect 11994 31236 12000 31864
rect 12308 31236 12314 31864
rect 11994 31210 12314 31236
rect 12994 31864 13314 31890
rect 12994 31236 13000 31864
rect 13308 31236 13314 31864
rect 12994 31210 13314 31236
rect 13994 31864 14314 31890
rect 13994 31236 14000 31864
rect 14308 31236 14314 31864
rect 13994 31210 14314 31236
rect 14994 31864 15314 31890
rect 14994 31236 15000 31864
rect 15308 31236 15314 31864
rect 14994 31210 15314 31236
rect 15994 31864 16314 31890
rect 15994 31236 16000 31864
rect 16308 31236 16314 31864
rect 15994 31210 16314 31236
rect 16994 31864 17314 31890
rect 16994 31236 17000 31864
rect 17308 31236 17314 31864
rect 16994 31210 17314 31236
rect 17994 31864 18314 31890
rect 17994 31236 18000 31864
rect 18308 31236 18314 31864
rect 17994 31210 18314 31236
rect 18994 31864 19314 31890
rect 18994 31236 19000 31864
rect 19308 31236 19314 31864
rect 18994 31210 19314 31236
rect 19994 31864 20314 31890
rect 19994 31236 20000 31864
rect 20308 31236 20314 31864
rect 19994 31210 20314 31236
rect 20994 31864 21314 31890
rect 20994 31236 21000 31864
rect 21308 31236 21314 31864
rect 20994 31210 21314 31236
rect 21994 31864 22314 31890
rect 21994 31236 22000 31864
rect 22308 31236 22314 31864
rect 21994 31210 22314 31236
rect 22994 31864 23314 31890
rect 22994 31236 23000 31864
rect 23308 31236 23314 31864
rect 22994 31210 23314 31236
rect 23994 31864 24314 31890
rect 23994 31236 24000 31864
rect 24308 31236 24314 31864
rect 23994 31210 24314 31236
rect 24994 31864 25314 31890
rect 24994 31236 25000 31864
rect 25308 31236 25314 31864
rect 24994 31210 25314 31236
rect 25994 31864 26314 31890
rect 25994 31236 26000 31864
rect 26308 31236 26314 31864
rect 25994 31210 26314 31236
rect 26994 31864 27314 31890
rect 26994 31236 27000 31864
rect 27308 31236 27314 31864
rect 26994 31210 27314 31236
rect 27994 31864 28314 31890
rect 27994 31236 28000 31864
rect 28308 31236 28314 31864
rect 27994 31210 28314 31236
rect 28994 31864 29314 31890
rect 28994 31236 29000 31864
rect 29308 31236 29314 31864
rect 28994 31210 29314 31236
rect 29994 31864 30314 31890
rect 29994 31236 30000 31864
rect 30308 31236 30314 31864
rect 29994 31210 30314 31236
rect 30994 31864 31314 31890
rect 30994 31236 31000 31864
rect 31308 31236 31314 31864
rect 30994 31210 31314 31236
rect 31994 31864 32314 31890
rect 31994 31236 32000 31864
rect 32308 31236 32314 31864
rect 31994 31210 32314 31236
rect 32994 31864 33314 31890
rect 32994 31236 33000 31864
rect 33308 31236 33314 31864
rect 32994 31210 33314 31236
rect 33994 31864 34314 31890
rect 33994 31236 34000 31864
rect 34308 31236 34314 31864
rect 33994 31210 34314 31236
rect 9654 31204 34654 31210
rect 9654 30896 9660 31204
rect 9968 31198 10340 31204
rect 10968 31198 11340 31204
rect 11968 31198 12340 31204
rect 12968 31198 13340 31204
rect 13968 31198 14340 31204
rect 14968 31198 15340 31204
rect 15968 31198 16340 31204
rect 16968 31198 17340 31204
rect 17968 31198 18340 31204
rect 18968 31198 19340 31204
rect 19968 31198 20340 31204
rect 20968 31198 21340 31204
rect 21968 31198 22340 31204
rect 22968 31198 23340 31204
rect 23968 31198 24340 31204
rect 24968 31198 25340 31204
rect 25968 31198 26340 31204
rect 26968 31198 27340 31204
rect 27968 31198 28340 31204
rect 28968 31198 29340 31204
rect 29968 31198 30340 31204
rect 30968 31198 31340 31204
rect 31968 31198 32340 31204
rect 32968 31198 33340 31204
rect 33968 31198 34340 31204
rect 9968 30902 10006 31198
rect 10302 30902 10340 31198
rect 10968 30902 11006 31198
rect 11302 30902 11340 31198
rect 11968 30902 12006 31198
rect 12302 30902 12340 31198
rect 12968 30902 13006 31198
rect 13302 30902 13340 31198
rect 13968 30902 14006 31198
rect 14302 30902 14340 31198
rect 14968 30902 15006 31198
rect 15302 30902 15340 31198
rect 15968 30902 16006 31198
rect 16302 30902 16340 31198
rect 16968 30902 17006 31198
rect 17302 30902 17340 31198
rect 17968 30902 18006 31198
rect 18302 30902 18340 31198
rect 18968 30902 19006 31198
rect 19302 30902 19340 31198
rect 19968 30902 20006 31198
rect 20302 30902 20340 31198
rect 20968 30902 21006 31198
rect 21302 30902 21340 31198
rect 21968 30902 22006 31198
rect 22302 30902 22340 31198
rect 22968 30902 23006 31198
rect 23302 30902 23340 31198
rect 23968 30902 24006 31198
rect 24302 30902 24340 31198
rect 24968 30902 25006 31198
rect 25302 30902 25340 31198
rect 25968 30902 26006 31198
rect 26302 30902 26340 31198
rect 26968 30902 27006 31198
rect 27302 30902 27340 31198
rect 27968 30902 28006 31198
rect 28302 30902 28340 31198
rect 28968 30902 29006 31198
rect 29302 30902 29340 31198
rect 29968 30902 30006 31198
rect 30302 30902 30340 31198
rect 30968 30902 31006 31198
rect 31302 30902 31340 31198
rect 31968 30902 32006 31198
rect 32302 30902 32340 31198
rect 32968 30902 33006 31198
rect 33302 30902 33340 31198
rect 33968 30902 34006 31198
rect 34302 30902 34340 31198
rect 9968 30896 10340 30902
rect 10968 30896 11340 30902
rect 11968 30896 12340 30902
rect 12968 30896 13340 30902
rect 13968 30896 14340 30902
rect 14968 30896 15340 30902
rect 15968 30896 16340 30902
rect 16968 30896 17340 30902
rect 17968 30896 18340 30902
rect 18968 30896 19340 30902
rect 19968 30896 20340 30902
rect 20968 30896 21340 30902
rect 21968 30896 22340 30902
rect 22968 30896 23340 30902
rect 23968 30896 24340 30902
rect 24968 30896 25340 30902
rect 25968 30896 26340 30902
rect 26968 30896 27340 30902
rect 27968 30896 28340 30902
rect 28968 30896 29340 30902
rect 29968 30896 30340 30902
rect 30968 30896 31340 30902
rect 31968 30896 32340 30902
rect 32968 30896 33340 30902
rect 33968 30896 34340 30902
rect 34648 30896 34654 31204
rect 9654 30890 34654 30896
rect 9994 30864 10314 30890
rect 9994 30236 10000 30864
rect 10308 30236 10314 30864
rect 9994 30210 10314 30236
rect 10994 30864 11314 30890
rect 10994 30236 11000 30864
rect 11308 30236 11314 30864
rect 10994 30210 11314 30236
rect 11994 30864 12314 30890
rect 11994 30236 12000 30864
rect 12308 30236 12314 30864
rect 11994 30210 12314 30236
rect 12994 30864 13314 30890
rect 12994 30236 13000 30864
rect 13308 30236 13314 30864
rect 12994 30210 13314 30236
rect 13994 30864 14314 30890
rect 13994 30236 14000 30864
rect 14308 30236 14314 30864
rect 13994 30210 14314 30236
rect 14994 30864 15314 30890
rect 14994 30236 15000 30864
rect 15308 30236 15314 30864
rect 14994 30210 15314 30236
rect 15994 30864 16314 30890
rect 15994 30236 16000 30864
rect 16308 30236 16314 30864
rect 15994 30210 16314 30236
rect 16994 30864 17314 30890
rect 16994 30236 17000 30864
rect 17308 30236 17314 30864
rect 16994 30210 17314 30236
rect 17994 30864 18314 30890
rect 17994 30236 18000 30864
rect 18308 30236 18314 30864
rect 17994 30210 18314 30236
rect 18994 30864 19314 30890
rect 18994 30236 19000 30864
rect 19308 30236 19314 30864
rect 18994 30210 19314 30236
rect 19994 30864 20314 30890
rect 19994 30236 20000 30864
rect 20308 30236 20314 30864
rect 19994 30210 20314 30236
rect 20994 30864 21314 30890
rect 20994 30236 21000 30864
rect 21308 30236 21314 30864
rect 20994 30210 21314 30236
rect 21994 30864 22314 30890
rect 21994 30236 22000 30864
rect 22308 30236 22314 30864
rect 21994 30210 22314 30236
rect 22994 30864 23314 30890
rect 22994 30236 23000 30864
rect 23308 30236 23314 30864
rect 22994 30210 23314 30236
rect 23994 30864 24314 30890
rect 23994 30236 24000 30864
rect 24308 30236 24314 30864
rect 23994 30210 24314 30236
rect 24994 30864 25314 30890
rect 24994 30236 25000 30864
rect 25308 30236 25314 30864
rect 24994 30210 25314 30236
rect 25994 30864 26314 30890
rect 25994 30236 26000 30864
rect 26308 30236 26314 30864
rect 25994 30210 26314 30236
rect 26994 30864 27314 30890
rect 26994 30236 27000 30864
rect 27308 30236 27314 30864
rect 26994 30210 27314 30236
rect 27994 30864 28314 30890
rect 27994 30236 28000 30864
rect 28308 30236 28314 30864
rect 27994 30210 28314 30236
rect 28994 30864 29314 30890
rect 28994 30236 29000 30864
rect 29308 30236 29314 30864
rect 28994 30210 29314 30236
rect 29994 30864 30314 30890
rect 29994 30236 30000 30864
rect 30308 30236 30314 30864
rect 29994 30210 30314 30236
rect 30994 30864 31314 30890
rect 30994 30236 31000 30864
rect 31308 30236 31314 30864
rect 30994 30210 31314 30236
rect 31994 30864 32314 30890
rect 31994 30236 32000 30864
rect 32308 30236 32314 30864
rect 31994 30210 32314 30236
rect 32994 30864 33314 30890
rect 32994 30236 33000 30864
rect 33308 30236 33314 30864
rect 32994 30210 33314 30236
rect 33994 30864 34314 30890
rect 33994 30236 34000 30864
rect 34308 30236 34314 30864
rect 33994 30210 34314 30236
rect 9654 30204 34654 30210
rect 9654 29896 9660 30204
rect 9968 30198 10340 30204
rect 10968 30198 11340 30204
rect 11968 30198 12340 30204
rect 12968 30198 13340 30204
rect 13968 30198 14340 30204
rect 14968 30198 15340 30204
rect 15968 30198 16340 30204
rect 16968 30198 17340 30204
rect 17968 30198 18340 30204
rect 18968 30198 19340 30204
rect 19968 30198 20340 30204
rect 20968 30198 21340 30204
rect 21968 30198 22340 30204
rect 22968 30198 23340 30204
rect 23968 30198 24340 30204
rect 24968 30198 25340 30204
rect 25968 30198 26340 30204
rect 26968 30198 27340 30204
rect 27968 30198 28340 30204
rect 28968 30198 29340 30204
rect 29968 30198 30340 30204
rect 30968 30198 31340 30204
rect 31968 30198 32340 30204
rect 32968 30198 33340 30204
rect 33968 30198 34340 30204
rect 9968 29902 10006 30198
rect 10302 29902 10340 30198
rect 10968 29902 11006 30198
rect 11302 29902 11340 30198
rect 11968 29902 12006 30198
rect 12302 29902 12340 30198
rect 12968 29902 13006 30198
rect 13302 29902 13340 30198
rect 13968 29902 14006 30198
rect 14302 29902 14340 30198
rect 14968 29902 15006 30198
rect 15302 29902 15340 30198
rect 15968 29902 16006 30198
rect 16302 29902 16340 30198
rect 16968 29902 17006 30198
rect 17302 29902 17340 30198
rect 17968 29902 18006 30198
rect 18302 29902 18340 30198
rect 18968 29902 19006 30198
rect 19302 29902 19340 30198
rect 19968 29902 20006 30198
rect 20302 29902 20340 30198
rect 20968 29902 21006 30198
rect 21302 29902 21340 30198
rect 21968 29902 22006 30198
rect 22302 29902 22340 30198
rect 22968 29902 23006 30198
rect 23302 29902 23340 30198
rect 23968 29902 24006 30198
rect 24302 29902 24340 30198
rect 24968 29902 25006 30198
rect 25302 29902 25340 30198
rect 25968 29902 26006 30198
rect 26302 29902 26340 30198
rect 26968 29902 27006 30198
rect 27302 29902 27340 30198
rect 27968 29902 28006 30198
rect 28302 29902 28340 30198
rect 28968 29902 29006 30198
rect 29302 29902 29340 30198
rect 29968 29902 30006 30198
rect 30302 29902 30340 30198
rect 30968 29902 31006 30198
rect 31302 29902 31340 30198
rect 31968 29902 32006 30198
rect 32302 29902 32340 30198
rect 32968 29902 33006 30198
rect 33302 29902 33340 30198
rect 33968 29902 34006 30198
rect 34302 29902 34340 30198
rect 9968 29896 10340 29902
rect 10968 29896 11340 29902
rect 11968 29896 12340 29902
rect 12968 29896 13340 29902
rect 13968 29896 14340 29902
rect 14968 29896 15340 29902
rect 15968 29896 16340 29902
rect 16968 29896 17340 29902
rect 17968 29896 18340 29902
rect 18968 29896 19340 29902
rect 19968 29896 20340 29902
rect 20968 29896 21340 29902
rect 21968 29896 22340 29902
rect 22968 29896 23340 29902
rect 23968 29896 24340 29902
rect 24968 29896 25340 29902
rect 25968 29896 26340 29902
rect 26968 29896 27340 29902
rect 27968 29896 28340 29902
rect 28968 29896 29340 29902
rect 29968 29896 30340 29902
rect 30968 29896 31340 29902
rect 31968 29896 32340 29902
rect 32968 29896 33340 29902
rect 33968 29896 34340 29902
rect 34648 29896 34654 30204
rect 9654 29890 34654 29896
rect 9994 29864 10314 29890
rect 9994 29236 10000 29864
rect 10308 29236 10314 29864
rect 9994 29210 10314 29236
rect 10994 29864 11314 29890
rect 10994 29236 11000 29864
rect 11308 29236 11314 29864
rect 10994 29210 11314 29236
rect 11994 29864 12314 29890
rect 11994 29236 12000 29864
rect 12308 29236 12314 29864
rect 11994 29210 12314 29236
rect 12994 29864 13314 29890
rect 12994 29236 13000 29864
rect 13308 29236 13314 29864
rect 12994 29210 13314 29236
rect 13994 29864 14314 29890
rect 13994 29236 14000 29864
rect 14308 29236 14314 29864
rect 13994 29210 14314 29236
rect 14994 29864 15314 29890
rect 14994 29236 15000 29864
rect 15308 29236 15314 29864
rect 14994 29210 15314 29236
rect 15994 29864 16314 29890
rect 15994 29236 16000 29864
rect 16308 29236 16314 29864
rect 15994 29210 16314 29236
rect 16994 29864 17314 29890
rect 16994 29236 17000 29864
rect 17308 29236 17314 29864
rect 16994 29210 17314 29236
rect 17994 29864 18314 29890
rect 17994 29236 18000 29864
rect 18308 29236 18314 29864
rect 17994 29210 18314 29236
rect 18994 29864 19314 29890
rect 18994 29236 19000 29864
rect 19308 29236 19314 29864
rect 18994 29210 19314 29236
rect 19994 29864 20314 29890
rect 19994 29236 20000 29864
rect 20308 29236 20314 29864
rect 19994 29210 20314 29236
rect 20994 29864 21314 29890
rect 20994 29236 21000 29864
rect 21308 29236 21314 29864
rect 20994 29210 21314 29236
rect 21994 29864 22314 29890
rect 21994 29236 22000 29864
rect 22308 29236 22314 29864
rect 21994 29210 22314 29236
rect 22994 29864 23314 29890
rect 22994 29236 23000 29864
rect 23308 29236 23314 29864
rect 22994 29210 23314 29236
rect 23994 29864 24314 29890
rect 23994 29236 24000 29864
rect 24308 29236 24314 29864
rect 23994 29210 24314 29236
rect 24994 29864 25314 29890
rect 24994 29236 25000 29864
rect 25308 29236 25314 29864
rect 24994 29210 25314 29236
rect 25994 29864 26314 29890
rect 25994 29236 26000 29864
rect 26308 29236 26314 29864
rect 25994 29210 26314 29236
rect 26994 29864 27314 29890
rect 26994 29236 27000 29864
rect 27308 29236 27314 29864
rect 26994 29210 27314 29236
rect 27994 29864 28314 29890
rect 27994 29236 28000 29864
rect 28308 29236 28314 29864
rect 27994 29210 28314 29236
rect 28994 29864 29314 29890
rect 28994 29236 29000 29864
rect 29308 29236 29314 29864
rect 28994 29210 29314 29236
rect 29994 29864 30314 29890
rect 29994 29236 30000 29864
rect 30308 29236 30314 29864
rect 29994 29210 30314 29236
rect 30994 29864 31314 29890
rect 30994 29236 31000 29864
rect 31308 29236 31314 29864
rect 30994 29210 31314 29236
rect 31994 29864 32314 29890
rect 31994 29236 32000 29864
rect 32308 29236 32314 29864
rect 31994 29210 32314 29236
rect 32994 29864 33314 29890
rect 32994 29236 33000 29864
rect 33308 29236 33314 29864
rect 32994 29210 33314 29236
rect 33994 29864 34314 29890
rect 33994 29236 34000 29864
rect 34308 29236 34314 29864
rect 33994 29210 34314 29236
rect 9654 29204 34654 29210
rect 9654 28896 9660 29204
rect 9968 29198 10340 29204
rect 10968 29198 11340 29204
rect 11968 29198 12340 29204
rect 12968 29198 13340 29204
rect 13968 29198 14340 29204
rect 14968 29198 15340 29204
rect 15968 29198 16340 29204
rect 16968 29198 17340 29204
rect 17968 29198 18340 29204
rect 18968 29198 19340 29204
rect 19968 29198 20340 29204
rect 20968 29198 21340 29204
rect 21968 29198 22340 29204
rect 22968 29198 23340 29204
rect 23968 29198 24340 29204
rect 24968 29198 25340 29204
rect 25968 29198 26340 29204
rect 26968 29198 27340 29204
rect 27968 29198 28340 29204
rect 28968 29198 29340 29204
rect 29968 29198 30340 29204
rect 30968 29198 31340 29204
rect 31968 29198 32340 29204
rect 32968 29198 33340 29204
rect 33968 29198 34340 29204
rect 9968 28902 10006 29198
rect 10302 28902 10340 29198
rect 10968 28902 11006 29198
rect 11302 28902 11340 29198
rect 11968 28902 12006 29198
rect 12302 28902 12340 29198
rect 12968 28902 13006 29198
rect 13302 28902 13340 29198
rect 13968 28902 14006 29198
rect 14302 28902 14340 29198
rect 14968 28902 15006 29198
rect 15302 28902 15340 29198
rect 15968 28902 16006 29198
rect 16302 28902 16340 29198
rect 16968 28902 17006 29198
rect 17302 28902 17340 29198
rect 17968 28902 18006 29198
rect 18302 28902 18340 29198
rect 18968 28902 19006 29198
rect 19302 28902 19340 29198
rect 19968 28902 20006 29198
rect 20302 28902 20340 29198
rect 20968 28902 21006 29198
rect 21302 28902 21340 29198
rect 21968 28902 22006 29198
rect 22302 28902 22340 29198
rect 22968 28902 23006 29198
rect 23302 28902 23340 29198
rect 23968 28902 24006 29198
rect 24302 28902 24340 29198
rect 24968 28902 25006 29198
rect 25302 28902 25340 29198
rect 25968 28902 26006 29198
rect 26302 28902 26340 29198
rect 26968 28902 27006 29198
rect 27302 28902 27340 29198
rect 27968 28902 28006 29198
rect 28302 28902 28340 29198
rect 28968 28902 29006 29198
rect 29302 28902 29340 29198
rect 29968 28902 30006 29198
rect 30302 28902 30340 29198
rect 30968 28902 31006 29198
rect 31302 28902 31340 29198
rect 31968 28902 32006 29198
rect 32302 28902 32340 29198
rect 32968 28902 33006 29198
rect 33302 28902 33340 29198
rect 33968 28902 34006 29198
rect 34302 28902 34340 29198
rect 9968 28896 10340 28902
rect 10968 28896 11340 28902
rect 11968 28896 12340 28902
rect 12968 28896 13340 28902
rect 13968 28896 14340 28902
rect 14968 28896 15340 28902
rect 15968 28896 16340 28902
rect 16968 28896 17340 28902
rect 17968 28896 18340 28902
rect 18968 28896 19340 28902
rect 19968 28896 20340 28902
rect 20968 28896 21340 28902
rect 21968 28896 22340 28902
rect 22968 28896 23340 28902
rect 23968 28896 24340 28902
rect 24968 28896 25340 28902
rect 25968 28896 26340 28902
rect 26968 28896 27340 28902
rect 27968 28896 28340 28902
rect 28968 28896 29340 28902
rect 29968 28896 30340 28902
rect 30968 28896 31340 28902
rect 31968 28896 32340 28902
rect 32968 28896 33340 28902
rect 33968 28896 34340 28902
rect 34648 28896 34654 29204
rect 9654 28890 34654 28896
rect 9994 28864 10314 28890
rect 9994 28556 10000 28864
rect 10308 28556 10314 28864
rect 9994 28550 10314 28556
rect 10994 28864 11314 28890
rect 10994 28556 11000 28864
rect 11308 28556 11314 28864
rect 10994 28550 11314 28556
rect 11994 28864 12314 28890
rect 11994 28556 12000 28864
rect 12308 28556 12314 28864
rect 11994 28550 12314 28556
rect 12994 28864 13314 28890
rect 12994 28556 13000 28864
rect 13308 28556 13314 28864
rect 12994 28550 13314 28556
rect 13994 28864 14314 28890
rect 13994 28556 14000 28864
rect 14308 28556 14314 28864
rect 13994 28550 14314 28556
rect 14994 28864 15314 28890
rect 14994 28556 15000 28864
rect 15308 28556 15314 28864
rect 14994 28550 15314 28556
rect 15994 28864 16314 28890
rect 15994 28556 16000 28864
rect 16308 28556 16314 28864
rect 15994 28550 16314 28556
rect 16994 28864 17314 28890
rect 16994 28556 17000 28864
rect 17308 28556 17314 28864
rect 16994 28550 17314 28556
rect 17994 28864 18314 28890
rect 17994 28556 18000 28864
rect 18308 28556 18314 28864
rect 17994 28550 18314 28556
rect 18994 28864 19314 28890
rect 18994 28556 19000 28864
rect 19308 28556 19314 28864
rect 18994 28550 19314 28556
rect 19994 28864 20314 28890
rect 19994 28556 20000 28864
rect 20308 28556 20314 28864
rect 19994 28550 20314 28556
rect 20994 28864 21314 28890
rect 20994 28556 21000 28864
rect 21308 28556 21314 28864
rect 20994 28550 21314 28556
rect 21994 28864 22314 28890
rect 21994 28556 22000 28864
rect 22308 28556 22314 28864
rect 21994 28550 22314 28556
rect 22994 28864 23314 28890
rect 22994 28556 23000 28864
rect 23308 28556 23314 28864
rect 22994 28550 23314 28556
rect 23994 28864 24314 28890
rect 23994 28556 24000 28864
rect 24308 28556 24314 28864
rect 23994 28550 24314 28556
rect 24994 28864 25314 28890
rect 24994 28556 25000 28864
rect 25308 28556 25314 28864
rect 24994 28550 25314 28556
rect 25994 28864 26314 28890
rect 25994 28556 26000 28864
rect 26308 28556 26314 28864
rect 25994 28550 26314 28556
rect 26994 28864 27314 28890
rect 26994 28556 27000 28864
rect 27308 28556 27314 28864
rect 26994 28550 27314 28556
rect 27994 28864 28314 28890
rect 27994 28556 28000 28864
rect 28308 28556 28314 28864
rect 27994 28550 28314 28556
rect 28994 28864 29314 28890
rect 28994 28556 29000 28864
rect 29308 28556 29314 28864
rect 28994 28550 29314 28556
rect 29994 28864 30314 28890
rect 29994 28556 30000 28864
rect 30308 28556 30314 28864
rect 29994 28550 30314 28556
rect 30994 28864 31314 28890
rect 30994 28556 31000 28864
rect 31308 28556 31314 28864
rect 30994 28550 31314 28556
rect 31994 28864 32314 28890
rect 31994 28556 32000 28864
rect 32308 28556 32314 28864
rect 31994 28550 32314 28556
rect 32994 28864 33314 28890
rect 32994 28556 33000 28864
rect 33308 28556 33314 28864
rect 32994 28550 33314 28556
rect 33994 28864 34314 28890
rect 33994 28556 34000 28864
rect 34308 28556 34314 28864
rect 33994 28550 34314 28556
rect 6620 25567 6638 26131
rect 7202 25567 7220 26131
rect 6620 25561 7220 25567
rect 20275 25954 32275 26000
rect 20275 25948 20324 25954
rect 32216 25948 32275 25954
rect -47625 25517 -47025 25523
rect -72825 16041 -72776 16047
rect -60884 16041 -60825 16047
rect -72825 16000 -60825 16041
rect 20275 16052 20322 25948
rect 32218 16052 32275 25948
rect 20275 16046 20324 16052
rect 32216 16046 32275 16052
rect 20275 16000 32275 16046
rect -21218 15124 -19298 15130
rect -21218 13856 -21212 15124
rect -19304 13856 -19298 15124
rect -21218 13850 -19298 13856
rect -42440 13820 -40660 13850
rect -42440 7880 -42408 13820
rect -40692 7880 -40660 13820
rect -42440 7850 -40660 7880
rect 110 13820 1890 13850
rect 110 7880 142 13820
rect 1858 7880 1890 13820
rect 110 7850 1890 7880
rect -42440 2308 -40660 2350
rect -42440 2298 -42378 2308
rect -40722 2298 -40660 2308
rect -42440 -2298 -42408 2298
rect -40692 -2298 -40660 2298
rect -42440 -2308 -42378 -2298
rect -40722 -2308 -40660 -2298
rect -42440 -2350 -40660 -2308
rect 110 2308 1890 2350
rect 110 2298 172 2308
rect 1828 2298 1890 2308
rect 110 -2298 142 2298
rect 1858 -2298 1890 2298
rect 110 -2308 172 -2298
rect 1828 -2308 1890 -2298
rect 110 -2350 1890 -2308
rect -42440 -7880 -40660 -7850
rect -42440 -13820 -42408 -7880
rect -40692 -13820 -40660 -7880
rect -42440 -13850 -40660 -13820
rect 110 -7880 1890 -7850
rect 110 -13820 142 -7880
rect 1858 -13820 1890 -7880
rect 110 -13850 1890 -13820
rect -72825 -16046 -60825 -16000
rect -72825 -16052 -72776 -16046
rect -60884 -16052 -60825 -16046
rect -72825 -25948 -72778 -16052
rect -60882 -25948 -60825 -16052
rect -72825 -25954 -72776 -25948
rect -60884 -25954 -60825 -25948
rect -72825 -26000 -60825 -25954
rect 20275 -16046 32275 -16000
rect 20275 -16052 20324 -16046
rect 32216 -16052 32275 -16046
rect 20275 -25948 20322 -16052
rect 32218 -25948 32275 -16052
rect 20275 -25954 20324 -25948
rect 32216 -25954 32275 -25948
rect 20275 -26000 32275 -25954
rect -74485 -28556 -74165 -28550
rect -74485 -28864 -74479 -28556
rect -74171 -28864 -74165 -28556
rect -74485 -28890 -74165 -28864
rect -73485 -28556 -73165 -28550
rect -73485 -28864 -73479 -28556
rect -73171 -28864 -73165 -28556
rect -73485 -28890 -73165 -28864
rect -72485 -28556 -72165 -28550
rect -72485 -28864 -72479 -28556
rect -72171 -28864 -72165 -28556
rect -72485 -28890 -72165 -28864
rect -71485 -28556 -71165 -28550
rect -71485 -28864 -71479 -28556
rect -71171 -28864 -71165 -28556
rect -71485 -28890 -71165 -28864
rect -70485 -28556 -70165 -28550
rect -70485 -28864 -70479 -28556
rect -70171 -28864 -70165 -28556
rect -70485 -28890 -70165 -28864
rect -69485 -28556 -69165 -28550
rect -69485 -28864 -69479 -28556
rect -69171 -28864 -69165 -28556
rect -69485 -28890 -69165 -28864
rect -68485 -28556 -68165 -28550
rect -68485 -28864 -68479 -28556
rect -68171 -28864 -68165 -28556
rect -68485 -28890 -68165 -28864
rect -67485 -28556 -67165 -28550
rect -67485 -28864 -67479 -28556
rect -67171 -28864 -67165 -28556
rect -67485 -28890 -67165 -28864
rect -66485 -28556 -66165 -28550
rect -66485 -28864 -66479 -28556
rect -66171 -28864 -66165 -28556
rect -66485 -28890 -66165 -28864
rect -65485 -28556 -65165 -28550
rect -65485 -28864 -65479 -28556
rect -65171 -28864 -65165 -28556
rect -65485 -28890 -65165 -28864
rect -64485 -28556 -64165 -28550
rect -64485 -28864 -64479 -28556
rect -64171 -28864 -64165 -28556
rect -64485 -28890 -64165 -28864
rect -63485 -28556 -63165 -28550
rect -63485 -28864 -63479 -28556
rect -63171 -28864 -63165 -28556
rect -63485 -28890 -63165 -28864
rect -62485 -28556 -62165 -28550
rect -62485 -28864 -62479 -28556
rect -62171 -28864 -62165 -28556
rect -62485 -28890 -62165 -28864
rect -61485 -28556 -61165 -28550
rect -61485 -28864 -61479 -28556
rect -61171 -28864 -61165 -28556
rect -61485 -28890 -61165 -28864
rect -60485 -28556 -60165 -28550
rect -60485 -28864 -60479 -28556
rect -60171 -28864 -60165 -28556
rect -60485 -28890 -60165 -28864
rect -59485 -28556 -59165 -28550
rect -59485 -28864 -59479 -28556
rect -59171 -28864 -59165 -28556
rect -59485 -28890 -59165 -28864
rect -58485 -28556 -58165 -28550
rect -58485 -28864 -58479 -28556
rect -58171 -28864 -58165 -28556
rect -58485 -28890 -58165 -28864
rect -57485 -28556 -57165 -28550
rect -57485 -28864 -57479 -28556
rect -57171 -28864 -57165 -28556
rect -57485 -28890 -57165 -28864
rect -56485 -28556 -56165 -28550
rect -56485 -28864 -56479 -28556
rect -56171 -28864 -56165 -28556
rect -56485 -28890 -56165 -28864
rect -55485 -28556 -55165 -28550
rect -55485 -28864 -55479 -28556
rect -55171 -28864 -55165 -28556
rect -55485 -28890 -55165 -28864
rect -54485 -28556 -54165 -28550
rect -54485 -28864 -54479 -28556
rect -54171 -28864 -54165 -28556
rect -54485 -28890 -54165 -28864
rect -53485 -28556 -53165 -28550
rect -53485 -28864 -53479 -28556
rect -53171 -28864 -53165 -28556
rect -53485 -28890 -53165 -28864
rect -52485 -28556 -52165 -28550
rect -52485 -28864 -52479 -28556
rect -52171 -28864 -52165 -28556
rect -52485 -28890 -52165 -28864
rect -51485 -28556 -51165 -28550
rect -51485 -28864 -51479 -28556
rect -51171 -28864 -51165 -28556
rect -51485 -28890 -51165 -28864
rect -50485 -28556 -50165 -28550
rect -50485 -28864 -50479 -28556
rect -50171 -28864 -50165 -28556
rect -50485 -28890 -50165 -28864
rect -49485 -28556 -49165 -28550
rect -49485 -28864 -49479 -28556
rect -49171 -28864 -49165 -28556
rect -49485 -28890 -49165 -28864
rect 8615 -28556 8935 -28550
rect 8615 -28864 8621 -28556
rect 8929 -28864 8935 -28556
rect 8615 -28890 8935 -28864
rect 9615 -28556 9935 -28550
rect 9615 -28864 9621 -28556
rect 9929 -28864 9935 -28556
rect 9615 -28890 9935 -28864
rect 10615 -28556 10935 -28550
rect 10615 -28864 10621 -28556
rect 10929 -28864 10935 -28556
rect 10615 -28890 10935 -28864
rect 11615 -28556 11935 -28550
rect 11615 -28864 11621 -28556
rect 11929 -28864 11935 -28556
rect 11615 -28890 11935 -28864
rect 12615 -28556 12935 -28550
rect 12615 -28864 12621 -28556
rect 12929 -28864 12935 -28556
rect 12615 -28890 12935 -28864
rect 13615 -28556 13935 -28550
rect 13615 -28864 13621 -28556
rect 13929 -28864 13935 -28556
rect 13615 -28890 13935 -28864
rect 14615 -28556 14935 -28550
rect 14615 -28864 14621 -28556
rect 14929 -28864 14935 -28556
rect 14615 -28890 14935 -28864
rect 15615 -28556 15935 -28550
rect 15615 -28864 15621 -28556
rect 15929 -28864 15935 -28556
rect 15615 -28890 15935 -28864
rect 16615 -28556 16935 -28550
rect 16615 -28864 16621 -28556
rect 16929 -28864 16935 -28556
rect 16615 -28890 16935 -28864
rect 17615 -28556 17935 -28550
rect 17615 -28864 17621 -28556
rect 17929 -28864 17935 -28556
rect 17615 -28890 17935 -28864
rect 18615 -28556 18935 -28550
rect 18615 -28864 18621 -28556
rect 18929 -28864 18935 -28556
rect 18615 -28890 18935 -28864
rect 19615 -28556 19935 -28550
rect 19615 -28864 19621 -28556
rect 19929 -28864 19935 -28556
rect 19615 -28890 19935 -28864
rect 20615 -28556 20935 -28550
rect 20615 -28864 20621 -28556
rect 20929 -28864 20935 -28556
rect 20615 -28890 20935 -28864
rect 21615 -28556 21935 -28550
rect 21615 -28864 21621 -28556
rect 21929 -28864 21935 -28556
rect 21615 -28890 21935 -28864
rect 22615 -28556 22935 -28550
rect 22615 -28864 22621 -28556
rect 22929 -28864 22935 -28556
rect 22615 -28890 22935 -28864
rect 23615 -28556 23935 -28550
rect 23615 -28864 23621 -28556
rect 23929 -28864 23935 -28556
rect 23615 -28890 23935 -28864
rect 24615 -28556 24935 -28550
rect 24615 -28864 24621 -28556
rect 24929 -28864 24935 -28556
rect 24615 -28890 24935 -28864
rect 25615 -28556 25935 -28550
rect 25615 -28864 25621 -28556
rect 25929 -28864 25935 -28556
rect 25615 -28890 25935 -28864
rect 26615 -28556 26935 -28550
rect 26615 -28864 26621 -28556
rect 26929 -28864 26935 -28556
rect 26615 -28890 26935 -28864
rect 27615 -28556 27935 -28550
rect 27615 -28864 27621 -28556
rect 27929 -28864 27935 -28556
rect 27615 -28890 27935 -28864
rect 28615 -28556 28935 -28550
rect 28615 -28864 28621 -28556
rect 28929 -28864 28935 -28556
rect 28615 -28890 28935 -28864
rect 29615 -28556 29935 -28550
rect 29615 -28864 29621 -28556
rect 29929 -28864 29935 -28556
rect 29615 -28890 29935 -28864
rect 30615 -28556 30935 -28550
rect 30615 -28864 30621 -28556
rect 30929 -28864 30935 -28556
rect 30615 -28890 30935 -28864
rect 31615 -28556 31935 -28550
rect 31615 -28864 31621 -28556
rect 31929 -28864 31935 -28556
rect 31615 -28890 31935 -28864
rect 32615 -28556 32935 -28550
rect 32615 -28864 32621 -28556
rect 32929 -28864 32935 -28556
rect 32615 -28890 32935 -28864
rect 33615 -28556 33935 -28550
rect 33615 -28864 33621 -28556
rect 33929 -28864 33935 -28556
rect 33615 -28890 33935 -28864
rect -74825 -28896 -48825 -28890
rect -74825 -29204 -74819 -28896
rect -74511 -28902 -74139 -28896
rect -73511 -28902 -73139 -28896
rect -72511 -28902 -72139 -28896
rect -71511 -28902 -71139 -28896
rect -70511 -28902 -70139 -28896
rect -69511 -28902 -69139 -28896
rect -68511 -28902 -68139 -28896
rect -67511 -28902 -67139 -28896
rect -66511 -28902 -66139 -28896
rect -65511 -28902 -65139 -28896
rect -64511 -28902 -64139 -28896
rect -63511 -28902 -63139 -28896
rect -62511 -28902 -62139 -28896
rect -61511 -28902 -61139 -28896
rect -60511 -28902 -60139 -28896
rect -59511 -28902 -59139 -28896
rect -58511 -28902 -58139 -28896
rect -57511 -28902 -57139 -28896
rect -56511 -28902 -56139 -28896
rect -55511 -28902 -55139 -28896
rect -54511 -28902 -54139 -28896
rect -53511 -28902 -53139 -28896
rect -52511 -28902 -52139 -28896
rect -51511 -28902 -51139 -28896
rect -50511 -28902 -50139 -28896
rect -49511 -28902 -49139 -28896
rect -74511 -29198 -74473 -28902
rect -74177 -29198 -74139 -28902
rect -73511 -29198 -73473 -28902
rect -73177 -29198 -73139 -28902
rect -72511 -29198 -72473 -28902
rect -72177 -29198 -72139 -28902
rect -71511 -29198 -71473 -28902
rect -71177 -29198 -71139 -28902
rect -70511 -29198 -70473 -28902
rect -70177 -29198 -70139 -28902
rect -69511 -29198 -69473 -28902
rect -69177 -29198 -69139 -28902
rect -68511 -29198 -68473 -28902
rect -68177 -29198 -68139 -28902
rect -67511 -29198 -67473 -28902
rect -67177 -29198 -67139 -28902
rect -66511 -29198 -66473 -28902
rect -66177 -29198 -66139 -28902
rect -65511 -29198 -65473 -28902
rect -65177 -29198 -65139 -28902
rect -64511 -29198 -64473 -28902
rect -64177 -29198 -64139 -28902
rect -63511 -29198 -63473 -28902
rect -63177 -29198 -63139 -28902
rect -62511 -29198 -62473 -28902
rect -62177 -29198 -62139 -28902
rect -61511 -29198 -61473 -28902
rect -61177 -29198 -61139 -28902
rect -60511 -29198 -60473 -28902
rect -60177 -29198 -60139 -28902
rect -59511 -29198 -59473 -28902
rect -59177 -29198 -59139 -28902
rect -58511 -29198 -58473 -28902
rect -58177 -29198 -58139 -28902
rect -57511 -29198 -57473 -28902
rect -57177 -29198 -57139 -28902
rect -56511 -29198 -56473 -28902
rect -56177 -29198 -56139 -28902
rect -55511 -29198 -55473 -28902
rect -55177 -29198 -55139 -28902
rect -54511 -29198 -54473 -28902
rect -54177 -29198 -54139 -28902
rect -53511 -29198 -53473 -28902
rect -53177 -29198 -53139 -28902
rect -52511 -29198 -52473 -28902
rect -52177 -29198 -52139 -28902
rect -51511 -29198 -51473 -28902
rect -51177 -29198 -51139 -28902
rect -50511 -29198 -50473 -28902
rect -50177 -29198 -50139 -28902
rect -49511 -29198 -49473 -28902
rect -49177 -29198 -49139 -28902
rect -74511 -29204 -74139 -29198
rect -73511 -29204 -73139 -29198
rect -72511 -29204 -72139 -29198
rect -71511 -29204 -71139 -29198
rect -70511 -29204 -70139 -29198
rect -69511 -29204 -69139 -29198
rect -68511 -29204 -68139 -29198
rect -67511 -29204 -67139 -29198
rect -66511 -29204 -66139 -29198
rect -65511 -29204 -65139 -29198
rect -64511 -29204 -64139 -29198
rect -63511 -29204 -63139 -29198
rect -62511 -29204 -62139 -29198
rect -61511 -29204 -61139 -29198
rect -60511 -29204 -60139 -29198
rect -59511 -29204 -59139 -29198
rect -58511 -29204 -58139 -29198
rect -57511 -29204 -57139 -29198
rect -56511 -29204 -56139 -29198
rect -55511 -29204 -55139 -29198
rect -54511 -29204 -54139 -29198
rect -53511 -29204 -53139 -29198
rect -52511 -29204 -52139 -29198
rect -51511 -29204 -51139 -29198
rect -50511 -29204 -50139 -29198
rect -49511 -29204 -49139 -29198
rect -48831 -29204 -48825 -28896
rect -74825 -29210 -48825 -29204
rect 8275 -28896 34275 -28890
rect 8275 -29204 8281 -28896
rect 8589 -28902 8961 -28896
rect 9589 -28902 9961 -28896
rect 10589 -28902 10961 -28896
rect 11589 -28902 11961 -28896
rect 12589 -28902 12961 -28896
rect 13589 -28902 13961 -28896
rect 14589 -28902 14961 -28896
rect 15589 -28902 15961 -28896
rect 16589 -28902 16961 -28896
rect 17589 -28902 17961 -28896
rect 18589 -28902 18961 -28896
rect 19589 -28902 19961 -28896
rect 20589 -28902 20961 -28896
rect 21589 -28902 21961 -28896
rect 22589 -28902 22961 -28896
rect 23589 -28902 23961 -28896
rect 24589 -28902 24961 -28896
rect 25589 -28902 25961 -28896
rect 26589 -28902 26961 -28896
rect 27589 -28902 27961 -28896
rect 28589 -28902 28961 -28896
rect 29589 -28902 29961 -28896
rect 30589 -28902 30961 -28896
rect 31589 -28902 31961 -28896
rect 32589 -28902 32961 -28896
rect 33589 -28902 33961 -28896
rect 8589 -29198 8627 -28902
rect 8923 -29198 8961 -28902
rect 9589 -29198 9627 -28902
rect 9923 -29198 9961 -28902
rect 10589 -29198 10627 -28902
rect 10923 -29198 10961 -28902
rect 11589 -29198 11627 -28902
rect 11923 -29198 11961 -28902
rect 12589 -29198 12627 -28902
rect 12923 -29198 12961 -28902
rect 13589 -29198 13627 -28902
rect 13923 -29198 13961 -28902
rect 14589 -29198 14627 -28902
rect 14923 -29198 14961 -28902
rect 15589 -29198 15627 -28902
rect 15923 -29198 15961 -28902
rect 16589 -29198 16627 -28902
rect 16923 -29198 16961 -28902
rect 17589 -29198 17627 -28902
rect 17923 -29198 17961 -28902
rect 18589 -29198 18627 -28902
rect 18923 -29198 18961 -28902
rect 19589 -29198 19627 -28902
rect 19923 -29198 19961 -28902
rect 20589 -29198 20627 -28902
rect 20923 -29198 20961 -28902
rect 21589 -29198 21627 -28902
rect 21923 -29198 21961 -28902
rect 22589 -29198 22627 -28902
rect 22923 -29198 22961 -28902
rect 23589 -29198 23627 -28902
rect 23923 -29198 23961 -28902
rect 24589 -29198 24627 -28902
rect 24923 -29198 24961 -28902
rect 25589 -29198 25627 -28902
rect 25923 -29198 25961 -28902
rect 26589 -29198 26627 -28902
rect 26923 -29198 26961 -28902
rect 27589 -29198 27627 -28902
rect 27923 -29198 27961 -28902
rect 28589 -29198 28627 -28902
rect 28923 -29198 28961 -28902
rect 29589 -29198 29627 -28902
rect 29923 -29198 29961 -28902
rect 30589 -29198 30627 -28902
rect 30923 -29198 30961 -28902
rect 31589 -29198 31627 -28902
rect 31923 -29198 31961 -28902
rect 32589 -29198 32627 -28902
rect 32923 -29198 32961 -28902
rect 33589 -29198 33627 -28902
rect 33923 -29198 33961 -28902
rect 8589 -29204 8961 -29198
rect 9589 -29204 9961 -29198
rect 10589 -29204 10961 -29198
rect 11589 -29204 11961 -29198
rect 12589 -29204 12961 -29198
rect 13589 -29204 13961 -29198
rect 14589 -29204 14961 -29198
rect 15589 -29204 15961 -29198
rect 16589 -29204 16961 -29198
rect 17589 -29204 17961 -29198
rect 18589 -29204 18961 -29198
rect 19589 -29204 19961 -29198
rect 20589 -29204 20961 -29198
rect 21589 -29204 21961 -29198
rect 22589 -29204 22961 -29198
rect 23589 -29204 23961 -29198
rect 24589 -29204 24961 -29198
rect 25589 -29204 25961 -29198
rect 26589 -29204 26961 -29198
rect 27589 -29204 27961 -29198
rect 28589 -29204 28961 -29198
rect 29589 -29204 29961 -29198
rect 30589 -29204 30961 -29198
rect 31589 -29204 31961 -29198
rect 32589 -29204 32961 -29198
rect 33589 -29204 33961 -29198
rect 34269 -29204 34275 -28896
rect 8275 -29210 34275 -29204
rect -74485 -29236 -74165 -29210
rect -74485 -29864 -74479 -29236
rect -74171 -29864 -74165 -29236
rect -74485 -29890 -74165 -29864
rect -73485 -29236 -73165 -29210
rect -73485 -29864 -73479 -29236
rect -73171 -29864 -73165 -29236
rect -73485 -29890 -73165 -29864
rect -72485 -29236 -72165 -29210
rect -72485 -29864 -72479 -29236
rect -72171 -29864 -72165 -29236
rect -72485 -29890 -72165 -29864
rect -71485 -29236 -71165 -29210
rect -71485 -29864 -71479 -29236
rect -71171 -29864 -71165 -29236
rect -71485 -29890 -71165 -29864
rect -70485 -29236 -70165 -29210
rect -70485 -29864 -70479 -29236
rect -70171 -29864 -70165 -29236
rect -70485 -29890 -70165 -29864
rect -69485 -29236 -69165 -29210
rect -69485 -29864 -69479 -29236
rect -69171 -29864 -69165 -29236
rect -69485 -29890 -69165 -29864
rect -68485 -29236 -68165 -29210
rect -68485 -29864 -68479 -29236
rect -68171 -29864 -68165 -29236
rect -68485 -29890 -68165 -29864
rect -67485 -29236 -67165 -29210
rect -67485 -29864 -67479 -29236
rect -67171 -29864 -67165 -29236
rect -67485 -29890 -67165 -29864
rect -66485 -29236 -66165 -29210
rect -66485 -29864 -66479 -29236
rect -66171 -29864 -66165 -29236
rect -66485 -29890 -66165 -29864
rect -65485 -29236 -65165 -29210
rect -65485 -29864 -65479 -29236
rect -65171 -29864 -65165 -29236
rect -65485 -29890 -65165 -29864
rect -64485 -29236 -64165 -29210
rect -64485 -29864 -64479 -29236
rect -64171 -29864 -64165 -29236
rect -64485 -29890 -64165 -29864
rect -63485 -29236 -63165 -29210
rect -63485 -29864 -63479 -29236
rect -63171 -29864 -63165 -29236
rect -63485 -29890 -63165 -29864
rect -62485 -29236 -62165 -29210
rect -62485 -29864 -62479 -29236
rect -62171 -29864 -62165 -29236
rect -62485 -29890 -62165 -29864
rect -61485 -29236 -61165 -29210
rect -61485 -29864 -61479 -29236
rect -61171 -29864 -61165 -29236
rect -61485 -29890 -61165 -29864
rect -60485 -29236 -60165 -29210
rect -60485 -29864 -60479 -29236
rect -60171 -29864 -60165 -29236
rect -60485 -29890 -60165 -29864
rect -59485 -29236 -59165 -29210
rect -59485 -29864 -59479 -29236
rect -59171 -29864 -59165 -29236
rect -59485 -29890 -59165 -29864
rect -58485 -29236 -58165 -29210
rect -58485 -29864 -58479 -29236
rect -58171 -29864 -58165 -29236
rect -58485 -29890 -58165 -29864
rect -57485 -29236 -57165 -29210
rect -57485 -29864 -57479 -29236
rect -57171 -29864 -57165 -29236
rect -57485 -29890 -57165 -29864
rect -56485 -29236 -56165 -29210
rect -56485 -29864 -56479 -29236
rect -56171 -29864 -56165 -29236
rect -56485 -29890 -56165 -29864
rect -55485 -29236 -55165 -29210
rect -55485 -29864 -55479 -29236
rect -55171 -29864 -55165 -29236
rect -55485 -29890 -55165 -29864
rect -54485 -29236 -54165 -29210
rect -54485 -29864 -54479 -29236
rect -54171 -29864 -54165 -29236
rect -54485 -29890 -54165 -29864
rect -53485 -29236 -53165 -29210
rect -53485 -29864 -53479 -29236
rect -53171 -29864 -53165 -29236
rect -53485 -29890 -53165 -29864
rect -52485 -29236 -52165 -29210
rect -52485 -29864 -52479 -29236
rect -52171 -29864 -52165 -29236
rect -52485 -29890 -52165 -29864
rect -51485 -29236 -51165 -29210
rect -51485 -29864 -51479 -29236
rect -51171 -29864 -51165 -29236
rect -51485 -29890 -51165 -29864
rect -50485 -29236 -50165 -29210
rect -50485 -29864 -50479 -29236
rect -50171 -29864 -50165 -29236
rect -50485 -29890 -50165 -29864
rect -49485 -29236 -49165 -29210
rect -49485 -29864 -49479 -29236
rect -49171 -29864 -49165 -29236
rect -49485 -29890 -49165 -29864
rect 8615 -29236 8935 -29210
rect 8615 -29864 8621 -29236
rect 8929 -29864 8935 -29236
rect 8615 -29890 8935 -29864
rect 9615 -29236 9935 -29210
rect 9615 -29864 9621 -29236
rect 9929 -29864 9935 -29236
rect 9615 -29890 9935 -29864
rect 10615 -29236 10935 -29210
rect 10615 -29864 10621 -29236
rect 10929 -29864 10935 -29236
rect 10615 -29890 10935 -29864
rect 11615 -29236 11935 -29210
rect 11615 -29864 11621 -29236
rect 11929 -29864 11935 -29236
rect 11615 -29890 11935 -29864
rect 12615 -29236 12935 -29210
rect 12615 -29864 12621 -29236
rect 12929 -29864 12935 -29236
rect 12615 -29890 12935 -29864
rect 13615 -29236 13935 -29210
rect 13615 -29864 13621 -29236
rect 13929 -29864 13935 -29236
rect 13615 -29890 13935 -29864
rect 14615 -29236 14935 -29210
rect 14615 -29864 14621 -29236
rect 14929 -29864 14935 -29236
rect 14615 -29890 14935 -29864
rect 15615 -29236 15935 -29210
rect 15615 -29864 15621 -29236
rect 15929 -29864 15935 -29236
rect 15615 -29890 15935 -29864
rect 16615 -29236 16935 -29210
rect 16615 -29864 16621 -29236
rect 16929 -29864 16935 -29236
rect 16615 -29890 16935 -29864
rect 17615 -29236 17935 -29210
rect 17615 -29864 17621 -29236
rect 17929 -29864 17935 -29236
rect 17615 -29890 17935 -29864
rect 18615 -29236 18935 -29210
rect 18615 -29864 18621 -29236
rect 18929 -29864 18935 -29236
rect 18615 -29890 18935 -29864
rect 19615 -29236 19935 -29210
rect 19615 -29864 19621 -29236
rect 19929 -29864 19935 -29236
rect 19615 -29890 19935 -29864
rect 20615 -29236 20935 -29210
rect 20615 -29864 20621 -29236
rect 20929 -29864 20935 -29236
rect 20615 -29890 20935 -29864
rect 21615 -29236 21935 -29210
rect 21615 -29864 21621 -29236
rect 21929 -29864 21935 -29236
rect 21615 -29890 21935 -29864
rect 22615 -29236 22935 -29210
rect 22615 -29864 22621 -29236
rect 22929 -29864 22935 -29236
rect 22615 -29890 22935 -29864
rect 23615 -29236 23935 -29210
rect 23615 -29864 23621 -29236
rect 23929 -29864 23935 -29236
rect 23615 -29890 23935 -29864
rect 24615 -29236 24935 -29210
rect 24615 -29864 24621 -29236
rect 24929 -29864 24935 -29236
rect 24615 -29890 24935 -29864
rect 25615 -29236 25935 -29210
rect 25615 -29864 25621 -29236
rect 25929 -29864 25935 -29236
rect 25615 -29890 25935 -29864
rect 26615 -29236 26935 -29210
rect 26615 -29864 26621 -29236
rect 26929 -29864 26935 -29236
rect 26615 -29890 26935 -29864
rect 27615 -29236 27935 -29210
rect 27615 -29864 27621 -29236
rect 27929 -29864 27935 -29236
rect 27615 -29890 27935 -29864
rect 28615 -29236 28935 -29210
rect 28615 -29864 28621 -29236
rect 28929 -29864 28935 -29236
rect 28615 -29890 28935 -29864
rect 29615 -29236 29935 -29210
rect 29615 -29864 29621 -29236
rect 29929 -29864 29935 -29236
rect 29615 -29890 29935 -29864
rect 30615 -29236 30935 -29210
rect 30615 -29864 30621 -29236
rect 30929 -29864 30935 -29236
rect 30615 -29890 30935 -29864
rect 31615 -29236 31935 -29210
rect 31615 -29864 31621 -29236
rect 31929 -29864 31935 -29236
rect 31615 -29890 31935 -29864
rect 32615 -29236 32935 -29210
rect 32615 -29864 32621 -29236
rect 32929 -29864 32935 -29236
rect 32615 -29890 32935 -29864
rect 33615 -29236 33935 -29210
rect 33615 -29864 33621 -29236
rect 33929 -29864 33935 -29236
rect 33615 -29890 33935 -29864
rect -74825 -29896 -48825 -29890
rect -74825 -30204 -74819 -29896
rect -74511 -29902 -74139 -29896
rect -73511 -29902 -73139 -29896
rect -72511 -29902 -72139 -29896
rect -71511 -29902 -71139 -29896
rect -70511 -29902 -70139 -29896
rect -69511 -29902 -69139 -29896
rect -68511 -29902 -68139 -29896
rect -67511 -29902 -67139 -29896
rect -66511 -29902 -66139 -29896
rect -65511 -29902 -65139 -29896
rect -64511 -29902 -64139 -29896
rect -63511 -29902 -63139 -29896
rect -62511 -29902 -62139 -29896
rect -61511 -29902 -61139 -29896
rect -60511 -29902 -60139 -29896
rect -59511 -29902 -59139 -29896
rect -58511 -29902 -58139 -29896
rect -57511 -29902 -57139 -29896
rect -56511 -29902 -56139 -29896
rect -55511 -29902 -55139 -29896
rect -54511 -29902 -54139 -29896
rect -53511 -29902 -53139 -29896
rect -52511 -29902 -52139 -29896
rect -51511 -29902 -51139 -29896
rect -50511 -29902 -50139 -29896
rect -49511 -29902 -49139 -29896
rect -74511 -30198 -74473 -29902
rect -74177 -30198 -74139 -29902
rect -73511 -30198 -73473 -29902
rect -73177 -30198 -73139 -29902
rect -72511 -30198 -72473 -29902
rect -72177 -30198 -72139 -29902
rect -71511 -30198 -71473 -29902
rect -71177 -30198 -71139 -29902
rect -70511 -30198 -70473 -29902
rect -70177 -30198 -70139 -29902
rect -69511 -30198 -69473 -29902
rect -69177 -30198 -69139 -29902
rect -68511 -30198 -68473 -29902
rect -68177 -30198 -68139 -29902
rect -67511 -30198 -67473 -29902
rect -67177 -30198 -67139 -29902
rect -66511 -30198 -66473 -29902
rect -66177 -30198 -66139 -29902
rect -65511 -30198 -65473 -29902
rect -65177 -30198 -65139 -29902
rect -64511 -30198 -64473 -29902
rect -64177 -30198 -64139 -29902
rect -63511 -30198 -63473 -29902
rect -63177 -30198 -63139 -29902
rect -62511 -30198 -62473 -29902
rect -62177 -30198 -62139 -29902
rect -61511 -30198 -61473 -29902
rect -61177 -30198 -61139 -29902
rect -60511 -30198 -60473 -29902
rect -60177 -30198 -60139 -29902
rect -59511 -30198 -59473 -29902
rect -59177 -30198 -59139 -29902
rect -58511 -30198 -58473 -29902
rect -58177 -30198 -58139 -29902
rect -57511 -30198 -57473 -29902
rect -57177 -30198 -57139 -29902
rect -56511 -30198 -56473 -29902
rect -56177 -30198 -56139 -29902
rect -55511 -30198 -55473 -29902
rect -55177 -30198 -55139 -29902
rect -54511 -30198 -54473 -29902
rect -54177 -30198 -54139 -29902
rect -53511 -30198 -53473 -29902
rect -53177 -30198 -53139 -29902
rect -52511 -30198 -52473 -29902
rect -52177 -30198 -52139 -29902
rect -51511 -30198 -51473 -29902
rect -51177 -30198 -51139 -29902
rect -50511 -30198 -50473 -29902
rect -50177 -30198 -50139 -29902
rect -49511 -30198 -49473 -29902
rect -49177 -30198 -49139 -29902
rect -74511 -30204 -74139 -30198
rect -73511 -30204 -73139 -30198
rect -72511 -30204 -72139 -30198
rect -71511 -30204 -71139 -30198
rect -70511 -30204 -70139 -30198
rect -69511 -30204 -69139 -30198
rect -68511 -30204 -68139 -30198
rect -67511 -30204 -67139 -30198
rect -66511 -30204 -66139 -30198
rect -65511 -30204 -65139 -30198
rect -64511 -30204 -64139 -30198
rect -63511 -30204 -63139 -30198
rect -62511 -30204 -62139 -30198
rect -61511 -30204 -61139 -30198
rect -60511 -30204 -60139 -30198
rect -59511 -30204 -59139 -30198
rect -58511 -30204 -58139 -30198
rect -57511 -30204 -57139 -30198
rect -56511 -30204 -56139 -30198
rect -55511 -30204 -55139 -30198
rect -54511 -30204 -54139 -30198
rect -53511 -30204 -53139 -30198
rect -52511 -30204 -52139 -30198
rect -51511 -30204 -51139 -30198
rect -50511 -30204 -50139 -30198
rect -49511 -30204 -49139 -30198
rect -48831 -30204 -48825 -29896
rect -74825 -30210 -48825 -30204
rect 8275 -29896 34275 -29890
rect 8275 -30204 8281 -29896
rect 8589 -29902 8961 -29896
rect 9589 -29902 9961 -29896
rect 10589 -29902 10961 -29896
rect 11589 -29902 11961 -29896
rect 12589 -29902 12961 -29896
rect 13589 -29902 13961 -29896
rect 14589 -29902 14961 -29896
rect 15589 -29902 15961 -29896
rect 16589 -29902 16961 -29896
rect 17589 -29902 17961 -29896
rect 18589 -29902 18961 -29896
rect 19589 -29902 19961 -29896
rect 20589 -29902 20961 -29896
rect 21589 -29902 21961 -29896
rect 22589 -29902 22961 -29896
rect 23589 -29902 23961 -29896
rect 24589 -29902 24961 -29896
rect 25589 -29902 25961 -29896
rect 26589 -29902 26961 -29896
rect 27589 -29902 27961 -29896
rect 28589 -29902 28961 -29896
rect 29589 -29902 29961 -29896
rect 30589 -29902 30961 -29896
rect 31589 -29902 31961 -29896
rect 32589 -29902 32961 -29896
rect 33589 -29902 33961 -29896
rect 8589 -30198 8627 -29902
rect 8923 -30198 8961 -29902
rect 9589 -30198 9627 -29902
rect 9923 -30198 9961 -29902
rect 10589 -30198 10627 -29902
rect 10923 -30198 10961 -29902
rect 11589 -30198 11627 -29902
rect 11923 -30198 11961 -29902
rect 12589 -30198 12627 -29902
rect 12923 -30198 12961 -29902
rect 13589 -30198 13627 -29902
rect 13923 -30198 13961 -29902
rect 14589 -30198 14627 -29902
rect 14923 -30198 14961 -29902
rect 15589 -30198 15627 -29902
rect 15923 -30198 15961 -29902
rect 16589 -30198 16627 -29902
rect 16923 -30198 16961 -29902
rect 17589 -30198 17627 -29902
rect 17923 -30198 17961 -29902
rect 18589 -30198 18627 -29902
rect 18923 -30198 18961 -29902
rect 19589 -30198 19627 -29902
rect 19923 -30198 19961 -29902
rect 20589 -30198 20627 -29902
rect 20923 -30198 20961 -29902
rect 21589 -30198 21627 -29902
rect 21923 -30198 21961 -29902
rect 22589 -30198 22627 -29902
rect 22923 -30198 22961 -29902
rect 23589 -30198 23627 -29902
rect 23923 -30198 23961 -29902
rect 24589 -30198 24627 -29902
rect 24923 -30198 24961 -29902
rect 25589 -30198 25627 -29902
rect 25923 -30198 25961 -29902
rect 26589 -30198 26627 -29902
rect 26923 -30198 26961 -29902
rect 27589 -30198 27627 -29902
rect 27923 -30198 27961 -29902
rect 28589 -30198 28627 -29902
rect 28923 -30198 28961 -29902
rect 29589 -30198 29627 -29902
rect 29923 -30198 29961 -29902
rect 30589 -30198 30627 -29902
rect 30923 -30198 30961 -29902
rect 31589 -30198 31627 -29902
rect 31923 -30198 31961 -29902
rect 32589 -30198 32627 -29902
rect 32923 -30198 32961 -29902
rect 33589 -30198 33627 -29902
rect 33923 -30198 33961 -29902
rect 8589 -30204 8961 -30198
rect 9589 -30204 9961 -30198
rect 10589 -30204 10961 -30198
rect 11589 -30204 11961 -30198
rect 12589 -30204 12961 -30198
rect 13589 -30204 13961 -30198
rect 14589 -30204 14961 -30198
rect 15589 -30204 15961 -30198
rect 16589 -30204 16961 -30198
rect 17589 -30204 17961 -30198
rect 18589 -30204 18961 -30198
rect 19589 -30204 19961 -30198
rect 20589 -30204 20961 -30198
rect 21589 -30204 21961 -30198
rect 22589 -30204 22961 -30198
rect 23589 -30204 23961 -30198
rect 24589 -30204 24961 -30198
rect 25589 -30204 25961 -30198
rect 26589 -30204 26961 -30198
rect 27589 -30204 27961 -30198
rect 28589 -30204 28961 -30198
rect 29589 -30204 29961 -30198
rect 30589 -30204 30961 -30198
rect 31589 -30204 31961 -30198
rect 32589 -30204 32961 -30198
rect 33589 -30204 33961 -30198
rect 34269 -30204 34275 -29896
rect 8275 -30210 34275 -30204
rect -74485 -30236 -74165 -30210
rect -74485 -30864 -74479 -30236
rect -74171 -30864 -74165 -30236
rect -74485 -30890 -74165 -30864
rect -73485 -30236 -73165 -30210
rect -73485 -30864 -73479 -30236
rect -73171 -30864 -73165 -30236
rect -73485 -30890 -73165 -30864
rect -72485 -30236 -72165 -30210
rect -72485 -30864 -72479 -30236
rect -72171 -30864 -72165 -30236
rect -72485 -30890 -72165 -30864
rect -71485 -30236 -71165 -30210
rect -71485 -30864 -71479 -30236
rect -71171 -30864 -71165 -30236
rect -71485 -30890 -71165 -30864
rect -70485 -30236 -70165 -30210
rect -70485 -30864 -70479 -30236
rect -70171 -30864 -70165 -30236
rect -70485 -30890 -70165 -30864
rect -69485 -30236 -69165 -30210
rect -69485 -30864 -69479 -30236
rect -69171 -30864 -69165 -30236
rect -69485 -30890 -69165 -30864
rect -68485 -30236 -68165 -30210
rect -68485 -30864 -68479 -30236
rect -68171 -30864 -68165 -30236
rect -68485 -30890 -68165 -30864
rect -67485 -30236 -67165 -30210
rect -67485 -30864 -67479 -30236
rect -67171 -30864 -67165 -30236
rect -67485 -30890 -67165 -30864
rect -66485 -30236 -66165 -30210
rect -66485 -30864 -66479 -30236
rect -66171 -30864 -66165 -30236
rect -66485 -30890 -66165 -30864
rect -65485 -30236 -65165 -30210
rect -65485 -30864 -65479 -30236
rect -65171 -30864 -65165 -30236
rect -65485 -30890 -65165 -30864
rect -64485 -30236 -64165 -30210
rect -64485 -30864 -64479 -30236
rect -64171 -30864 -64165 -30236
rect -64485 -30890 -64165 -30864
rect -63485 -30236 -63165 -30210
rect -63485 -30864 -63479 -30236
rect -63171 -30864 -63165 -30236
rect -63485 -30890 -63165 -30864
rect -62485 -30236 -62165 -30210
rect -62485 -30864 -62479 -30236
rect -62171 -30864 -62165 -30236
rect -62485 -30890 -62165 -30864
rect -61485 -30236 -61165 -30210
rect -61485 -30864 -61479 -30236
rect -61171 -30864 -61165 -30236
rect -61485 -30890 -61165 -30864
rect -60485 -30236 -60165 -30210
rect -60485 -30864 -60479 -30236
rect -60171 -30864 -60165 -30236
rect -60485 -30890 -60165 -30864
rect -59485 -30236 -59165 -30210
rect -59485 -30864 -59479 -30236
rect -59171 -30864 -59165 -30236
rect -59485 -30890 -59165 -30864
rect -58485 -30236 -58165 -30210
rect -58485 -30864 -58479 -30236
rect -58171 -30864 -58165 -30236
rect -58485 -30890 -58165 -30864
rect -57485 -30236 -57165 -30210
rect -57485 -30864 -57479 -30236
rect -57171 -30864 -57165 -30236
rect -57485 -30890 -57165 -30864
rect -56485 -30236 -56165 -30210
rect -56485 -30864 -56479 -30236
rect -56171 -30864 -56165 -30236
rect -56485 -30890 -56165 -30864
rect -55485 -30236 -55165 -30210
rect -55485 -30864 -55479 -30236
rect -55171 -30864 -55165 -30236
rect -55485 -30890 -55165 -30864
rect -54485 -30236 -54165 -30210
rect -54485 -30864 -54479 -30236
rect -54171 -30864 -54165 -30236
rect -54485 -30890 -54165 -30864
rect -53485 -30236 -53165 -30210
rect -53485 -30864 -53479 -30236
rect -53171 -30864 -53165 -30236
rect -53485 -30890 -53165 -30864
rect -52485 -30236 -52165 -30210
rect -52485 -30864 -52479 -30236
rect -52171 -30864 -52165 -30236
rect -52485 -30890 -52165 -30864
rect -51485 -30236 -51165 -30210
rect -51485 -30864 -51479 -30236
rect -51171 -30864 -51165 -30236
rect -51485 -30890 -51165 -30864
rect -50485 -30236 -50165 -30210
rect -50485 -30864 -50479 -30236
rect -50171 -30864 -50165 -30236
rect -50485 -30890 -50165 -30864
rect -49485 -30236 -49165 -30210
rect -49485 -30864 -49479 -30236
rect -49171 -30864 -49165 -30236
rect -49485 -30890 -49165 -30864
rect 8615 -30236 8935 -30210
rect 8615 -30864 8621 -30236
rect 8929 -30864 8935 -30236
rect 8615 -30890 8935 -30864
rect 9615 -30236 9935 -30210
rect 9615 -30864 9621 -30236
rect 9929 -30864 9935 -30236
rect 9615 -30890 9935 -30864
rect 10615 -30236 10935 -30210
rect 10615 -30864 10621 -30236
rect 10929 -30864 10935 -30236
rect 10615 -30890 10935 -30864
rect 11615 -30236 11935 -30210
rect 11615 -30864 11621 -30236
rect 11929 -30864 11935 -30236
rect 11615 -30890 11935 -30864
rect 12615 -30236 12935 -30210
rect 12615 -30864 12621 -30236
rect 12929 -30864 12935 -30236
rect 12615 -30890 12935 -30864
rect 13615 -30236 13935 -30210
rect 13615 -30864 13621 -30236
rect 13929 -30864 13935 -30236
rect 13615 -30890 13935 -30864
rect 14615 -30236 14935 -30210
rect 14615 -30864 14621 -30236
rect 14929 -30864 14935 -30236
rect 14615 -30890 14935 -30864
rect 15615 -30236 15935 -30210
rect 15615 -30864 15621 -30236
rect 15929 -30864 15935 -30236
rect 15615 -30890 15935 -30864
rect 16615 -30236 16935 -30210
rect 16615 -30864 16621 -30236
rect 16929 -30864 16935 -30236
rect 16615 -30890 16935 -30864
rect 17615 -30236 17935 -30210
rect 17615 -30864 17621 -30236
rect 17929 -30864 17935 -30236
rect 17615 -30890 17935 -30864
rect 18615 -30236 18935 -30210
rect 18615 -30864 18621 -30236
rect 18929 -30864 18935 -30236
rect 18615 -30890 18935 -30864
rect 19615 -30236 19935 -30210
rect 19615 -30864 19621 -30236
rect 19929 -30864 19935 -30236
rect 19615 -30890 19935 -30864
rect 20615 -30236 20935 -30210
rect 20615 -30864 20621 -30236
rect 20929 -30864 20935 -30236
rect 20615 -30890 20935 -30864
rect 21615 -30236 21935 -30210
rect 21615 -30864 21621 -30236
rect 21929 -30864 21935 -30236
rect 21615 -30890 21935 -30864
rect 22615 -30236 22935 -30210
rect 22615 -30864 22621 -30236
rect 22929 -30864 22935 -30236
rect 22615 -30890 22935 -30864
rect 23615 -30236 23935 -30210
rect 23615 -30864 23621 -30236
rect 23929 -30864 23935 -30236
rect 23615 -30890 23935 -30864
rect 24615 -30236 24935 -30210
rect 24615 -30864 24621 -30236
rect 24929 -30864 24935 -30236
rect 24615 -30890 24935 -30864
rect 25615 -30236 25935 -30210
rect 25615 -30864 25621 -30236
rect 25929 -30864 25935 -30236
rect 25615 -30890 25935 -30864
rect 26615 -30236 26935 -30210
rect 26615 -30864 26621 -30236
rect 26929 -30864 26935 -30236
rect 26615 -30890 26935 -30864
rect 27615 -30236 27935 -30210
rect 27615 -30864 27621 -30236
rect 27929 -30864 27935 -30236
rect 27615 -30890 27935 -30864
rect 28615 -30236 28935 -30210
rect 28615 -30864 28621 -30236
rect 28929 -30864 28935 -30236
rect 28615 -30890 28935 -30864
rect 29615 -30236 29935 -30210
rect 29615 -30864 29621 -30236
rect 29929 -30864 29935 -30236
rect 29615 -30890 29935 -30864
rect 30615 -30236 30935 -30210
rect 30615 -30864 30621 -30236
rect 30929 -30864 30935 -30236
rect 30615 -30890 30935 -30864
rect 31615 -30236 31935 -30210
rect 31615 -30864 31621 -30236
rect 31929 -30864 31935 -30236
rect 31615 -30890 31935 -30864
rect 32615 -30236 32935 -30210
rect 32615 -30864 32621 -30236
rect 32929 -30864 32935 -30236
rect 32615 -30890 32935 -30864
rect 33615 -30236 33935 -30210
rect 33615 -30864 33621 -30236
rect 33929 -30864 33935 -30236
rect 33615 -30890 33935 -30864
rect -74825 -30896 -48825 -30890
rect -74825 -31204 -74819 -30896
rect -74511 -30902 -74139 -30896
rect -73511 -30902 -73139 -30896
rect -72511 -30902 -72139 -30896
rect -71511 -30902 -71139 -30896
rect -70511 -30902 -70139 -30896
rect -69511 -30902 -69139 -30896
rect -68511 -30902 -68139 -30896
rect -67511 -30902 -67139 -30896
rect -66511 -30902 -66139 -30896
rect -65511 -30902 -65139 -30896
rect -64511 -30902 -64139 -30896
rect -63511 -30902 -63139 -30896
rect -62511 -30902 -62139 -30896
rect -61511 -30902 -61139 -30896
rect -60511 -30902 -60139 -30896
rect -59511 -30902 -59139 -30896
rect -58511 -30902 -58139 -30896
rect -57511 -30902 -57139 -30896
rect -56511 -30902 -56139 -30896
rect -55511 -30902 -55139 -30896
rect -54511 -30902 -54139 -30896
rect -53511 -30902 -53139 -30896
rect -52511 -30902 -52139 -30896
rect -51511 -30902 -51139 -30896
rect -50511 -30902 -50139 -30896
rect -49511 -30902 -49139 -30896
rect -74511 -31198 -74473 -30902
rect -74177 -31198 -74139 -30902
rect -73511 -31198 -73473 -30902
rect -73177 -31198 -73139 -30902
rect -72511 -31198 -72473 -30902
rect -72177 -31198 -72139 -30902
rect -71511 -31198 -71473 -30902
rect -71177 -31198 -71139 -30902
rect -70511 -31198 -70473 -30902
rect -70177 -31198 -70139 -30902
rect -69511 -31198 -69473 -30902
rect -69177 -31198 -69139 -30902
rect -68511 -31198 -68473 -30902
rect -68177 -31198 -68139 -30902
rect -67511 -31198 -67473 -30902
rect -67177 -31198 -67139 -30902
rect -66511 -31198 -66473 -30902
rect -66177 -31198 -66139 -30902
rect -65511 -31198 -65473 -30902
rect -65177 -31198 -65139 -30902
rect -64511 -31198 -64473 -30902
rect -64177 -31198 -64139 -30902
rect -63511 -31198 -63473 -30902
rect -63177 -31198 -63139 -30902
rect -62511 -31198 -62473 -30902
rect -62177 -31198 -62139 -30902
rect -61511 -31198 -61473 -30902
rect -61177 -31198 -61139 -30902
rect -60511 -31198 -60473 -30902
rect -60177 -31198 -60139 -30902
rect -59511 -31198 -59473 -30902
rect -59177 -31198 -59139 -30902
rect -58511 -31198 -58473 -30902
rect -58177 -31198 -58139 -30902
rect -57511 -31198 -57473 -30902
rect -57177 -31198 -57139 -30902
rect -56511 -31198 -56473 -30902
rect -56177 -31198 -56139 -30902
rect -55511 -31198 -55473 -30902
rect -55177 -31198 -55139 -30902
rect -54511 -31198 -54473 -30902
rect -54177 -31198 -54139 -30902
rect -53511 -31198 -53473 -30902
rect -53177 -31198 -53139 -30902
rect -52511 -31198 -52473 -30902
rect -52177 -31198 -52139 -30902
rect -51511 -31198 -51473 -30902
rect -51177 -31198 -51139 -30902
rect -50511 -31198 -50473 -30902
rect -50177 -31198 -50139 -30902
rect -49511 -31198 -49473 -30902
rect -49177 -31198 -49139 -30902
rect -74511 -31204 -74139 -31198
rect -73511 -31204 -73139 -31198
rect -72511 -31204 -72139 -31198
rect -71511 -31204 -71139 -31198
rect -70511 -31204 -70139 -31198
rect -69511 -31204 -69139 -31198
rect -68511 -31204 -68139 -31198
rect -67511 -31204 -67139 -31198
rect -66511 -31204 -66139 -31198
rect -65511 -31204 -65139 -31198
rect -64511 -31204 -64139 -31198
rect -63511 -31204 -63139 -31198
rect -62511 -31204 -62139 -31198
rect -61511 -31204 -61139 -31198
rect -60511 -31204 -60139 -31198
rect -59511 -31204 -59139 -31198
rect -58511 -31204 -58139 -31198
rect -57511 -31204 -57139 -31198
rect -56511 -31204 -56139 -31198
rect -55511 -31204 -55139 -31198
rect -54511 -31204 -54139 -31198
rect -53511 -31204 -53139 -31198
rect -52511 -31204 -52139 -31198
rect -51511 -31204 -51139 -31198
rect -50511 -31204 -50139 -31198
rect -49511 -31204 -49139 -31198
rect -48831 -31204 -48825 -30896
rect -74825 -31210 -48825 -31204
rect 8275 -30896 34275 -30890
rect 8275 -31204 8281 -30896
rect 8589 -30902 8961 -30896
rect 9589 -30902 9961 -30896
rect 10589 -30902 10961 -30896
rect 11589 -30902 11961 -30896
rect 12589 -30902 12961 -30896
rect 13589 -30902 13961 -30896
rect 14589 -30902 14961 -30896
rect 15589 -30902 15961 -30896
rect 16589 -30902 16961 -30896
rect 17589 -30902 17961 -30896
rect 18589 -30902 18961 -30896
rect 19589 -30902 19961 -30896
rect 20589 -30902 20961 -30896
rect 21589 -30902 21961 -30896
rect 22589 -30902 22961 -30896
rect 23589 -30902 23961 -30896
rect 24589 -30902 24961 -30896
rect 25589 -30902 25961 -30896
rect 26589 -30902 26961 -30896
rect 27589 -30902 27961 -30896
rect 28589 -30902 28961 -30896
rect 29589 -30902 29961 -30896
rect 30589 -30902 30961 -30896
rect 31589 -30902 31961 -30896
rect 32589 -30902 32961 -30896
rect 33589 -30902 33961 -30896
rect 8589 -31198 8627 -30902
rect 8923 -31198 8961 -30902
rect 9589 -31198 9627 -30902
rect 9923 -31198 9961 -30902
rect 10589 -31198 10627 -30902
rect 10923 -31198 10961 -30902
rect 11589 -31198 11627 -30902
rect 11923 -31198 11961 -30902
rect 12589 -31198 12627 -30902
rect 12923 -31198 12961 -30902
rect 13589 -31198 13627 -30902
rect 13923 -31198 13961 -30902
rect 14589 -31198 14627 -30902
rect 14923 -31198 14961 -30902
rect 15589 -31198 15627 -30902
rect 15923 -31198 15961 -30902
rect 16589 -31198 16627 -30902
rect 16923 -31198 16961 -30902
rect 17589 -31198 17627 -30902
rect 17923 -31198 17961 -30902
rect 18589 -31198 18627 -30902
rect 18923 -31198 18961 -30902
rect 19589 -31198 19627 -30902
rect 19923 -31198 19961 -30902
rect 20589 -31198 20627 -30902
rect 20923 -31198 20961 -30902
rect 21589 -31198 21627 -30902
rect 21923 -31198 21961 -30902
rect 22589 -31198 22627 -30902
rect 22923 -31198 22961 -30902
rect 23589 -31198 23627 -30902
rect 23923 -31198 23961 -30902
rect 24589 -31198 24627 -30902
rect 24923 -31198 24961 -30902
rect 25589 -31198 25627 -30902
rect 25923 -31198 25961 -30902
rect 26589 -31198 26627 -30902
rect 26923 -31198 26961 -30902
rect 27589 -31198 27627 -30902
rect 27923 -31198 27961 -30902
rect 28589 -31198 28627 -30902
rect 28923 -31198 28961 -30902
rect 29589 -31198 29627 -30902
rect 29923 -31198 29961 -30902
rect 30589 -31198 30627 -30902
rect 30923 -31198 30961 -30902
rect 31589 -31198 31627 -30902
rect 31923 -31198 31961 -30902
rect 32589 -31198 32627 -30902
rect 32923 -31198 32961 -30902
rect 33589 -31198 33627 -30902
rect 33923 -31198 33961 -30902
rect 8589 -31204 8961 -31198
rect 9589 -31204 9961 -31198
rect 10589 -31204 10961 -31198
rect 11589 -31204 11961 -31198
rect 12589 -31204 12961 -31198
rect 13589 -31204 13961 -31198
rect 14589 -31204 14961 -31198
rect 15589 -31204 15961 -31198
rect 16589 -31204 16961 -31198
rect 17589 -31204 17961 -31198
rect 18589 -31204 18961 -31198
rect 19589 -31204 19961 -31198
rect 20589 -31204 20961 -31198
rect 21589 -31204 21961 -31198
rect 22589 -31204 22961 -31198
rect 23589 -31204 23961 -31198
rect 24589 -31204 24961 -31198
rect 25589 -31204 25961 -31198
rect 26589 -31204 26961 -31198
rect 27589 -31204 27961 -31198
rect 28589 -31204 28961 -31198
rect 29589 -31204 29961 -31198
rect 30589 -31204 30961 -31198
rect 31589 -31204 31961 -31198
rect 32589 -31204 32961 -31198
rect 33589 -31204 33961 -31198
rect 34269 -31204 34275 -30896
rect 8275 -31210 34275 -31204
rect -74485 -31236 -74165 -31210
rect -74485 -31864 -74479 -31236
rect -74171 -31864 -74165 -31236
rect -74485 -31890 -74165 -31864
rect -73485 -31236 -73165 -31210
rect -73485 -31864 -73479 -31236
rect -73171 -31864 -73165 -31236
rect -73485 -31890 -73165 -31864
rect -72485 -31236 -72165 -31210
rect -72485 -31864 -72479 -31236
rect -72171 -31864 -72165 -31236
rect -72485 -31890 -72165 -31864
rect -71485 -31236 -71165 -31210
rect -71485 -31864 -71479 -31236
rect -71171 -31864 -71165 -31236
rect -71485 -31890 -71165 -31864
rect -70485 -31236 -70165 -31210
rect -70485 -31864 -70479 -31236
rect -70171 -31864 -70165 -31236
rect -70485 -31890 -70165 -31864
rect -69485 -31236 -69165 -31210
rect -69485 -31864 -69479 -31236
rect -69171 -31864 -69165 -31236
rect -69485 -31890 -69165 -31864
rect -68485 -31236 -68165 -31210
rect -68485 -31864 -68479 -31236
rect -68171 -31864 -68165 -31236
rect -68485 -31890 -68165 -31864
rect -67485 -31236 -67165 -31210
rect -67485 -31864 -67479 -31236
rect -67171 -31864 -67165 -31236
rect -67485 -31890 -67165 -31864
rect -66485 -31236 -66165 -31210
rect -66485 -31864 -66479 -31236
rect -66171 -31864 -66165 -31236
rect -66485 -31890 -66165 -31864
rect -65485 -31236 -65165 -31210
rect -65485 -31864 -65479 -31236
rect -65171 -31864 -65165 -31236
rect -65485 -31890 -65165 -31864
rect -64485 -31236 -64165 -31210
rect -64485 -31864 -64479 -31236
rect -64171 -31864 -64165 -31236
rect -64485 -31890 -64165 -31864
rect -63485 -31236 -63165 -31210
rect -63485 -31864 -63479 -31236
rect -63171 -31864 -63165 -31236
rect -63485 -31890 -63165 -31864
rect -62485 -31236 -62165 -31210
rect -62485 -31864 -62479 -31236
rect -62171 -31864 -62165 -31236
rect -62485 -31890 -62165 -31864
rect -61485 -31236 -61165 -31210
rect -61485 -31864 -61479 -31236
rect -61171 -31864 -61165 -31236
rect -61485 -31890 -61165 -31864
rect -60485 -31236 -60165 -31210
rect -60485 -31864 -60479 -31236
rect -60171 -31864 -60165 -31236
rect -60485 -31890 -60165 -31864
rect -59485 -31236 -59165 -31210
rect -59485 -31864 -59479 -31236
rect -59171 -31864 -59165 -31236
rect -59485 -31890 -59165 -31864
rect -58485 -31236 -58165 -31210
rect -58485 -31864 -58479 -31236
rect -58171 -31864 -58165 -31236
rect -58485 -31890 -58165 -31864
rect -57485 -31236 -57165 -31210
rect -57485 -31864 -57479 -31236
rect -57171 -31864 -57165 -31236
rect -57485 -31890 -57165 -31864
rect -56485 -31236 -56165 -31210
rect -56485 -31864 -56479 -31236
rect -56171 -31864 -56165 -31236
rect -56485 -31890 -56165 -31864
rect -55485 -31236 -55165 -31210
rect -55485 -31864 -55479 -31236
rect -55171 -31864 -55165 -31236
rect -55485 -31890 -55165 -31864
rect -54485 -31236 -54165 -31210
rect -54485 -31864 -54479 -31236
rect -54171 -31864 -54165 -31236
rect -54485 -31890 -54165 -31864
rect -53485 -31236 -53165 -31210
rect -53485 -31864 -53479 -31236
rect -53171 -31864 -53165 -31236
rect -53485 -31890 -53165 -31864
rect -52485 -31236 -52165 -31210
rect -52485 -31864 -52479 -31236
rect -52171 -31864 -52165 -31236
rect -52485 -31890 -52165 -31864
rect -51485 -31236 -51165 -31210
rect -51485 -31864 -51479 -31236
rect -51171 -31864 -51165 -31236
rect -51485 -31890 -51165 -31864
rect -50485 -31236 -50165 -31210
rect -50485 -31864 -50479 -31236
rect -50171 -31864 -50165 -31236
rect -50485 -31890 -50165 -31864
rect -49485 -31236 -49165 -31210
rect -49485 -31864 -49479 -31236
rect -49171 -31864 -49165 -31236
rect -49485 -31890 -49165 -31864
rect 8615 -31236 8935 -31210
rect 8615 -31864 8621 -31236
rect 8929 -31864 8935 -31236
rect 8615 -31890 8935 -31864
rect 9615 -31236 9935 -31210
rect 9615 -31864 9621 -31236
rect 9929 -31864 9935 -31236
rect 9615 -31890 9935 -31864
rect 10615 -31236 10935 -31210
rect 10615 -31864 10621 -31236
rect 10929 -31864 10935 -31236
rect 10615 -31890 10935 -31864
rect 11615 -31236 11935 -31210
rect 11615 -31864 11621 -31236
rect 11929 -31864 11935 -31236
rect 11615 -31890 11935 -31864
rect 12615 -31236 12935 -31210
rect 12615 -31864 12621 -31236
rect 12929 -31864 12935 -31236
rect 12615 -31890 12935 -31864
rect 13615 -31236 13935 -31210
rect 13615 -31864 13621 -31236
rect 13929 -31864 13935 -31236
rect 13615 -31890 13935 -31864
rect 14615 -31236 14935 -31210
rect 14615 -31864 14621 -31236
rect 14929 -31864 14935 -31236
rect 14615 -31890 14935 -31864
rect 15615 -31236 15935 -31210
rect 15615 -31864 15621 -31236
rect 15929 -31864 15935 -31236
rect 15615 -31890 15935 -31864
rect 16615 -31236 16935 -31210
rect 16615 -31864 16621 -31236
rect 16929 -31864 16935 -31236
rect 16615 -31890 16935 -31864
rect 17615 -31236 17935 -31210
rect 17615 -31864 17621 -31236
rect 17929 -31864 17935 -31236
rect 17615 -31890 17935 -31864
rect 18615 -31236 18935 -31210
rect 18615 -31864 18621 -31236
rect 18929 -31864 18935 -31236
rect 18615 -31890 18935 -31864
rect 19615 -31236 19935 -31210
rect 19615 -31864 19621 -31236
rect 19929 -31864 19935 -31236
rect 19615 -31890 19935 -31864
rect 20615 -31236 20935 -31210
rect 20615 -31864 20621 -31236
rect 20929 -31864 20935 -31236
rect 20615 -31890 20935 -31864
rect 21615 -31236 21935 -31210
rect 21615 -31864 21621 -31236
rect 21929 -31864 21935 -31236
rect 21615 -31890 21935 -31864
rect 22615 -31236 22935 -31210
rect 22615 -31864 22621 -31236
rect 22929 -31864 22935 -31236
rect 22615 -31890 22935 -31864
rect 23615 -31236 23935 -31210
rect 23615 -31864 23621 -31236
rect 23929 -31864 23935 -31236
rect 23615 -31890 23935 -31864
rect 24615 -31236 24935 -31210
rect 24615 -31864 24621 -31236
rect 24929 -31864 24935 -31236
rect 24615 -31890 24935 -31864
rect 25615 -31236 25935 -31210
rect 25615 -31864 25621 -31236
rect 25929 -31864 25935 -31236
rect 25615 -31890 25935 -31864
rect 26615 -31236 26935 -31210
rect 26615 -31864 26621 -31236
rect 26929 -31864 26935 -31236
rect 26615 -31890 26935 -31864
rect 27615 -31236 27935 -31210
rect 27615 -31864 27621 -31236
rect 27929 -31864 27935 -31236
rect 27615 -31890 27935 -31864
rect 28615 -31236 28935 -31210
rect 28615 -31864 28621 -31236
rect 28929 -31864 28935 -31236
rect 28615 -31890 28935 -31864
rect 29615 -31236 29935 -31210
rect 29615 -31864 29621 -31236
rect 29929 -31864 29935 -31236
rect 29615 -31890 29935 -31864
rect 30615 -31236 30935 -31210
rect 30615 -31864 30621 -31236
rect 30929 -31864 30935 -31236
rect 30615 -31890 30935 -31864
rect 31615 -31236 31935 -31210
rect 31615 -31864 31621 -31236
rect 31929 -31864 31935 -31236
rect 31615 -31890 31935 -31864
rect 32615 -31236 32935 -31210
rect 32615 -31864 32621 -31236
rect 32929 -31864 32935 -31236
rect 32615 -31890 32935 -31864
rect 33615 -31236 33935 -31210
rect 33615 -31864 33621 -31236
rect 33929 -31864 33935 -31236
rect 33615 -31890 33935 -31864
rect -74825 -31896 -48825 -31890
rect -74825 -32204 -74819 -31896
rect -74511 -31902 -74139 -31896
rect -73511 -31902 -73139 -31896
rect -72511 -31902 -72139 -31896
rect -71511 -31902 -71139 -31896
rect -70511 -31902 -70139 -31896
rect -69511 -31902 -69139 -31896
rect -68511 -31902 -68139 -31896
rect -67511 -31902 -67139 -31896
rect -66511 -31902 -66139 -31896
rect -65511 -31902 -65139 -31896
rect -64511 -31902 -64139 -31896
rect -63511 -31902 -63139 -31896
rect -62511 -31902 -62139 -31896
rect -61511 -31902 -61139 -31896
rect -60511 -31902 -60139 -31896
rect -59511 -31902 -59139 -31896
rect -58511 -31902 -58139 -31896
rect -57511 -31902 -57139 -31896
rect -56511 -31902 -56139 -31896
rect -55511 -31902 -55139 -31896
rect -54511 -31902 -54139 -31896
rect -53511 -31902 -53139 -31896
rect -52511 -31902 -52139 -31896
rect -51511 -31902 -51139 -31896
rect -50511 -31902 -50139 -31896
rect -49511 -31902 -49139 -31896
rect -74511 -32198 -74473 -31902
rect -74177 -32198 -74139 -31902
rect -73511 -32198 -73473 -31902
rect -73177 -32198 -73139 -31902
rect -72511 -32198 -72473 -31902
rect -72177 -32198 -72139 -31902
rect -71511 -32198 -71473 -31902
rect -71177 -32198 -71139 -31902
rect -70511 -32198 -70473 -31902
rect -70177 -32198 -70139 -31902
rect -69511 -32198 -69473 -31902
rect -69177 -32198 -69139 -31902
rect -68511 -32198 -68473 -31902
rect -68177 -32198 -68139 -31902
rect -67511 -32198 -67473 -31902
rect -67177 -32198 -67139 -31902
rect -66511 -32198 -66473 -31902
rect -66177 -32198 -66139 -31902
rect -65511 -32198 -65473 -31902
rect -65177 -32198 -65139 -31902
rect -64511 -32198 -64473 -31902
rect -64177 -32198 -64139 -31902
rect -63511 -32198 -63473 -31902
rect -63177 -32198 -63139 -31902
rect -62511 -32198 -62473 -31902
rect -62177 -32198 -62139 -31902
rect -61511 -32198 -61473 -31902
rect -61177 -32198 -61139 -31902
rect -60511 -32198 -60473 -31902
rect -60177 -32198 -60139 -31902
rect -59511 -32198 -59473 -31902
rect -59177 -32198 -59139 -31902
rect -58511 -32198 -58473 -31902
rect -58177 -32198 -58139 -31902
rect -57511 -32198 -57473 -31902
rect -57177 -32198 -57139 -31902
rect -56511 -32198 -56473 -31902
rect -56177 -32198 -56139 -31902
rect -55511 -32198 -55473 -31902
rect -55177 -32198 -55139 -31902
rect -54511 -32198 -54473 -31902
rect -54177 -32198 -54139 -31902
rect -53511 -32198 -53473 -31902
rect -53177 -32198 -53139 -31902
rect -52511 -32198 -52473 -31902
rect -52177 -32198 -52139 -31902
rect -51511 -32198 -51473 -31902
rect -51177 -32198 -51139 -31902
rect -50511 -32198 -50473 -31902
rect -50177 -32198 -50139 -31902
rect -49511 -32198 -49473 -31902
rect -49177 -32198 -49139 -31902
rect -74511 -32204 -74139 -32198
rect -73511 -32204 -73139 -32198
rect -72511 -32204 -72139 -32198
rect -71511 -32204 -71139 -32198
rect -70511 -32204 -70139 -32198
rect -69511 -32204 -69139 -32198
rect -68511 -32204 -68139 -32198
rect -67511 -32204 -67139 -32198
rect -66511 -32204 -66139 -32198
rect -65511 -32204 -65139 -32198
rect -64511 -32204 -64139 -32198
rect -63511 -32204 -63139 -32198
rect -62511 -32204 -62139 -32198
rect -61511 -32204 -61139 -32198
rect -60511 -32204 -60139 -32198
rect -59511 -32204 -59139 -32198
rect -58511 -32204 -58139 -32198
rect -57511 -32204 -57139 -32198
rect -56511 -32204 -56139 -32198
rect -55511 -32204 -55139 -32198
rect -54511 -32204 -54139 -32198
rect -53511 -32204 -53139 -32198
rect -52511 -32204 -52139 -32198
rect -51511 -32204 -51139 -32198
rect -50511 -32204 -50139 -32198
rect -49511 -32204 -49139 -32198
rect -48831 -32204 -48825 -31896
rect -74825 -32210 -48825 -32204
rect 8275 -31896 34275 -31890
rect 8275 -32204 8281 -31896
rect 8589 -31902 8961 -31896
rect 9589 -31902 9961 -31896
rect 10589 -31902 10961 -31896
rect 11589 -31902 11961 -31896
rect 12589 -31902 12961 -31896
rect 13589 -31902 13961 -31896
rect 14589 -31902 14961 -31896
rect 15589 -31902 15961 -31896
rect 16589 -31902 16961 -31896
rect 17589 -31902 17961 -31896
rect 18589 -31902 18961 -31896
rect 19589 -31902 19961 -31896
rect 20589 -31902 20961 -31896
rect 21589 -31902 21961 -31896
rect 22589 -31902 22961 -31896
rect 23589 -31902 23961 -31896
rect 24589 -31902 24961 -31896
rect 25589 -31902 25961 -31896
rect 26589 -31902 26961 -31896
rect 27589 -31902 27961 -31896
rect 28589 -31902 28961 -31896
rect 29589 -31902 29961 -31896
rect 30589 -31902 30961 -31896
rect 31589 -31902 31961 -31896
rect 32589 -31902 32961 -31896
rect 33589 -31902 33961 -31896
rect 8589 -32198 8627 -31902
rect 8923 -32198 8961 -31902
rect 9589 -32198 9627 -31902
rect 9923 -32198 9961 -31902
rect 10589 -32198 10627 -31902
rect 10923 -32198 10961 -31902
rect 11589 -32198 11627 -31902
rect 11923 -32198 11961 -31902
rect 12589 -32198 12627 -31902
rect 12923 -32198 12961 -31902
rect 13589 -32198 13627 -31902
rect 13923 -32198 13961 -31902
rect 14589 -32198 14627 -31902
rect 14923 -32198 14961 -31902
rect 15589 -32198 15627 -31902
rect 15923 -32198 15961 -31902
rect 16589 -32198 16627 -31902
rect 16923 -32198 16961 -31902
rect 17589 -32198 17627 -31902
rect 17923 -32198 17961 -31902
rect 18589 -32198 18627 -31902
rect 18923 -32198 18961 -31902
rect 19589 -32198 19627 -31902
rect 19923 -32198 19961 -31902
rect 20589 -32198 20627 -31902
rect 20923 -32198 20961 -31902
rect 21589 -32198 21627 -31902
rect 21923 -32198 21961 -31902
rect 22589 -32198 22627 -31902
rect 22923 -32198 22961 -31902
rect 23589 -32198 23627 -31902
rect 23923 -32198 23961 -31902
rect 24589 -32198 24627 -31902
rect 24923 -32198 24961 -31902
rect 25589 -32198 25627 -31902
rect 25923 -32198 25961 -31902
rect 26589 -32198 26627 -31902
rect 26923 -32198 26961 -31902
rect 27589 -32198 27627 -31902
rect 27923 -32198 27961 -31902
rect 28589 -32198 28627 -31902
rect 28923 -32198 28961 -31902
rect 29589 -32198 29627 -31902
rect 29923 -32198 29961 -31902
rect 30589 -32198 30627 -31902
rect 30923 -32198 30961 -31902
rect 31589 -32198 31627 -31902
rect 31923 -32198 31961 -31902
rect 32589 -32198 32627 -31902
rect 32923 -32198 32961 -31902
rect 33589 -32198 33627 -31902
rect 33923 -32198 33961 -31902
rect 8589 -32204 8961 -32198
rect 9589 -32204 9961 -32198
rect 10589 -32204 10961 -32198
rect 11589 -32204 11961 -32198
rect 12589 -32204 12961 -32198
rect 13589 -32204 13961 -32198
rect 14589 -32204 14961 -32198
rect 15589 -32204 15961 -32198
rect 16589 -32204 16961 -32198
rect 17589 -32204 17961 -32198
rect 18589 -32204 18961 -32198
rect 19589 -32204 19961 -32198
rect 20589 -32204 20961 -32198
rect 21589 -32204 21961 -32198
rect 22589 -32204 22961 -32198
rect 23589 -32204 23961 -32198
rect 24589 -32204 24961 -32198
rect 25589 -32204 25961 -32198
rect 26589 -32204 26961 -32198
rect 27589 -32204 27961 -32198
rect 28589 -32204 28961 -32198
rect 29589 -32204 29961 -32198
rect 30589 -32204 30961 -32198
rect 31589 -32204 31961 -32198
rect 32589 -32204 32961 -32198
rect 33589 -32204 33961 -32198
rect 34269 -32204 34275 -31896
rect 8275 -32210 34275 -32204
rect -74485 -32236 -74165 -32210
rect -74485 -32864 -74479 -32236
rect -74171 -32864 -74165 -32236
rect -74485 -32890 -74165 -32864
rect -73485 -32236 -73165 -32210
rect -73485 -32864 -73479 -32236
rect -73171 -32864 -73165 -32236
rect -73485 -32890 -73165 -32864
rect -72485 -32236 -72165 -32210
rect -72485 -32864 -72479 -32236
rect -72171 -32864 -72165 -32236
rect -72485 -32890 -72165 -32864
rect -71485 -32236 -71165 -32210
rect -71485 -32864 -71479 -32236
rect -71171 -32864 -71165 -32236
rect -71485 -32890 -71165 -32864
rect -70485 -32236 -70165 -32210
rect -70485 -32864 -70479 -32236
rect -70171 -32864 -70165 -32236
rect -70485 -32890 -70165 -32864
rect -69485 -32236 -69165 -32210
rect -69485 -32864 -69479 -32236
rect -69171 -32864 -69165 -32236
rect -69485 -32890 -69165 -32864
rect -68485 -32236 -68165 -32210
rect -68485 -32864 -68479 -32236
rect -68171 -32864 -68165 -32236
rect -68485 -32890 -68165 -32864
rect -67485 -32236 -67165 -32210
rect -67485 -32864 -67479 -32236
rect -67171 -32864 -67165 -32236
rect -67485 -32890 -67165 -32864
rect -66485 -32236 -66165 -32210
rect -66485 -32864 -66479 -32236
rect -66171 -32864 -66165 -32236
rect -66485 -32890 -66165 -32864
rect -65485 -32236 -65165 -32210
rect -65485 -32864 -65479 -32236
rect -65171 -32864 -65165 -32236
rect -65485 -32890 -65165 -32864
rect -64485 -32236 -64165 -32210
rect -64485 -32864 -64479 -32236
rect -64171 -32864 -64165 -32236
rect -64485 -32890 -64165 -32864
rect -63485 -32236 -63165 -32210
rect -63485 -32864 -63479 -32236
rect -63171 -32864 -63165 -32236
rect -63485 -32890 -63165 -32864
rect -62485 -32236 -62165 -32210
rect -62485 -32864 -62479 -32236
rect -62171 -32864 -62165 -32236
rect -62485 -32890 -62165 -32864
rect -61485 -32236 -61165 -32210
rect -61485 -32864 -61479 -32236
rect -61171 -32864 -61165 -32236
rect -61485 -32890 -61165 -32864
rect -60485 -32236 -60165 -32210
rect -60485 -32864 -60479 -32236
rect -60171 -32864 -60165 -32236
rect -60485 -32890 -60165 -32864
rect -59485 -32236 -59165 -32210
rect -59485 -32864 -59479 -32236
rect -59171 -32864 -59165 -32236
rect -59485 -32890 -59165 -32864
rect -58485 -32236 -58165 -32210
rect -58485 -32864 -58479 -32236
rect -58171 -32864 -58165 -32236
rect -58485 -32890 -58165 -32864
rect -57485 -32236 -57165 -32210
rect -57485 -32864 -57479 -32236
rect -57171 -32864 -57165 -32236
rect -57485 -32890 -57165 -32864
rect -56485 -32236 -56165 -32210
rect -56485 -32864 -56479 -32236
rect -56171 -32864 -56165 -32236
rect -56485 -32890 -56165 -32864
rect -55485 -32236 -55165 -32210
rect -55485 -32864 -55479 -32236
rect -55171 -32864 -55165 -32236
rect -55485 -32890 -55165 -32864
rect -54485 -32236 -54165 -32210
rect -54485 -32864 -54479 -32236
rect -54171 -32864 -54165 -32236
rect -54485 -32890 -54165 -32864
rect -53485 -32236 -53165 -32210
rect -53485 -32864 -53479 -32236
rect -53171 -32864 -53165 -32236
rect -53485 -32890 -53165 -32864
rect -52485 -32236 -52165 -32210
rect -52485 -32864 -52479 -32236
rect -52171 -32864 -52165 -32236
rect -52485 -32890 -52165 -32864
rect -51485 -32236 -51165 -32210
rect -51485 -32864 -51479 -32236
rect -51171 -32864 -51165 -32236
rect -51485 -32890 -51165 -32864
rect -50485 -32236 -50165 -32210
rect -50485 -32864 -50479 -32236
rect -50171 -32864 -50165 -32236
rect -50485 -32890 -50165 -32864
rect -49485 -32236 -49165 -32210
rect -49485 -32864 -49479 -32236
rect -49171 -32864 -49165 -32236
rect 8615 -32236 8935 -32210
rect -49485 -32890 -49165 -32864
rect -46275 -32602 -36275 -32550
rect -46275 -32604 -46228 -32602
rect -36332 -32604 -36275 -32602
rect -74825 -32896 -48825 -32890
rect -74825 -33204 -74819 -32896
rect -74511 -32902 -74139 -32896
rect -73511 -32902 -73139 -32896
rect -72511 -32902 -72139 -32896
rect -71511 -32902 -71139 -32896
rect -70511 -32902 -70139 -32896
rect -69511 -32902 -69139 -32896
rect -68511 -32902 -68139 -32896
rect -67511 -32902 -67139 -32896
rect -66511 -32902 -66139 -32896
rect -65511 -32902 -65139 -32896
rect -64511 -32902 -64139 -32896
rect -63511 -32902 -63139 -32896
rect -62511 -32902 -62139 -32896
rect -61511 -32902 -61139 -32896
rect -60511 -32902 -60139 -32896
rect -59511 -32902 -59139 -32896
rect -58511 -32902 -58139 -32896
rect -57511 -32902 -57139 -32896
rect -56511 -32902 -56139 -32896
rect -55511 -32902 -55139 -32896
rect -54511 -32902 -54139 -32896
rect -53511 -32902 -53139 -32896
rect -52511 -32902 -52139 -32896
rect -51511 -32902 -51139 -32896
rect -50511 -32902 -50139 -32896
rect -49511 -32902 -49139 -32896
rect -74511 -33198 -74473 -32902
rect -74177 -33198 -74139 -32902
rect -73511 -33198 -73473 -32902
rect -73177 -33198 -73139 -32902
rect -72511 -33198 -72473 -32902
rect -72177 -33198 -72139 -32902
rect -71511 -33198 -71473 -32902
rect -71177 -33198 -71139 -32902
rect -70511 -33198 -70473 -32902
rect -70177 -33198 -70139 -32902
rect -69511 -33198 -69473 -32902
rect -69177 -33198 -69139 -32902
rect -68511 -33198 -68473 -32902
rect -68177 -33198 -68139 -32902
rect -67511 -33198 -67473 -32902
rect -67177 -33198 -67139 -32902
rect -66511 -33198 -66473 -32902
rect -66177 -33198 -66139 -32902
rect -65511 -33198 -65473 -32902
rect -65177 -33198 -65139 -32902
rect -64511 -33198 -64473 -32902
rect -64177 -33198 -64139 -32902
rect -63511 -33198 -63473 -32902
rect -63177 -33198 -63139 -32902
rect -62511 -33198 -62473 -32902
rect -62177 -33198 -62139 -32902
rect -61511 -33198 -61473 -32902
rect -61177 -33198 -61139 -32902
rect -60511 -33198 -60473 -32902
rect -60177 -33198 -60139 -32902
rect -59511 -33198 -59473 -32902
rect -59177 -33198 -59139 -32902
rect -58511 -33198 -58473 -32902
rect -58177 -33198 -58139 -32902
rect -57511 -33198 -57473 -32902
rect -57177 -33198 -57139 -32902
rect -56511 -33198 -56473 -32902
rect -56177 -33198 -56139 -32902
rect -55511 -33198 -55473 -32902
rect -55177 -33198 -55139 -32902
rect -54511 -33198 -54473 -32902
rect -54177 -33198 -54139 -32902
rect -53511 -33198 -53473 -32902
rect -53177 -33198 -53139 -32902
rect -52511 -33198 -52473 -32902
rect -52177 -33198 -52139 -32902
rect -51511 -33198 -51473 -32902
rect -51177 -33198 -51139 -32902
rect -50511 -33198 -50473 -32902
rect -50177 -33198 -50139 -32902
rect -49511 -33198 -49473 -32902
rect -49177 -33198 -49139 -32902
rect -74511 -33204 -74139 -33198
rect -73511 -33204 -73139 -33198
rect -72511 -33204 -72139 -33198
rect -71511 -33204 -71139 -33198
rect -70511 -33204 -70139 -33198
rect -69511 -33204 -69139 -33198
rect -68511 -33204 -68139 -33198
rect -67511 -33204 -67139 -33198
rect -66511 -33204 -66139 -33198
rect -65511 -33204 -65139 -33198
rect -64511 -33204 -64139 -33198
rect -63511 -33204 -63139 -33198
rect -62511 -33204 -62139 -33198
rect -61511 -33204 -61139 -33198
rect -60511 -33204 -60139 -33198
rect -59511 -33204 -59139 -33198
rect -58511 -33204 -58139 -33198
rect -57511 -33204 -57139 -33198
rect -56511 -33204 -56139 -33198
rect -55511 -33204 -55139 -33198
rect -54511 -33204 -54139 -33198
rect -53511 -33204 -53139 -33198
rect -52511 -33204 -52139 -33198
rect -51511 -33204 -51139 -33198
rect -50511 -33204 -50139 -33198
rect -49511 -33204 -49139 -33198
rect -48831 -33204 -48825 -32896
rect -74825 -33210 -48825 -33204
rect -74485 -33236 -74165 -33210
rect -74485 -33864 -74479 -33236
rect -74171 -33864 -74165 -33236
rect -74485 -33890 -74165 -33864
rect -73485 -33236 -73165 -33210
rect -73485 -33864 -73479 -33236
rect -73171 -33864 -73165 -33236
rect -73485 -33890 -73165 -33864
rect -72485 -33236 -72165 -33210
rect -72485 -33864 -72479 -33236
rect -72171 -33864 -72165 -33236
rect -72485 -33890 -72165 -33864
rect -71485 -33236 -71165 -33210
rect -71485 -33864 -71479 -33236
rect -71171 -33864 -71165 -33236
rect -71485 -33890 -71165 -33864
rect -70485 -33236 -70165 -33210
rect -70485 -33864 -70479 -33236
rect -70171 -33864 -70165 -33236
rect -70485 -33890 -70165 -33864
rect -69485 -33236 -69165 -33210
rect -69485 -33864 -69479 -33236
rect -69171 -33864 -69165 -33236
rect -69485 -33890 -69165 -33864
rect -68485 -33236 -68165 -33210
rect -68485 -33864 -68479 -33236
rect -68171 -33864 -68165 -33236
rect -68485 -33890 -68165 -33864
rect -67485 -33236 -67165 -33210
rect -67485 -33864 -67479 -33236
rect -67171 -33864 -67165 -33236
rect -67485 -33890 -67165 -33864
rect -66485 -33236 -66165 -33210
rect -66485 -33864 -66479 -33236
rect -66171 -33864 -66165 -33236
rect -66485 -33890 -66165 -33864
rect -65485 -33236 -65165 -33210
rect -65485 -33864 -65479 -33236
rect -65171 -33864 -65165 -33236
rect -65485 -33890 -65165 -33864
rect -64485 -33236 -64165 -33210
rect -64485 -33864 -64479 -33236
rect -64171 -33864 -64165 -33236
rect -64485 -33890 -64165 -33864
rect -63485 -33236 -63165 -33210
rect -63485 -33864 -63479 -33236
rect -63171 -33864 -63165 -33236
rect -63485 -33890 -63165 -33864
rect -62485 -33236 -62165 -33210
rect -62485 -33864 -62479 -33236
rect -62171 -33864 -62165 -33236
rect -62485 -33890 -62165 -33864
rect -61485 -33236 -61165 -33210
rect -61485 -33864 -61479 -33236
rect -61171 -33864 -61165 -33236
rect -61485 -33890 -61165 -33864
rect -60485 -33236 -60165 -33210
rect -60485 -33864 -60479 -33236
rect -60171 -33864 -60165 -33236
rect -60485 -33890 -60165 -33864
rect -59485 -33236 -59165 -33210
rect -59485 -33864 -59479 -33236
rect -59171 -33864 -59165 -33236
rect -59485 -33890 -59165 -33864
rect -58485 -33236 -58165 -33210
rect -58485 -33864 -58479 -33236
rect -58171 -33864 -58165 -33236
rect -58485 -33890 -58165 -33864
rect -57485 -33236 -57165 -33210
rect -57485 -33864 -57479 -33236
rect -57171 -33864 -57165 -33236
rect -57485 -33890 -57165 -33864
rect -56485 -33236 -56165 -33210
rect -56485 -33864 -56479 -33236
rect -56171 -33864 -56165 -33236
rect -56485 -33890 -56165 -33864
rect -55485 -33236 -55165 -33210
rect -55485 -33864 -55479 -33236
rect -55171 -33864 -55165 -33236
rect -55485 -33890 -55165 -33864
rect -54485 -33236 -54165 -33210
rect -54485 -33864 -54479 -33236
rect -54171 -33864 -54165 -33236
rect -54485 -33890 -54165 -33864
rect -53485 -33236 -53165 -33210
rect -53485 -33864 -53479 -33236
rect -53171 -33864 -53165 -33236
rect -53485 -33890 -53165 -33864
rect -52485 -33236 -52165 -33210
rect -52485 -33864 -52479 -33236
rect -52171 -33864 -52165 -33236
rect -52485 -33890 -52165 -33864
rect -51485 -33236 -51165 -33210
rect -51485 -33864 -51479 -33236
rect -51171 -33864 -51165 -33236
rect -51485 -33890 -51165 -33864
rect -50485 -33236 -50165 -33210
rect -50485 -33864 -50479 -33236
rect -50171 -33864 -50165 -33236
rect -50485 -33890 -50165 -33864
rect -49485 -33236 -49165 -33210
rect -49485 -33864 -49479 -33236
rect -49171 -33864 -49165 -33236
rect -49485 -33890 -49165 -33864
rect -74825 -33896 -48825 -33890
rect -74825 -34204 -74819 -33896
rect -74511 -33902 -74139 -33896
rect -73511 -33902 -73139 -33896
rect -72511 -33902 -72139 -33896
rect -71511 -33902 -71139 -33896
rect -70511 -33902 -70139 -33896
rect -69511 -33902 -69139 -33896
rect -68511 -33902 -68139 -33896
rect -67511 -33902 -67139 -33896
rect -66511 -33902 -66139 -33896
rect -65511 -33902 -65139 -33896
rect -64511 -33902 -64139 -33896
rect -63511 -33902 -63139 -33896
rect -62511 -33902 -62139 -33896
rect -61511 -33902 -61139 -33896
rect -60511 -33902 -60139 -33896
rect -59511 -33902 -59139 -33896
rect -58511 -33902 -58139 -33896
rect -57511 -33902 -57139 -33896
rect -56511 -33902 -56139 -33896
rect -55511 -33902 -55139 -33896
rect -54511 -33902 -54139 -33896
rect -53511 -33902 -53139 -33896
rect -52511 -33902 -52139 -33896
rect -51511 -33902 -51139 -33896
rect -50511 -33902 -50139 -33896
rect -49511 -33902 -49139 -33896
rect -74511 -34198 -74473 -33902
rect -74177 -34198 -74139 -33902
rect -73511 -34198 -73473 -33902
rect -73177 -34198 -73139 -33902
rect -72511 -34198 -72473 -33902
rect -72177 -34198 -72139 -33902
rect -71511 -34198 -71473 -33902
rect -71177 -34198 -71139 -33902
rect -70511 -34198 -70473 -33902
rect -70177 -34198 -70139 -33902
rect -69511 -34198 -69473 -33902
rect -69177 -34198 -69139 -33902
rect -68511 -34198 -68473 -33902
rect -68177 -34198 -68139 -33902
rect -67511 -34198 -67473 -33902
rect -67177 -34198 -67139 -33902
rect -66511 -34198 -66473 -33902
rect -66177 -34198 -66139 -33902
rect -65511 -34198 -65473 -33902
rect -65177 -34198 -65139 -33902
rect -64511 -34198 -64473 -33902
rect -64177 -34198 -64139 -33902
rect -63511 -34198 -63473 -33902
rect -63177 -34198 -63139 -33902
rect -62511 -34198 -62473 -33902
rect -62177 -34198 -62139 -33902
rect -61511 -34198 -61473 -33902
rect -61177 -34198 -61139 -33902
rect -60511 -34198 -60473 -33902
rect -60177 -34198 -60139 -33902
rect -59511 -34198 -59473 -33902
rect -59177 -34198 -59139 -33902
rect -58511 -34198 -58473 -33902
rect -58177 -34198 -58139 -33902
rect -57511 -34198 -57473 -33902
rect -57177 -34198 -57139 -33902
rect -56511 -34198 -56473 -33902
rect -56177 -34198 -56139 -33902
rect -55511 -34198 -55473 -33902
rect -55177 -34198 -55139 -33902
rect -54511 -34198 -54473 -33902
rect -54177 -34198 -54139 -33902
rect -53511 -34198 -53473 -33902
rect -53177 -34198 -53139 -33902
rect -52511 -34198 -52473 -33902
rect -52177 -34198 -52139 -33902
rect -51511 -34198 -51473 -33902
rect -51177 -34198 -51139 -33902
rect -50511 -34198 -50473 -33902
rect -50177 -34198 -50139 -33902
rect -49511 -34198 -49473 -33902
rect -49177 -34198 -49139 -33902
rect -74511 -34204 -74139 -34198
rect -73511 -34204 -73139 -34198
rect -72511 -34204 -72139 -34198
rect -71511 -34204 -71139 -34198
rect -70511 -34204 -70139 -34198
rect -69511 -34204 -69139 -34198
rect -68511 -34204 -68139 -34198
rect -67511 -34204 -67139 -34198
rect -66511 -34204 -66139 -34198
rect -65511 -34204 -65139 -34198
rect -64511 -34204 -64139 -34198
rect -63511 -34204 -63139 -34198
rect -62511 -34204 -62139 -34198
rect -61511 -34204 -61139 -34198
rect -60511 -34204 -60139 -34198
rect -59511 -34204 -59139 -34198
rect -58511 -34204 -58139 -34198
rect -57511 -34204 -57139 -34198
rect -56511 -34204 -56139 -34198
rect -55511 -34204 -55139 -34198
rect -54511 -34204 -54139 -34198
rect -53511 -34204 -53139 -34198
rect -52511 -34204 -52139 -34198
rect -51511 -34204 -51139 -34198
rect -50511 -34204 -50139 -34198
rect -49511 -34204 -49139 -34198
rect -48831 -34204 -48825 -33896
rect -74825 -34210 -48825 -34204
rect -74485 -34236 -74165 -34210
rect -74485 -34864 -74479 -34236
rect -74171 -34864 -74165 -34236
rect -74485 -34890 -74165 -34864
rect -73485 -34236 -73165 -34210
rect -73485 -34864 -73479 -34236
rect -73171 -34864 -73165 -34236
rect -73485 -34890 -73165 -34864
rect -72485 -34236 -72165 -34210
rect -72485 -34864 -72479 -34236
rect -72171 -34864 -72165 -34236
rect -72485 -34890 -72165 -34864
rect -71485 -34236 -71165 -34210
rect -71485 -34864 -71479 -34236
rect -71171 -34864 -71165 -34236
rect -71485 -34890 -71165 -34864
rect -70485 -34236 -70165 -34210
rect -70485 -34864 -70479 -34236
rect -70171 -34864 -70165 -34236
rect -70485 -34890 -70165 -34864
rect -69485 -34236 -69165 -34210
rect -69485 -34864 -69479 -34236
rect -69171 -34864 -69165 -34236
rect -69485 -34890 -69165 -34864
rect -68485 -34236 -68165 -34210
rect -68485 -34864 -68479 -34236
rect -68171 -34864 -68165 -34236
rect -68485 -34890 -68165 -34864
rect -67485 -34236 -67165 -34210
rect -67485 -34864 -67479 -34236
rect -67171 -34864 -67165 -34236
rect -67485 -34890 -67165 -34864
rect -66485 -34236 -66165 -34210
rect -66485 -34864 -66479 -34236
rect -66171 -34864 -66165 -34236
rect -66485 -34890 -66165 -34864
rect -65485 -34236 -65165 -34210
rect -65485 -34864 -65479 -34236
rect -65171 -34864 -65165 -34236
rect -65485 -34890 -65165 -34864
rect -64485 -34236 -64165 -34210
rect -64485 -34864 -64479 -34236
rect -64171 -34864 -64165 -34236
rect -64485 -34890 -64165 -34864
rect -63485 -34236 -63165 -34210
rect -63485 -34864 -63479 -34236
rect -63171 -34864 -63165 -34236
rect -63485 -34890 -63165 -34864
rect -62485 -34236 -62165 -34210
rect -62485 -34864 -62479 -34236
rect -62171 -34864 -62165 -34236
rect -62485 -34890 -62165 -34864
rect -61485 -34236 -61165 -34210
rect -61485 -34864 -61479 -34236
rect -61171 -34864 -61165 -34236
rect -61485 -34890 -61165 -34864
rect -60485 -34236 -60165 -34210
rect -60485 -34864 -60479 -34236
rect -60171 -34864 -60165 -34236
rect -60485 -34890 -60165 -34864
rect -59485 -34236 -59165 -34210
rect -59485 -34864 -59479 -34236
rect -59171 -34864 -59165 -34236
rect -59485 -34890 -59165 -34864
rect -58485 -34236 -58165 -34210
rect -58485 -34864 -58479 -34236
rect -58171 -34864 -58165 -34236
rect -58485 -34890 -58165 -34864
rect -57485 -34236 -57165 -34210
rect -57485 -34864 -57479 -34236
rect -57171 -34864 -57165 -34236
rect -57485 -34890 -57165 -34864
rect -56485 -34236 -56165 -34210
rect -56485 -34864 -56479 -34236
rect -56171 -34864 -56165 -34236
rect -56485 -34890 -56165 -34864
rect -55485 -34236 -55165 -34210
rect -55485 -34864 -55479 -34236
rect -55171 -34864 -55165 -34236
rect -55485 -34890 -55165 -34864
rect -54485 -34236 -54165 -34210
rect -54485 -34864 -54479 -34236
rect -54171 -34864 -54165 -34236
rect -54485 -34890 -54165 -34864
rect -53485 -34236 -53165 -34210
rect -53485 -34864 -53479 -34236
rect -53171 -34864 -53165 -34236
rect -53485 -34890 -53165 -34864
rect -52485 -34236 -52165 -34210
rect -52485 -34864 -52479 -34236
rect -52171 -34864 -52165 -34236
rect -52485 -34890 -52165 -34864
rect -51485 -34236 -51165 -34210
rect -51485 -34864 -51479 -34236
rect -51171 -34864 -51165 -34236
rect -51485 -34890 -51165 -34864
rect -50485 -34236 -50165 -34210
rect -50485 -34864 -50479 -34236
rect -50171 -34864 -50165 -34236
rect -50485 -34890 -50165 -34864
rect -49485 -34236 -49165 -34210
rect -49485 -34864 -49479 -34236
rect -49171 -34864 -49165 -34236
rect -49485 -34890 -49165 -34864
rect -74825 -34896 -48825 -34890
rect -74825 -35204 -74819 -34896
rect -74511 -34902 -74139 -34896
rect -73511 -34902 -73139 -34896
rect -72511 -34902 -72139 -34896
rect -71511 -34902 -71139 -34896
rect -70511 -34902 -70139 -34896
rect -69511 -34902 -69139 -34896
rect -68511 -34902 -68139 -34896
rect -67511 -34902 -67139 -34896
rect -66511 -34902 -66139 -34896
rect -65511 -34902 -65139 -34896
rect -64511 -34902 -64139 -34896
rect -63511 -34902 -63139 -34896
rect -62511 -34902 -62139 -34896
rect -61511 -34902 -61139 -34896
rect -60511 -34902 -60139 -34896
rect -59511 -34902 -59139 -34896
rect -58511 -34902 -58139 -34896
rect -57511 -34902 -57139 -34896
rect -56511 -34902 -56139 -34896
rect -55511 -34902 -55139 -34896
rect -54511 -34902 -54139 -34896
rect -53511 -34902 -53139 -34896
rect -52511 -34902 -52139 -34896
rect -51511 -34902 -51139 -34896
rect -50511 -34902 -50139 -34896
rect -49511 -34902 -49139 -34896
rect -74511 -35198 -74473 -34902
rect -74177 -35198 -74139 -34902
rect -73511 -35198 -73473 -34902
rect -73177 -35198 -73139 -34902
rect -72511 -35198 -72473 -34902
rect -72177 -35198 -72139 -34902
rect -71511 -35198 -71473 -34902
rect -71177 -35198 -71139 -34902
rect -70511 -35198 -70473 -34902
rect -70177 -35198 -70139 -34902
rect -69511 -35198 -69473 -34902
rect -69177 -35198 -69139 -34902
rect -68511 -35198 -68473 -34902
rect -68177 -35198 -68139 -34902
rect -67511 -35198 -67473 -34902
rect -67177 -35198 -67139 -34902
rect -66511 -35198 -66473 -34902
rect -66177 -35198 -66139 -34902
rect -65511 -35198 -65473 -34902
rect -65177 -35198 -65139 -34902
rect -64511 -35198 -64473 -34902
rect -64177 -35198 -64139 -34902
rect -63511 -35198 -63473 -34902
rect -63177 -35198 -63139 -34902
rect -62511 -35198 -62473 -34902
rect -62177 -35198 -62139 -34902
rect -61511 -35198 -61473 -34902
rect -61177 -35198 -61139 -34902
rect -60511 -35198 -60473 -34902
rect -60177 -35198 -60139 -34902
rect -59511 -35198 -59473 -34902
rect -59177 -35198 -59139 -34902
rect -58511 -35198 -58473 -34902
rect -58177 -35198 -58139 -34902
rect -57511 -35198 -57473 -34902
rect -57177 -35198 -57139 -34902
rect -56511 -35198 -56473 -34902
rect -56177 -35198 -56139 -34902
rect -55511 -35198 -55473 -34902
rect -55177 -35198 -55139 -34902
rect -54511 -35198 -54473 -34902
rect -54177 -35198 -54139 -34902
rect -53511 -35198 -53473 -34902
rect -53177 -35198 -53139 -34902
rect -52511 -35198 -52473 -34902
rect -52177 -35198 -52139 -34902
rect -51511 -35198 -51473 -34902
rect -51177 -35198 -51139 -34902
rect -50511 -35198 -50473 -34902
rect -50177 -35198 -50139 -34902
rect -49511 -35198 -49473 -34902
rect -49177 -35198 -49139 -34902
rect -74511 -35204 -74139 -35198
rect -73511 -35204 -73139 -35198
rect -72511 -35204 -72139 -35198
rect -71511 -35204 -71139 -35198
rect -70511 -35204 -70139 -35198
rect -69511 -35204 -69139 -35198
rect -68511 -35204 -68139 -35198
rect -67511 -35204 -67139 -35198
rect -66511 -35204 -66139 -35198
rect -65511 -35204 -65139 -35198
rect -64511 -35204 -64139 -35198
rect -63511 -35204 -63139 -35198
rect -62511 -35204 -62139 -35198
rect -61511 -35204 -61139 -35198
rect -60511 -35204 -60139 -35198
rect -59511 -35204 -59139 -35198
rect -58511 -35204 -58139 -35198
rect -57511 -35204 -57139 -35198
rect -56511 -35204 -56139 -35198
rect -55511 -35204 -55139 -35198
rect -54511 -35204 -54139 -35198
rect -53511 -35204 -53139 -35198
rect -52511 -35204 -52139 -35198
rect -51511 -35204 -51139 -35198
rect -50511 -35204 -50139 -35198
rect -49511 -35204 -49139 -35198
rect -48831 -35204 -48825 -34896
rect -74825 -35210 -48825 -35204
rect -74485 -35236 -74165 -35210
rect -74485 -35864 -74479 -35236
rect -74171 -35864 -74165 -35236
rect -74485 -35890 -74165 -35864
rect -73485 -35236 -73165 -35210
rect -73485 -35864 -73479 -35236
rect -73171 -35864 -73165 -35236
rect -73485 -35890 -73165 -35864
rect -72485 -35236 -72165 -35210
rect -72485 -35864 -72479 -35236
rect -72171 -35864 -72165 -35236
rect -72485 -35890 -72165 -35864
rect -71485 -35236 -71165 -35210
rect -71485 -35864 -71479 -35236
rect -71171 -35864 -71165 -35236
rect -71485 -35890 -71165 -35864
rect -70485 -35236 -70165 -35210
rect -70485 -35864 -70479 -35236
rect -70171 -35864 -70165 -35236
rect -70485 -35890 -70165 -35864
rect -69485 -35236 -69165 -35210
rect -69485 -35864 -69479 -35236
rect -69171 -35864 -69165 -35236
rect -69485 -35890 -69165 -35864
rect -68485 -35236 -68165 -35210
rect -68485 -35864 -68479 -35236
rect -68171 -35864 -68165 -35236
rect -68485 -35890 -68165 -35864
rect -67485 -35236 -67165 -35210
rect -67485 -35864 -67479 -35236
rect -67171 -35864 -67165 -35236
rect -67485 -35890 -67165 -35864
rect -66485 -35236 -66165 -35210
rect -66485 -35864 -66479 -35236
rect -66171 -35864 -66165 -35236
rect -66485 -35890 -66165 -35864
rect -65485 -35236 -65165 -35210
rect -65485 -35864 -65479 -35236
rect -65171 -35864 -65165 -35236
rect -65485 -35890 -65165 -35864
rect -64485 -35236 -64165 -35210
rect -64485 -35864 -64479 -35236
rect -64171 -35864 -64165 -35236
rect -64485 -35890 -64165 -35864
rect -63485 -35236 -63165 -35210
rect -63485 -35864 -63479 -35236
rect -63171 -35864 -63165 -35236
rect -63485 -35890 -63165 -35864
rect -62485 -35236 -62165 -35210
rect -62485 -35864 -62479 -35236
rect -62171 -35864 -62165 -35236
rect -62485 -35890 -62165 -35864
rect -61485 -35236 -61165 -35210
rect -61485 -35864 -61479 -35236
rect -61171 -35864 -61165 -35236
rect -61485 -35890 -61165 -35864
rect -60485 -35236 -60165 -35210
rect -60485 -35864 -60479 -35236
rect -60171 -35864 -60165 -35236
rect -60485 -35890 -60165 -35864
rect -59485 -35236 -59165 -35210
rect -59485 -35864 -59479 -35236
rect -59171 -35864 -59165 -35236
rect -59485 -35890 -59165 -35864
rect -58485 -35236 -58165 -35210
rect -58485 -35864 -58479 -35236
rect -58171 -35864 -58165 -35236
rect -58485 -35890 -58165 -35864
rect -57485 -35236 -57165 -35210
rect -57485 -35864 -57479 -35236
rect -57171 -35864 -57165 -35236
rect -57485 -35890 -57165 -35864
rect -56485 -35236 -56165 -35210
rect -56485 -35864 -56479 -35236
rect -56171 -35864 -56165 -35236
rect -56485 -35890 -56165 -35864
rect -55485 -35236 -55165 -35210
rect -55485 -35864 -55479 -35236
rect -55171 -35864 -55165 -35236
rect -55485 -35890 -55165 -35864
rect -54485 -35236 -54165 -35210
rect -54485 -35864 -54479 -35236
rect -54171 -35864 -54165 -35236
rect -54485 -35890 -54165 -35864
rect -53485 -35236 -53165 -35210
rect -53485 -35864 -53479 -35236
rect -53171 -35864 -53165 -35236
rect -53485 -35890 -53165 -35864
rect -52485 -35236 -52165 -35210
rect -52485 -35864 -52479 -35236
rect -52171 -35864 -52165 -35236
rect -52485 -35890 -52165 -35864
rect -51485 -35236 -51165 -35210
rect -51485 -35864 -51479 -35236
rect -51171 -35864 -51165 -35236
rect -51485 -35890 -51165 -35864
rect -50485 -35236 -50165 -35210
rect -50485 -35864 -50479 -35236
rect -50171 -35864 -50165 -35236
rect -50485 -35890 -50165 -35864
rect -49485 -35236 -49165 -35210
rect -49485 -35864 -49479 -35236
rect -49171 -35864 -49165 -35236
rect -49485 -35890 -49165 -35864
rect -74825 -35896 -48825 -35890
rect -74825 -36204 -74819 -35896
rect -74511 -35902 -74139 -35896
rect -73511 -35902 -73139 -35896
rect -72511 -35902 -72139 -35896
rect -71511 -35902 -71139 -35896
rect -70511 -35902 -70139 -35896
rect -69511 -35902 -69139 -35896
rect -68511 -35902 -68139 -35896
rect -67511 -35902 -67139 -35896
rect -66511 -35902 -66139 -35896
rect -65511 -35902 -65139 -35896
rect -64511 -35902 -64139 -35896
rect -63511 -35902 -63139 -35896
rect -62511 -35902 -62139 -35896
rect -61511 -35902 -61139 -35896
rect -60511 -35902 -60139 -35896
rect -59511 -35902 -59139 -35896
rect -58511 -35902 -58139 -35896
rect -57511 -35902 -57139 -35896
rect -56511 -35902 -56139 -35896
rect -55511 -35902 -55139 -35896
rect -54511 -35902 -54139 -35896
rect -53511 -35902 -53139 -35896
rect -52511 -35902 -52139 -35896
rect -51511 -35902 -51139 -35896
rect -50511 -35902 -50139 -35896
rect -49511 -35902 -49139 -35896
rect -74511 -36198 -74473 -35902
rect -74177 -36198 -74139 -35902
rect -73511 -36198 -73473 -35902
rect -73177 -36198 -73139 -35902
rect -72511 -36198 -72473 -35902
rect -72177 -36198 -72139 -35902
rect -71511 -36198 -71473 -35902
rect -71177 -36198 -71139 -35902
rect -70511 -36198 -70473 -35902
rect -70177 -36198 -70139 -35902
rect -69511 -36198 -69473 -35902
rect -69177 -36198 -69139 -35902
rect -68511 -36198 -68473 -35902
rect -68177 -36198 -68139 -35902
rect -67511 -36198 -67473 -35902
rect -67177 -36198 -67139 -35902
rect -66511 -36198 -66473 -35902
rect -66177 -36198 -66139 -35902
rect -65511 -36198 -65473 -35902
rect -65177 -36198 -65139 -35902
rect -64511 -36198 -64473 -35902
rect -64177 -36198 -64139 -35902
rect -63511 -36198 -63473 -35902
rect -63177 -36198 -63139 -35902
rect -62511 -36198 -62473 -35902
rect -62177 -36198 -62139 -35902
rect -61511 -36198 -61473 -35902
rect -61177 -36198 -61139 -35902
rect -60511 -36198 -60473 -35902
rect -60177 -36198 -60139 -35902
rect -59511 -36198 -59473 -35902
rect -59177 -36198 -59139 -35902
rect -58511 -36198 -58473 -35902
rect -58177 -36198 -58139 -35902
rect -57511 -36198 -57473 -35902
rect -57177 -36198 -57139 -35902
rect -56511 -36198 -56473 -35902
rect -56177 -36198 -56139 -35902
rect -55511 -36198 -55473 -35902
rect -55177 -36198 -55139 -35902
rect -54511 -36198 -54473 -35902
rect -54177 -36198 -54139 -35902
rect -53511 -36198 -53473 -35902
rect -53177 -36198 -53139 -35902
rect -52511 -36198 -52473 -35902
rect -52177 -36198 -52139 -35902
rect -51511 -36198 -51473 -35902
rect -51177 -36198 -51139 -35902
rect -50511 -36198 -50473 -35902
rect -50177 -36198 -50139 -35902
rect -49511 -36198 -49473 -35902
rect -49177 -36198 -49139 -35902
rect -74511 -36204 -74139 -36198
rect -73511 -36204 -73139 -36198
rect -72511 -36204 -72139 -36198
rect -71511 -36204 -71139 -36198
rect -70511 -36204 -70139 -36198
rect -69511 -36204 -69139 -36198
rect -68511 -36204 -68139 -36198
rect -67511 -36204 -67139 -36198
rect -66511 -36204 -66139 -36198
rect -65511 -36204 -65139 -36198
rect -64511 -36204 -64139 -36198
rect -63511 -36204 -63139 -36198
rect -62511 -36204 -62139 -36198
rect -61511 -36204 -61139 -36198
rect -60511 -36204 -60139 -36198
rect -59511 -36204 -59139 -36198
rect -58511 -36204 -58139 -36198
rect -57511 -36204 -57139 -36198
rect -56511 -36204 -56139 -36198
rect -55511 -36204 -55139 -36198
rect -54511 -36204 -54139 -36198
rect -53511 -36204 -53139 -36198
rect -52511 -36204 -52139 -36198
rect -51511 -36204 -51139 -36198
rect -50511 -36204 -50139 -36198
rect -49511 -36204 -49139 -36198
rect -48831 -36204 -48825 -35896
rect -74825 -36210 -48825 -36204
rect -74485 -36236 -74165 -36210
rect -74485 -36864 -74479 -36236
rect -74171 -36864 -74165 -36236
rect -74485 -36890 -74165 -36864
rect -73485 -36236 -73165 -36210
rect -73485 -36864 -73479 -36236
rect -73171 -36864 -73165 -36236
rect -73485 -36890 -73165 -36864
rect -72485 -36236 -72165 -36210
rect -72485 -36864 -72479 -36236
rect -72171 -36864 -72165 -36236
rect -72485 -36890 -72165 -36864
rect -71485 -36236 -71165 -36210
rect -71485 -36864 -71479 -36236
rect -71171 -36864 -71165 -36236
rect -71485 -36890 -71165 -36864
rect -70485 -36236 -70165 -36210
rect -70485 -36864 -70479 -36236
rect -70171 -36864 -70165 -36236
rect -70485 -36890 -70165 -36864
rect -69485 -36236 -69165 -36210
rect -69485 -36864 -69479 -36236
rect -69171 -36864 -69165 -36236
rect -69485 -36890 -69165 -36864
rect -68485 -36236 -68165 -36210
rect -68485 -36864 -68479 -36236
rect -68171 -36864 -68165 -36236
rect -68485 -36890 -68165 -36864
rect -67485 -36236 -67165 -36210
rect -67485 -36864 -67479 -36236
rect -67171 -36864 -67165 -36236
rect -67485 -36890 -67165 -36864
rect -66485 -36236 -66165 -36210
rect -66485 -36864 -66479 -36236
rect -66171 -36864 -66165 -36236
rect -66485 -36890 -66165 -36864
rect -65485 -36236 -65165 -36210
rect -65485 -36864 -65479 -36236
rect -65171 -36864 -65165 -36236
rect -65485 -36890 -65165 -36864
rect -64485 -36236 -64165 -36210
rect -64485 -36864 -64479 -36236
rect -64171 -36864 -64165 -36236
rect -64485 -36890 -64165 -36864
rect -63485 -36236 -63165 -36210
rect -63485 -36864 -63479 -36236
rect -63171 -36864 -63165 -36236
rect -63485 -36890 -63165 -36864
rect -62485 -36236 -62165 -36210
rect -62485 -36864 -62479 -36236
rect -62171 -36864 -62165 -36236
rect -62485 -36890 -62165 -36864
rect -61485 -36236 -61165 -36210
rect -61485 -36864 -61479 -36236
rect -61171 -36864 -61165 -36236
rect -61485 -36890 -61165 -36864
rect -60485 -36236 -60165 -36210
rect -60485 -36864 -60479 -36236
rect -60171 -36864 -60165 -36236
rect -60485 -36890 -60165 -36864
rect -59485 -36236 -59165 -36210
rect -59485 -36864 -59479 -36236
rect -59171 -36864 -59165 -36236
rect -59485 -36890 -59165 -36864
rect -58485 -36236 -58165 -36210
rect -58485 -36864 -58479 -36236
rect -58171 -36864 -58165 -36236
rect -58485 -36890 -58165 -36864
rect -57485 -36236 -57165 -36210
rect -57485 -36864 -57479 -36236
rect -57171 -36864 -57165 -36236
rect -57485 -36890 -57165 -36864
rect -56485 -36236 -56165 -36210
rect -56485 -36864 -56479 -36236
rect -56171 -36864 -56165 -36236
rect -56485 -36890 -56165 -36864
rect -55485 -36236 -55165 -36210
rect -55485 -36864 -55479 -36236
rect -55171 -36864 -55165 -36236
rect -55485 -36890 -55165 -36864
rect -54485 -36236 -54165 -36210
rect -54485 -36864 -54479 -36236
rect -54171 -36864 -54165 -36236
rect -54485 -36890 -54165 -36864
rect -53485 -36236 -53165 -36210
rect -53485 -36864 -53479 -36236
rect -53171 -36864 -53165 -36236
rect -53485 -36890 -53165 -36864
rect -52485 -36236 -52165 -36210
rect -52485 -36864 -52479 -36236
rect -52171 -36864 -52165 -36236
rect -52485 -36890 -52165 -36864
rect -51485 -36236 -51165 -36210
rect -51485 -36864 -51479 -36236
rect -51171 -36864 -51165 -36236
rect -51485 -36890 -51165 -36864
rect -50485 -36236 -50165 -36210
rect -50485 -36864 -50479 -36236
rect -50171 -36864 -50165 -36236
rect -50485 -36890 -50165 -36864
rect -49485 -36236 -49165 -36210
rect -49485 -36864 -49479 -36236
rect -49171 -36864 -49165 -36236
rect -49485 -36890 -49165 -36864
rect -74825 -36896 -48825 -36890
rect -74825 -37204 -74819 -36896
rect -74511 -36902 -74139 -36896
rect -73511 -36902 -73139 -36896
rect -72511 -36902 -72139 -36896
rect -71511 -36902 -71139 -36896
rect -70511 -36902 -70139 -36896
rect -69511 -36902 -69139 -36896
rect -68511 -36902 -68139 -36896
rect -67511 -36902 -67139 -36896
rect -66511 -36902 -66139 -36896
rect -65511 -36902 -65139 -36896
rect -64511 -36902 -64139 -36896
rect -63511 -36902 -63139 -36896
rect -62511 -36902 -62139 -36896
rect -61511 -36902 -61139 -36896
rect -60511 -36902 -60139 -36896
rect -59511 -36902 -59139 -36896
rect -58511 -36902 -58139 -36896
rect -57511 -36902 -57139 -36896
rect -56511 -36902 -56139 -36896
rect -55511 -36902 -55139 -36896
rect -54511 -36902 -54139 -36896
rect -53511 -36902 -53139 -36896
rect -52511 -36902 -52139 -36896
rect -51511 -36902 -51139 -36896
rect -50511 -36902 -50139 -36896
rect -49511 -36902 -49139 -36896
rect -74511 -37198 -74473 -36902
rect -74177 -37198 -74139 -36902
rect -73511 -37198 -73473 -36902
rect -73177 -37198 -73139 -36902
rect -72511 -37198 -72473 -36902
rect -72177 -37198 -72139 -36902
rect -71511 -37198 -71473 -36902
rect -71177 -37198 -71139 -36902
rect -70511 -37198 -70473 -36902
rect -70177 -37198 -70139 -36902
rect -69511 -37198 -69473 -36902
rect -69177 -37198 -69139 -36902
rect -68511 -37198 -68473 -36902
rect -68177 -37198 -68139 -36902
rect -67511 -37198 -67473 -36902
rect -67177 -37198 -67139 -36902
rect -66511 -37198 -66473 -36902
rect -66177 -37198 -66139 -36902
rect -65511 -37198 -65473 -36902
rect -65177 -37198 -65139 -36902
rect -64511 -37198 -64473 -36902
rect -64177 -37198 -64139 -36902
rect -63511 -37198 -63473 -36902
rect -63177 -37198 -63139 -36902
rect -62511 -37198 -62473 -36902
rect -62177 -37198 -62139 -36902
rect -61511 -37198 -61473 -36902
rect -61177 -37198 -61139 -36902
rect -60511 -37198 -60473 -36902
rect -60177 -37198 -60139 -36902
rect -59511 -37198 -59473 -36902
rect -59177 -37198 -59139 -36902
rect -58511 -37198 -58473 -36902
rect -58177 -37198 -58139 -36902
rect -57511 -37198 -57473 -36902
rect -57177 -37198 -57139 -36902
rect -56511 -37198 -56473 -36902
rect -56177 -37198 -56139 -36902
rect -55511 -37198 -55473 -36902
rect -55177 -37198 -55139 -36902
rect -54511 -37198 -54473 -36902
rect -54177 -37198 -54139 -36902
rect -53511 -37198 -53473 -36902
rect -53177 -37198 -53139 -36902
rect -52511 -37198 -52473 -36902
rect -52177 -37198 -52139 -36902
rect -51511 -37198 -51473 -36902
rect -51177 -37198 -51139 -36902
rect -50511 -37198 -50473 -36902
rect -50177 -37198 -50139 -36902
rect -49511 -37198 -49473 -36902
rect -49177 -37198 -49139 -36902
rect -74511 -37204 -74139 -37198
rect -73511 -37204 -73139 -37198
rect -72511 -37204 -72139 -37198
rect -71511 -37204 -71139 -37198
rect -70511 -37204 -70139 -37198
rect -69511 -37204 -69139 -37198
rect -68511 -37204 -68139 -37198
rect -67511 -37204 -67139 -37198
rect -66511 -37204 -66139 -37198
rect -65511 -37204 -65139 -37198
rect -64511 -37204 -64139 -37198
rect -63511 -37204 -63139 -37198
rect -62511 -37204 -62139 -37198
rect -61511 -37204 -61139 -37198
rect -60511 -37204 -60139 -37198
rect -59511 -37204 -59139 -37198
rect -58511 -37204 -58139 -37198
rect -57511 -37204 -57139 -37198
rect -56511 -37204 -56139 -37198
rect -55511 -37204 -55139 -37198
rect -54511 -37204 -54139 -37198
rect -53511 -37204 -53139 -37198
rect -52511 -37204 -52139 -37198
rect -51511 -37204 -51139 -37198
rect -50511 -37204 -50139 -37198
rect -49511 -37204 -49139 -37198
rect -48831 -37204 -48825 -36896
rect -74825 -37210 -48825 -37204
rect -74485 -37236 -74165 -37210
rect -74485 -37864 -74479 -37236
rect -74171 -37864 -74165 -37236
rect -74485 -37890 -74165 -37864
rect -73485 -37236 -73165 -37210
rect -73485 -37864 -73479 -37236
rect -73171 -37864 -73165 -37236
rect -73485 -37890 -73165 -37864
rect -72485 -37236 -72165 -37210
rect -72485 -37864 -72479 -37236
rect -72171 -37864 -72165 -37236
rect -72485 -37890 -72165 -37864
rect -71485 -37236 -71165 -37210
rect -71485 -37864 -71479 -37236
rect -71171 -37864 -71165 -37236
rect -71485 -37890 -71165 -37864
rect -70485 -37236 -70165 -37210
rect -70485 -37864 -70479 -37236
rect -70171 -37864 -70165 -37236
rect -70485 -37890 -70165 -37864
rect -69485 -37236 -69165 -37210
rect -69485 -37864 -69479 -37236
rect -69171 -37864 -69165 -37236
rect -69485 -37890 -69165 -37864
rect -68485 -37236 -68165 -37210
rect -68485 -37864 -68479 -37236
rect -68171 -37864 -68165 -37236
rect -68485 -37890 -68165 -37864
rect -67485 -37236 -67165 -37210
rect -67485 -37864 -67479 -37236
rect -67171 -37864 -67165 -37236
rect -67485 -37890 -67165 -37864
rect -66485 -37236 -66165 -37210
rect -66485 -37864 -66479 -37236
rect -66171 -37864 -66165 -37236
rect -66485 -37890 -66165 -37864
rect -65485 -37236 -65165 -37210
rect -65485 -37864 -65479 -37236
rect -65171 -37864 -65165 -37236
rect -65485 -37890 -65165 -37864
rect -64485 -37236 -64165 -37210
rect -64485 -37864 -64479 -37236
rect -64171 -37864 -64165 -37236
rect -64485 -37890 -64165 -37864
rect -63485 -37236 -63165 -37210
rect -63485 -37864 -63479 -37236
rect -63171 -37864 -63165 -37236
rect -63485 -37890 -63165 -37864
rect -62485 -37236 -62165 -37210
rect -62485 -37864 -62479 -37236
rect -62171 -37864 -62165 -37236
rect -62485 -37890 -62165 -37864
rect -61485 -37236 -61165 -37210
rect -61485 -37864 -61479 -37236
rect -61171 -37864 -61165 -37236
rect -61485 -37890 -61165 -37864
rect -60485 -37236 -60165 -37210
rect -60485 -37864 -60479 -37236
rect -60171 -37864 -60165 -37236
rect -60485 -37890 -60165 -37864
rect -59485 -37236 -59165 -37210
rect -59485 -37864 -59479 -37236
rect -59171 -37864 -59165 -37236
rect -59485 -37890 -59165 -37864
rect -58485 -37236 -58165 -37210
rect -58485 -37864 -58479 -37236
rect -58171 -37864 -58165 -37236
rect -58485 -37890 -58165 -37864
rect -57485 -37236 -57165 -37210
rect -57485 -37864 -57479 -37236
rect -57171 -37864 -57165 -37236
rect -57485 -37890 -57165 -37864
rect -56485 -37236 -56165 -37210
rect -56485 -37864 -56479 -37236
rect -56171 -37864 -56165 -37236
rect -56485 -37890 -56165 -37864
rect -55485 -37236 -55165 -37210
rect -55485 -37864 -55479 -37236
rect -55171 -37864 -55165 -37236
rect -55485 -37890 -55165 -37864
rect -54485 -37236 -54165 -37210
rect -54485 -37864 -54479 -37236
rect -54171 -37864 -54165 -37236
rect -54485 -37890 -54165 -37864
rect -53485 -37236 -53165 -37210
rect -53485 -37864 -53479 -37236
rect -53171 -37864 -53165 -37236
rect -53485 -37890 -53165 -37864
rect -52485 -37236 -52165 -37210
rect -52485 -37864 -52479 -37236
rect -52171 -37864 -52165 -37236
rect -52485 -37890 -52165 -37864
rect -51485 -37236 -51165 -37210
rect -51485 -37864 -51479 -37236
rect -51171 -37864 -51165 -37236
rect -51485 -37890 -51165 -37864
rect -50485 -37236 -50165 -37210
rect -50485 -37864 -50479 -37236
rect -50171 -37864 -50165 -37236
rect -50485 -37890 -50165 -37864
rect -49485 -37236 -49165 -37210
rect -49485 -37864 -49479 -37236
rect -49171 -37864 -49165 -37236
rect -49485 -37890 -49165 -37864
rect -74825 -37896 -48825 -37890
rect -74825 -38204 -74819 -37896
rect -74511 -37902 -74139 -37896
rect -73511 -37902 -73139 -37896
rect -72511 -37902 -72139 -37896
rect -71511 -37902 -71139 -37896
rect -70511 -37902 -70139 -37896
rect -69511 -37902 -69139 -37896
rect -68511 -37902 -68139 -37896
rect -67511 -37902 -67139 -37896
rect -66511 -37902 -66139 -37896
rect -65511 -37902 -65139 -37896
rect -64511 -37902 -64139 -37896
rect -63511 -37902 -63139 -37896
rect -62511 -37902 -62139 -37896
rect -61511 -37902 -61139 -37896
rect -60511 -37902 -60139 -37896
rect -59511 -37902 -59139 -37896
rect -58511 -37902 -58139 -37896
rect -57511 -37902 -57139 -37896
rect -56511 -37902 -56139 -37896
rect -55511 -37902 -55139 -37896
rect -54511 -37902 -54139 -37896
rect -53511 -37902 -53139 -37896
rect -52511 -37902 -52139 -37896
rect -51511 -37902 -51139 -37896
rect -50511 -37902 -50139 -37896
rect -49511 -37902 -49139 -37896
rect -74511 -38198 -74473 -37902
rect -74177 -38198 -74139 -37902
rect -73511 -38198 -73473 -37902
rect -73177 -38198 -73139 -37902
rect -72511 -38198 -72473 -37902
rect -72177 -38198 -72139 -37902
rect -71511 -38198 -71473 -37902
rect -71177 -38198 -71139 -37902
rect -70511 -38198 -70473 -37902
rect -70177 -38198 -70139 -37902
rect -69511 -38198 -69473 -37902
rect -69177 -38198 -69139 -37902
rect -68511 -38198 -68473 -37902
rect -68177 -38198 -68139 -37902
rect -67511 -38198 -67473 -37902
rect -67177 -38198 -67139 -37902
rect -66511 -38198 -66473 -37902
rect -66177 -38198 -66139 -37902
rect -65511 -38198 -65473 -37902
rect -65177 -38198 -65139 -37902
rect -64511 -38198 -64473 -37902
rect -64177 -38198 -64139 -37902
rect -63511 -38198 -63473 -37902
rect -63177 -38198 -63139 -37902
rect -62511 -38198 -62473 -37902
rect -62177 -38198 -62139 -37902
rect -61511 -38198 -61473 -37902
rect -61177 -38198 -61139 -37902
rect -60511 -38198 -60473 -37902
rect -60177 -38198 -60139 -37902
rect -59511 -38198 -59473 -37902
rect -59177 -38198 -59139 -37902
rect -58511 -38198 -58473 -37902
rect -58177 -38198 -58139 -37902
rect -57511 -38198 -57473 -37902
rect -57177 -38198 -57139 -37902
rect -56511 -38198 -56473 -37902
rect -56177 -38198 -56139 -37902
rect -55511 -38198 -55473 -37902
rect -55177 -38198 -55139 -37902
rect -54511 -38198 -54473 -37902
rect -54177 -38198 -54139 -37902
rect -53511 -38198 -53473 -37902
rect -53177 -38198 -53139 -37902
rect -52511 -38198 -52473 -37902
rect -52177 -38198 -52139 -37902
rect -51511 -38198 -51473 -37902
rect -51177 -38198 -51139 -37902
rect -50511 -38198 -50473 -37902
rect -50177 -38198 -50139 -37902
rect -49511 -38198 -49473 -37902
rect -49177 -38198 -49139 -37902
rect -74511 -38204 -74139 -38198
rect -73511 -38204 -73139 -38198
rect -72511 -38204 -72139 -38198
rect -71511 -38204 -71139 -38198
rect -70511 -38204 -70139 -38198
rect -69511 -38204 -69139 -38198
rect -68511 -38204 -68139 -38198
rect -67511 -38204 -67139 -38198
rect -66511 -38204 -66139 -38198
rect -65511 -38204 -65139 -38198
rect -64511 -38204 -64139 -38198
rect -63511 -38204 -63139 -38198
rect -62511 -38204 -62139 -38198
rect -61511 -38204 -61139 -38198
rect -60511 -38204 -60139 -38198
rect -59511 -38204 -59139 -38198
rect -58511 -38204 -58139 -38198
rect -57511 -38204 -57139 -38198
rect -56511 -38204 -56139 -38198
rect -55511 -38204 -55139 -38198
rect -54511 -38204 -54139 -38198
rect -53511 -38204 -53139 -38198
rect -52511 -38204 -52139 -38198
rect -51511 -38204 -51139 -38198
rect -50511 -38204 -50139 -38198
rect -49511 -38204 -49139 -38198
rect -48831 -38204 -48825 -37896
rect -74825 -38210 -48825 -38204
rect -74485 -38236 -74165 -38210
rect -74485 -38864 -74479 -38236
rect -74171 -38864 -74165 -38236
rect -74485 -38890 -74165 -38864
rect -73485 -38236 -73165 -38210
rect -73485 -38864 -73479 -38236
rect -73171 -38864 -73165 -38236
rect -73485 -38890 -73165 -38864
rect -72485 -38236 -72165 -38210
rect -72485 -38864 -72479 -38236
rect -72171 -38864 -72165 -38236
rect -72485 -38890 -72165 -38864
rect -71485 -38236 -71165 -38210
rect -71485 -38864 -71479 -38236
rect -71171 -38864 -71165 -38236
rect -71485 -38890 -71165 -38864
rect -70485 -38236 -70165 -38210
rect -70485 -38864 -70479 -38236
rect -70171 -38864 -70165 -38236
rect -70485 -38890 -70165 -38864
rect -69485 -38236 -69165 -38210
rect -69485 -38864 -69479 -38236
rect -69171 -38864 -69165 -38236
rect -69485 -38890 -69165 -38864
rect -68485 -38236 -68165 -38210
rect -68485 -38864 -68479 -38236
rect -68171 -38864 -68165 -38236
rect -68485 -38890 -68165 -38864
rect -67485 -38236 -67165 -38210
rect -67485 -38864 -67479 -38236
rect -67171 -38864 -67165 -38236
rect -67485 -38890 -67165 -38864
rect -66485 -38236 -66165 -38210
rect -66485 -38864 -66479 -38236
rect -66171 -38864 -66165 -38236
rect -66485 -38890 -66165 -38864
rect -65485 -38236 -65165 -38210
rect -65485 -38864 -65479 -38236
rect -65171 -38864 -65165 -38236
rect -65485 -38890 -65165 -38864
rect -64485 -38236 -64165 -38210
rect -64485 -38864 -64479 -38236
rect -64171 -38864 -64165 -38236
rect -64485 -38890 -64165 -38864
rect -63485 -38236 -63165 -38210
rect -63485 -38864 -63479 -38236
rect -63171 -38864 -63165 -38236
rect -63485 -38890 -63165 -38864
rect -62485 -38236 -62165 -38210
rect -62485 -38864 -62479 -38236
rect -62171 -38864 -62165 -38236
rect -62485 -38890 -62165 -38864
rect -61485 -38236 -61165 -38210
rect -61485 -38864 -61479 -38236
rect -61171 -38864 -61165 -38236
rect -61485 -38890 -61165 -38864
rect -60485 -38236 -60165 -38210
rect -60485 -38864 -60479 -38236
rect -60171 -38864 -60165 -38236
rect -60485 -38890 -60165 -38864
rect -59485 -38236 -59165 -38210
rect -59485 -38864 -59479 -38236
rect -59171 -38864 -59165 -38236
rect -59485 -38890 -59165 -38864
rect -58485 -38236 -58165 -38210
rect -58485 -38864 -58479 -38236
rect -58171 -38864 -58165 -38236
rect -58485 -38890 -58165 -38864
rect -57485 -38236 -57165 -38210
rect -57485 -38864 -57479 -38236
rect -57171 -38864 -57165 -38236
rect -57485 -38890 -57165 -38864
rect -56485 -38236 -56165 -38210
rect -56485 -38864 -56479 -38236
rect -56171 -38864 -56165 -38236
rect -56485 -38890 -56165 -38864
rect -55485 -38236 -55165 -38210
rect -55485 -38864 -55479 -38236
rect -55171 -38864 -55165 -38236
rect -55485 -38890 -55165 -38864
rect -54485 -38236 -54165 -38210
rect -54485 -38864 -54479 -38236
rect -54171 -38864 -54165 -38236
rect -54485 -38890 -54165 -38864
rect -53485 -38236 -53165 -38210
rect -53485 -38864 -53479 -38236
rect -53171 -38864 -53165 -38236
rect -53485 -38890 -53165 -38864
rect -52485 -38236 -52165 -38210
rect -52485 -38864 -52479 -38236
rect -52171 -38864 -52165 -38236
rect -52485 -38890 -52165 -38864
rect -51485 -38236 -51165 -38210
rect -51485 -38864 -51479 -38236
rect -51171 -38864 -51165 -38236
rect -51485 -38890 -51165 -38864
rect -50485 -38236 -50165 -38210
rect -50485 -38864 -50479 -38236
rect -50171 -38864 -50165 -38236
rect -50485 -38890 -50165 -38864
rect -49485 -38236 -49165 -38210
rect -49485 -38864 -49479 -38236
rect -49171 -38864 -49165 -38236
rect -49485 -38890 -49165 -38864
rect -74825 -38896 -48825 -38890
rect -74825 -39204 -74819 -38896
rect -74511 -38902 -74139 -38896
rect -73511 -38902 -73139 -38896
rect -72511 -38902 -72139 -38896
rect -71511 -38902 -71139 -38896
rect -70511 -38902 -70139 -38896
rect -69511 -38902 -69139 -38896
rect -68511 -38902 -68139 -38896
rect -67511 -38902 -67139 -38896
rect -66511 -38902 -66139 -38896
rect -65511 -38902 -65139 -38896
rect -64511 -38902 -64139 -38896
rect -63511 -38902 -63139 -38896
rect -62511 -38902 -62139 -38896
rect -61511 -38902 -61139 -38896
rect -60511 -38902 -60139 -38896
rect -59511 -38902 -59139 -38896
rect -58511 -38902 -58139 -38896
rect -57511 -38902 -57139 -38896
rect -56511 -38902 -56139 -38896
rect -55511 -38902 -55139 -38896
rect -54511 -38902 -54139 -38896
rect -53511 -38902 -53139 -38896
rect -52511 -38902 -52139 -38896
rect -51511 -38902 -51139 -38896
rect -50511 -38902 -50139 -38896
rect -49511 -38902 -49139 -38896
rect -74511 -39198 -74473 -38902
rect -74177 -39198 -74139 -38902
rect -73511 -39198 -73473 -38902
rect -73177 -39198 -73139 -38902
rect -72511 -39198 -72473 -38902
rect -72177 -39198 -72139 -38902
rect -71511 -39198 -71473 -38902
rect -71177 -39198 -71139 -38902
rect -70511 -39198 -70473 -38902
rect -70177 -39198 -70139 -38902
rect -69511 -39198 -69473 -38902
rect -69177 -39198 -69139 -38902
rect -68511 -39198 -68473 -38902
rect -68177 -39198 -68139 -38902
rect -67511 -39198 -67473 -38902
rect -67177 -39198 -67139 -38902
rect -66511 -39198 -66473 -38902
rect -66177 -39198 -66139 -38902
rect -65511 -39198 -65473 -38902
rect -65177 -39198 -65139 -38902
rect -64511 -39198 -64473 -38902
rect -64177 -39198 -64139 -38902
rect -63511 -39198 -63473 -38902
rect -63177 -39198 -63139 -38902
rect -62511 -39198 -62473 -38902
rect -62177 -39198 -62139 -38902
rect -61511 -39198 -61473 -38902
rect -61177 -39198 -61139 -38902
rect -60511 -39198 -60473 -38902
rect -60177 -39198 -60139 -38902
rect -59511 -39198 -59473 -38902
rect -59177 -39198 -59139 -38902
rect -58511 -39198 -58473 -38902
rect -58177 -39198 -58139 -38902
rect -57511 -39198 -57473 -38902
rect -57177 -39198 -57139 -38902
rect -56511 -39198 -56473 -38902
rect -56177 -39198 -56139 -38902
rect -55511 -39198 -55473 -38902
rect -55177 -39198 -55139 -38902
rect -54511 -39198 -54473 -38902
rect -54177 -39198 -54139 -38902
rect -53511 -39198 -53473 -38902
rect -53177 -39198 -53139 -38902
rect -52511 -39198 -52473 -38902
rect -52177 -39198 -52139 -38902
rect -51511 -39198 -51473 -38902
rect -51177 -39198 -51139 -38902
rect -50511 -39198 -50473 -38902
rect -50177 -39198 -50139 -38902
rect -49511 -39198 -49473 -38902
rect -49177 -39198 -49139 -38902
rect -74511 -39204 -74139 -39198
rect -73511 -39204 -73139 -39198
rect -72511 -39204 -72139 -39198
rect -71511 -39204 -71139 -39198
rect -70511 -39204 -70139 -39198
rect -69511 -39204 -69139 -39198
rect -68511 -39204 -68139 -39198
rect -67511 -39204 -67139 -39198
rect -66511 -39204 -66139 -39198
rect -65511 -39204 -65139 -39198
rect -64511 -39204 -64139 -39198
rect -63511 -39204 -63139 -39198
rect -62511 -39204 -62139 -39198
rect -61511 -39204 -61139 -39198
rect -60511 -39204 -60139 -39198
rect -59511 -39204 -59139 -39198
rect -58511 -39204 -58139 -39198
rect -57511 -39204 -57139 -39198
rect -56511 -39204 -56139 -39198
rect -55511 -39204 -55139 -39198
rect -54511 -39204 -54139 -39198
rect -53511 -39204 -53139 -39198
rect -52511 -39204 -52139 -39198
rect -51511 -39204 -51139 -39198
rect -50511 -39204 -50139 -39198
rect -49511 -39204 -49139 -39198
rect -48831 -39204 -48825 -38896
rect -74825 -39210 -48825 -39204
rect -74485 -39236 -74165 -39210
rect -74485 -39864 -74479 -39236
rect -74171 -39864 -74165 -39236
rect -74485 -39890 -74165 -39864
rect -73485 -39236 -73165 -39210
rect -73485 -39864 -73479 -39236
rect -73171 -39864 -73165 -39236
rect -73485 -39890 -73165 -39864
rect -72485 -39236 -72165 -39210
rect -72485 -39864 -72479 -39236
rect -72171 -39864 -72165 -39236
rect -72485 -39890 -72165 -39864
rect -71485 -39236 -71165 -39210
rect -71485 -39864 -71479 -39236
rect -71171 -39864 -71165 -39236
rect -71485 -39890 -71165 -39864
rect -70485 -39236 -70165 -39210
rect -70485 -39864 -70479 -39236
rect -70171 -39864 -70165 -39236
rect -70485 -39890 -70165 -39864
rect -69485 -39236 -69165 -39210
rect -69485 -39864 -69479 -39236
rect -69171 -39864 -69165 -39236
rect -69485 -39890 -69165 -39864
rect -68485 -39236 -68165 -39210
rect -68485 -39864 -68479 -39236
rect -68171 -39864 -68165 -39236
rect -68485 -39890 -68165 -39864
rect -67485 -39236 -67165 -39210
rect -67485 -39864 -67479 -39236
rect -67171 -39864 -67165 -39236
rect -67485 -39890 -67165 -39864
rect -66485 -39236 -66165 -39210
rect -66485 -39864 -66479 -39236
rect -66171 -39864 -66165 -39236
rect -66485 -39890 -66165 -39864
rect -65485 -39236 -65165 -39210
rect -65485 -39864 -65479 -39236
rect -65171 -39864 -65165 -39236
rect -65485 -39890 -65165 -39864
rect -64485 -39236 -64165 -39210
rect -64485 -39864 -64479 -39236
rect -64171 -39864 -64165 -39236
rect -64485 -39890 -64165 -39864
rect -63485 -39236 -63165 -39210
rect -63485 -39864 -63479 -39236
rect -63171 -39864 -63165 -39236
rect -63485 -39890 -63165 -39864
rect -62485 -39236 -62165 -39210
rect -62485 -39864 -62479 -39236
rect -62171 -39864 -62165 -39236
rect -62485 -39890 -62165 -39864
rect -61485 -39236 -61165 -39210
rect -61485 -39864 -61479 -39236
rect -61171 -39864 -61165 -39236
rect -61485 -39890 -61165 -39864
rect -60485 -39236 -60165 -39210
rect -60485 -39864 -60479 -39236
rect -60171 -39864 -60165 -39236
rect -60485 -39890 -60165 -39864
rect -59485 -39236 -59165 -39210
rect -59485 -39864 -59479 -39236
rect -59171 -39864 -59165 -39236
rect -59485 -39890 -59165 -39864
rect -58485 -39236 -58165 -39210
rect -58485 -39864 -58479 -39236
rect -58171 -39864 -58165 -39236
rect -58485 -39890 -58165 -39864
rect -57485 -39236 -57165 -39210
rect -57485 -39864 -57479 -39236
rect -57171 -39864 -57165 -39236
rect -57485 -39890 -57165 -39864
rect -56485 -39236 -56165 -39210
rect -56485 -39864 -56479 -39236
rect -56171 -39864 -56165 -39236
rect -56485 -39890 -56165 -39864
rect -55485 -39236 -55165 -39210
rect -55485 -39864 -55479 -39236
rect -55171 -39864 -55165 -39236
rect -55485 -39890 -55165 -39864
rect -54485 -39236 -54165 -39210
rect -54485 -39864 -54479 -39236
rect -54171 -39864 -54165 -39236
rect -54485 -39890 -54165 -39864
rect -53485 -39236 -53165 -39210
rect -53485 -39864 -53479 -39236
rect -53171 -39864 -53165 -39236
rect -53485 -39890 -53165 -39864
rect -52485 -39236 -52165 -39210
rect -52485 -39864 -52479 -39236
rect -52171 -39864 -52165 -39236
rect -52485 -39890 -52165 -39864
rect -51485 -39236 -51165 -39210
rect -51485 -39864 -51479 -39236
rect -51171 -39864 -51165 -39236
rect -51485 -39890 -51165 -39864
rect -50485 -39236 -50165 -39210
rect -50485 -39864 -50479 -39236
rect -50171 -39864 -50165 -39236
rect -50485 -39890 -50165 -39864
rect -49485 -39236 -49165 -39210
rect -49485 -39864 -49479 -39236
rect -49171 -39864 -49165 -39236
rect -49485 -39890 -49165 -39864
rect -74825 -39896 -48825 -39890
rect -74825 -40204 -74819 -39896
rect -74511 -39902 -74139 -39896
rect -73511 -39902 -73139 -39896
rect -72511 -39902 -72139 -39896
rect -71511 -39902 -71139 -39896
rect -70511 -39902 -70139 -39896
rect -69511 -39902 -69139 -39896
rect -68511 -39902 -68139 -39896
rect -67511 -39902 -67139 -39896
rect -66511 -39902 -66139 -39896
rect -65511 -39902 -65139 -39896
rect -64511 -39902 -64139 -39896
rect -63511 -39902 -63139 -39896
rect -62511 -39902 -62139 -39896
rect -61511 -39902 -61139 -39896
rect -60511 -39902 -60139 -39896
rect -59511 -39902 -59139 -39896
rect -58511 -39902 -58139 -39896
rect -57511 -39902 -57139 -39896
rect -56511 -39902 -56139 -39896
rect -55511 -39902 -55139 -39896
rect -54511 -39902 -54139 -39896
rect -53511 -39902 -53139 -39896
rect -52511 -39902 -52139 -39896
rect -51511 -39902 -51139 -39896
rect -50511 -39902 -50139 -39896
rect -49511 -39902 -49139 -39896
rect -74511 -40198 -74473 -39902
rect -74177 -40198 -74139 -39902
rect -73511 -40198 -73473 -39902
rect -73177 -40198 -73139 -39902
rect -72511 -40198 -72473 -39902
rect -72177 -40198 -72139 -39902
rect -71511 -40198 -71473 -39902
rect -71177 -40198 -71139 -39902
rect -70511 -40198 -70473 -39902
rect -70177 -40198 -70139 -39902
rect -69511 -40198 -69473 -39902
rect -69177 -40198 -69139 -39902
rect -68511 -40198 -68473 -39902
rect -68177 -40198 -68139 -39902
rect -67511 -40198 -67473 -39902
rect -67177 -40198 -67139 -39902
rect -66511 -40198 -66473 -39902
rect -66177 -40198 -66139 -39902
rect -65511 -40198 -65473 -39902
rect -65177 -40198 -65139 -39902
rect -64511 -40198 -64473 -39902
rect -64177 -40198 -64139 -39902
rect -63511 -40198 -63473 -39902
rect -63177 -40198 -63139 -39902
rect -62511 -40198 -62473 -39902
rect -62177 -40198 -62139 -39902
rect -61511 -40198 -61473 -39902
rect -61177 -40198 -61139 -39902
rect -60511 -40198 -60473 -39902
rect -60177 -40198 -60139 -39902
rect -59511 -40198 -59473 -39902
rect -59177 -40198 -59139 -39902
rect -58511 -40198 -58473 -39902
rect -58177 -40198 -58139 -39902
rect -57511 -40198 -57473 -39902
rect -57177 -40198 -57139 -39902
rect -56511 -40198 -56473 -39902
rect -56177 -40198 -56139 -39902
rect -55511 -40198 -55473 -39902
rect -55177 -40198 -55139 -39902
rect -54511 -40198 -54473 -39902
rect -54177 -40198 -54139 -39902
rect -53511 -40198 -53473 -39902
rect -53177 -40198 -53139 -39902
rect -52511 -40198 -52473 -39902
rect -52177 -40198 -52139 -39902
rect -51511 -40198 -51473 -39902
rect -51177 -40198 -51139 -39902
rect -50511 -40198 -50473 -39902
rect -50177 -40198 -50139 -39902
rect -49511 -40198 -49473 -39902
rect -49177 -40198 -49139 -39902
rect -74511 -40204 -74139 -40198
rect -73511 -40204 -73139 -40198
rect -72511 -40204 -72139 -40198
rect -71511 -40204 -71139 -40198
rect -70511 -40204 -70139 -40198
rect -69511 -40204 -69139 -40198
rect -68511 -40204 -68139 -40198
rect -67511 -40204 -67139 -40198
rect -66511 -40204 -66139 -40198
rect -65511 -40204 -65139 -40198
rect -64511 -40204 -64139 -40198
rect -63511 -40204 -63139 -40198
rect -62511 -40204 -62139 -40198
rect -61511 -40204 -61139 -40198
rect -60511 -40204 -60139 -40198
rect -59511 -40204 -59139 -40198
rect -58511 -40204 -58139 -40198
rect -57511 -40204 -57139 -40198
rect -56511 -40204 -56139 -40198
rect -55511 -40204 -55139 -40198
rect -54511 -40204 -54139 -40198
rect -53511 -40204 -53139 -40198
rect -52511 -40204 -52139 -40198
rect -51511 -40204 -51139 -40198
rect -50511 -40204 -50139 -40198
rect -49511 -40204 -49139 -40198
rect -48831 -40204 -48825 -39896
rect -74825 -40210 -48825 -40204
rect -74485 -40236 -74165 -40210
rect -74485 -40864 -74479 -40236
rect -74171 -40864 -74165 -40236
rect -74485 -40890 -74165 -40864
rect -73485 -40236 -73165 -40210
rect -73485 -40864 -73479 -40236
rect -73171 -40864 -73165 -40236
rect -73485 -40890 -73165 -40864
rect -72485 -40236 -72165 -40210
rect -72485 -40864 -72479 -40236
rect -72171 -40864 -72165 -40236
rect -72485 -40890 -72165 -40864
rect -71485 -40236 -71165 -40210
rect -71485 -40864 -71479 -40236
rect -71171 -40864 -71165 -40236
rect -71485 -40890 -71165 -40864
rect -70485 -40236 -70165 -40210
rect -70485 -40864 -70479 -40236
rect -70171 -40864 -70165 -40236
rect -70485 -40890 -70165 -40864
rect -69485 -40236 -69165 -40210
rect -69485 -40864 -69479 -40236
rect -69171 -40864 -69165 -40236
rect -69485 -40890 -69165 -40864
rect -68485 -40236 -68165 -40210
rect -68485 -40864 -68479 -40236
rect -68171 -40864 -68165 -40236
rect -68485 -40890 -68165 -40864
rect -67485 -40236 -67165 -40210
rect -67485 -40864 -67479 -40236
rect -67171 -40864 -67165 -40236
rect -67485 -40890 -67165 -40864
rect -66485 -40236 -66165 -40210
rect -66485 -40864 -66479 -40236
rect -66171 -40864 -66165 -40236
rect -66485 -40890 -66165 -40864
rect -65485 -40236 -65165 -40210
rect -65485 -40864 -65479 -40236
rect -65171 -40864 -65165 -40236
rect -65485 -40890 -65165 -40864
rect -64485 -40236 -64165 -40210
rect -64485 -40864 -64479 -40236
rect -64171 -40864 -64165 -40236
rect -64485 -40890 -64165 -40864
rect -63485 -40236 -63165 -40210
rect -63485 -40864 -63479 -40236
rect -63171 -40864 -63165 -40236
rect -63485 -40890 -63165 -40864
rect -62485 -40236 -62165 -40210
rect -62485 -40864 -62479 -40236
rect -62171 -40864 -62165 -40236
rect -62485 -40890 -62165 -40864
rect -61485 -40236 -61165 -40210
rect -61485 -40864 -61479 -40236
rect -61171 -40864 -61165 -40236
rect -61485 -40890 -61165 -40864
rect -60485 -40236 -60165 -40210
rect -60485 -40864 -60479 -40236
rect -60171 -40864 -60165 -40236
rect -60485 -40890 -60165 -40864
rect -59485 -40236 -59165 -40210
rect -59485 -40864 -59479 -40236
rect -59171 -40864 -59165 -40236
rect -59485 -40890 -59165 -40864
rect -58485 -40236 -58165 -40210
rect -58485 -40864 -58479 -40236
rect -58171 -40864 -58165 -40236
rect -58485 -40890 -58165 -40864
rect -57485 -40236 -57165 -40210
rect -57485 -40864 -57479 -40236
rect -57171 -40864 -57165 -40236
rect -57485 -40890 -57165 -40864
rect -56485 -40236 -56165 -40210
rect -56485 -40864 -56479 -40236
rect -56171 -40864 -56165 -40236
rect -56485 -40890 -56165 -40864
rect -55485 -40236 -55165 -40210
rect -55485 -40864 -55479 -40236
rect -55171 -40864 -55165 -40236
rect -55485 -40890 -55165 -40864
rect -54485 -40236 -54165 -40210
rect -54485 -40864 -54479 -40236
rect -54171 -40864 -54165 -40236
rect -54485 -40890 -54165 -40864
rect -53485 -40236 -53165 -40210
rect -53485 -40864 -53479 -40236
rect -53171 -40864 -53165 -40236
rect -53485 -40890 -53165 -40864
rect -52485 -40236 -52165 -40210
rect -52485 -40864 -52479 -40236
rect -52171 -40864 -52165 -40236
rect -52485 -40890 -52165 -40864
rect -51485 -40236 -51165 -40210
rect -51485 -40864 -51479 -40236
rect -51171 -40864 -51165 -40236
rect -51485 -40890 -51165 -40864
rect -50485 -40236 -50165 -40210
rect -50485 -40864 -50479 -40236
rect -50171 -40864 -50165 -40236
rect -50485 -40890 -50165 -40864
rect -49485 -40236 -49165 -40210
rect -49485 -40864 -49479 -40236
rect -49171 -40864 -49165 -40236
rect -49485 -40890 -49165 -40864
rect -74825 -40896 -48825 -40890
rect -74825 -41204 -74819 -40896
rect -74511 -40902 -74139 -40896
rect -73511 -40902 -73139 -40896
rect -72511 -40902 -72139 -40896
rect -71511 -40902 -71139 -40896
rect -70511 -40902 -70139 -40896
rect -69511 -40902 -69139 -40896
rect -68511 -40902 -68139 -40896
rect -67511 -40902 -67139 -40896
rect -66511 -40902 -66139 -40896
rect -65511 -40902 -65139 -40896
rect -64511 -40902 -64139 -40896
rect -63511 -40902 -63139 -40896
rect -62511 -40902 -62139 -40896
rect -61511 -40902 -61139 -40896
rect -60511 -40902 -60139 -40896
rect -59511 -40902 -59139 -40896
rect -58511 -40902 -58139 -40896
rect -57511 -40902 -57139 -40896
rect -56511 -40902 -56139 -40896
rect -55511 -40902 -55139 -40896
rect -54511 -40902 -54139 -40896
rect -53511 -40902 -53139 -40896
rect -52511 -40902 -52139 -40896
rect -51511 -40902 -51139 -40896
rect -50511 -40902 -50139 -40896
rect -49511 -40902 -49139 -40896
rect -74511 -41198 -74473 -40902
rect -74177 -41198 -74139 -40902
rect -73511 -41198 -73473 -40902
rect -73177 -41198 -73139 -40902
rect -72511 -41198 -72473 -40902
rect -72177 -41198 -72139 -40902
rect -71511 -41198 -71473 -40902
rect -71177 -41198 -71139 -40902
rect -70511 -41198 -70473 -40902
rect -70177 -41198 -70139 -40902
rect -69511 -41198 -69473 -40902
rect -69177 -41198 -69139 -40902
rect -68511 -41198 -68473 -40902
rect -68177 -41198 -68139 -40902
rect -67511 -41198 -67473 -40902
rect -67177 -41198 -67139 -40902
rect -66511 -41198 -66473 -40902
rect -66177 -41198 -66139 -40902
rect -65511 -41198 -65473 -40902
rect -65177 -41198 -65139 -40902
rect -64511 -41198 -64473 -40902
rect -64177 -41198 -64139 -40902
rect -63511 -41198 -63473 -40902
rect -63177 -41198 -63139 -40902
rect -62511 -41198 -62473 -40902
rect -62177 -41198 -62139 -40902
rect -61511 -41198 -61473 -40902
rect -61177 -41198 -61139 -40902
rect -60511 -41198 -60473 -40902
rect -60177 -41198 -60139 -40902
rect -59511 -41198 -59473 -40902
rect -59177 -41198 -59139 -40902
rect -58511 -41198 -58473 -40902
rect -58177 -41198 -58139 -40902
rect -57511 -41198 -57473 -40902
rect -57177 -41198 -57139 -40902
rect -56511 -41198 -56473 -40902
rect -56177 -41198 -56139 -40902
rect -55511 -41198 -55473 -40902
rect -55177 -41198 -55139 -40902
rect -54511 -41198 -54473 -40902
rect -54177 -41198 -54139 -40902
rect -53511 -41198 -53473 -40902
rect -53177 -41198 -53139 -40902
rect -52511 -41198 -52473 -40902
rect -52177 -41198 -52139 -40902
rect -51511 -41198 -51473 -40902
rect -51177 -41198 -51139 -40902
rect -50511 -41198 -50473 -40902
rect -50177 -41198 -50139 -40902
rect -49511 -41198 -49473 -40902
rect -49177 -41198 -49139 -40902
rect -74511 -41204 -74139 -41198
rect -73511 -41204 -73139 -41198
rect -72511 -41204 -72139 -41198
rect -71511 -41204 -71139 -41198
rect -70511 -41204 -70139 -41198
rect -69511 -41204 -69139 -41198
rect -68511 -41204 -68139 -41198
rect -67511 -41204 -67139 -41198
rect -66511 -41204 -66139 -41198
rect -65511 -41204 -65139 -41198
rect -64511 -41204 -64139 -41198
rect -63511 -41204 -63139 -41198
rect -62511 -41204 -62139 -41198
rect -61511 -41204 -61139 -41198
rect -60511 -41204 -60139 -41198
rect -59511 -41204 -59139 -41198
rect -58511 -41204 -58139 -41198
rect -57511 -41204 -57139 -41198
rect -56511 -41204 -56139 -41198
rect -55511 -41204 -55139 -41198
rect -54511 -41204 -54139 -41198
rect -53511 -41204 -53139 -41198
rect -52511 -41204 -52139 -41198
rect -51511 -41204 -51139 -41198
rect -50511 -41204 -50139 -41198
rect -49511 -41204 -49139 -41198
rect -48831 -41204 -48825 -40896
rect -74825 -41210 -48825 -41204
rect -74485 -41236 -74165 -41210
rect -74485 -41864 -74479 -41236
rect -74171 -41864 -74165 -41236
rect -74485 -41890 -74165 -41864
rect -73485 -41236 -73165 -41210
rect -73485 -41864 -73479 -41236
rect -73171 -41864 -73165 -41236
rect -73485 -41890 -73165 -41864
rect -72485 -41236 -72165 -41210
rect -72485 -41864 -72479 -41236
rect -72171 -41864 -72165 -41236
rect -72485 -41890 -72165 -41864
rect -71485 -41236 -71165 -41210
rect -71485 -41864 -71479 -41236
rect -71171 -41864 -71165 -41236
rect -71485 -41890 -71165 -41864
rect -70485 -41236 -70165 -41210
rect -70485 -41864 -70479 -41236
rect -70171 -41864 -70165 -41236
rect -70485 -41890 -70165 -41864
rect -69485 -41236 -69165 -41210
rect -69485 -41864 -69479 -41236
rect -69171 -41864 -69165 -41236
rect -69485 -41890 -69165 -41864
rect -68485 -41236 -68165 -41210
rect -68485 -41864 -68479 -41236
rect -68171 -41864 -68165 -41236
rect -68485 -41890 -68165 -41864
rect -67485 -41236 -67165 -41210
rect -67485 -41864 -67479 -41236
rect -67171 -41864 -67165 -41236
rect -67485 -41890 -67165 -41864
rect -66485 -41236 -66165 -41210
rect -66485 -41864 -66479 -41236
rect -66171 -41864 -66165 -41236
rect -66485 -41890 -66165 -41864
rect -65485 -41236 -65165 -41210
rect -65485 -41864 -65479 -41236
rect -65171 -41864 -65165 -41236
rect -65485 -41890 -65165 -41864
rect -64485 -41236 -64165 -41210
rect -64485 -41864 -64479 -41236
rect -64171 -41864 -64165 -41236
rect -64485 -41890 -64165 -41864
rect -63485 -41236 -63165 -41210
rect -63485 -41864 -63479 -41236
rect -63171 -41864 -63165 -41236
rect -63485 -41890 -63165 -41864
rect -62485 -41236 -62165 -41210
rect -62485 -41864 -62479 -41236
rect -62171 -41864 -62165 -41236
rect -62485 -41890 -62165 -41864
rect -61485 -41236 -61165 -41210
rect -61485 -41864 -61479 -41236
rect -61171 -41864 -61165 -41236
rect -61485 -41890 -61165 -41864
rect -60485 -41236 -60165 -41210
rect -60485 -41864 -60479 -41236
rect -60171 -41864 -60165 -41236
rect -60485 -41890 -60165 -41864
rect -59485 -41236 -59165 -41210
rect -59485 -41864 -59479 -41236
rect -59171 -41864 -59165 -41236
rect -59485 -41890 -59165 -41864
rect -58485 -41236 -58165 -41210
rect -58485 -41864 -58479 -41236
rect -58171 -41864 -58165 -41236
rect -58485 -41890 -58165 -41864
rect -57485 -41236 -57165 -41210
rect -57485 -41864 -57479 -41236
rect -57171 -41864 -57165 -41236
rect -57485 -41890 -57165 -41864
rect -56485 -41236 -56165 -41210
rect -56485 -41864 -56479 -41236
rect -56171 -41864 -56165 -41236
rect -56485 -41890 -56165 -41864
rect -55485 -41236 -55165 -41210
rect -55485 -41864 -55479 -41236
rect -55171 -41864 -55165 -41236
rect -55485 -41890 -55165 -41864
rect -54485 -41236 -54165 -41210
rect -54485 -41864 -54479 -41236
rect -54171 -41864 -54165 -41236
rect -54485 -41890 -54165 -41864
rect -53485 -41236 -53165 -41210
rect -53485 -41864 -53479 -41236
rect -53171 -41864 -53165 -41236
rect -53485 -41890 -53165 -41864
rect -52485 -41236 -52165 -41210
rect -52485 -41864 -52479 -41236
rect -52171 -41864 -52165 -41236
rect -52485 -41890 -52165 -41864
rect -51485 -41236 -51165 -41210
rect -51485 -41864 -51479 -41236
rect -51171 -41864 -51165 -41236
rect -51485 -41890 -51165 -41864
rect -50485 -41236 -50165 -41210
rect -50485 -41864 -50479 -41236
rect -50171 -41864 -50165 -41236
rect -50485 -41890 -50165 -41864
rect -49485 -41236 -49165 -41210
rect -49485 -41864 -49479 -41236
rect -49171 -41864 -49165 -41236
rect -49485 -41890 -49165 -41864
rect -74825 -41896 -48825 -41890
rect -74825 -42204 -74819 -41896
rect -74511 -41902 -74139 -41896
rect -73511 -41902 -73139 -41896
rect -72511 -41902 -72139 -41896
rect -71511 -41902 -71139 -41896
rect -70511 -41902 -70139 -41896
rect -69511 -41902 -69139 -41896
rect -68511 -41902 -68139 -41896
rect -67511 -41902 -67139 -41896
rect -66511 -41902 -66139 -41896
rect -65511 -41902 -65139 -41896
rect -64511 -41902 -64139 -41896
rect -63511 -41902 -63139 -41896
rect -62511 -41902 -62139 -41896
rect -61511 -41902 -61139 -41896
rect -60511 -41902 -60139 -41896
rect -59511 -41902 -59139 -41896
rect -58511 -41902 -58139 -41896
rect -57511 -41902 -57139 -41896
rect -56511 -41902 -56139 -41896
rect -55511 -41902 -55139 -41896
rect -54511 -41902 -54139 -41896
rect -53511 -41902 -53139 -41896
rect -52511 -41902 -52139 -41896
rect -51511 -41902 -51139 -41896
rect -50511 -41902 -50139 -41896
rect -49511 -41902 -49139 -41896
rect -74511 -42198 -74473 -41902
rect -74177 -42198 -74139 -41902
rect -73511 -42198 -73473 -41902
rect -73177 -42198 -73139 -41902
rect -72511 -42198 -72473 -41902
rect -72177 -42198 -72139 -41902
rect -71511 -42198 -71473 -41902
rect -71177 -42198 -71139 -41902
rect -70511 -42198 -70473 -41902
rect -70177 -42198 -70139 -41902
rect -69511 -42198 -69473 -41902
rect -69177 -42198 -69139 -41902
rect -68511 -42198 -68473 -41902
rect -68177 -42198 -68139 -41902
rect -67511 -42198 -67473 -41902
rect -67177 -42198 -67139 -41902
rect -66511 -42198 -66473 -41902
rect -66177 -42198 -66139 -41902
rect -65511 -42198 -65473 -41902
rect -65177 -42198 -65139 -41902
rect -64511 -42198 -64473 -41902
rect -64177 -42198 -64139 -41902
rect -63511 -42198 -63473 -41902
rect -63177 -42198 -63139 -41902
rect -62511 -42198 -62473 -41902
rect -62177 -42198 -62139 -41902
rect -61511 -42198 -61473 -41902
rect -61177 -42198 -61139 -41902
rect -60511 -42198 -60473 -41902
rect -60177 -42198 -60139 -41902
rect -59511 -42198 -59473 -41902
rect -59177 -42198 -59139 -41902
rect -58511 -42198 -58473 -41902
rect -58177 -42198 -58139 -41902
rect -57511 -42198 -57473 -41902
rect -57177 -42198 -57139 -41902
rect -56511 -42198 -56473 -41902
rect -56177 -42198 -56139 -41902
rect -55511 -42198 -55473 -41902
rect -55177 -42198 -55139 -41902
rect -54511 -42198 -54473 -41902
rect -54177 -42198 -54139 -41902
rect -53511 -42198 -53473 -41902
rect -53177 -42198 -53139 -41902
rect -52511 -42198 -52473 -41902
rect -52177 -42198 -52139 -41902
rect -51511 -42198 -51473 -41902
rect -51177 -42198 -51139 -41902
rect -50511 -42198 -50473 -41902
rect -50177 -42198 -50139 -41902
rect -49511 -42198 -49473 -41902
rect -49177 -42198 -49139 -41902
rect -74511 -42204 -74139 -42198
rect -73511 -42204 -73139 -42198
rect -72511 -42204 -72139 -42198
rect -71511 -42204 -71139 -42198
rect -70511 -42204 -70139 -42198
rect -69511 -42204 -69139 -42198
rect -68511 -42204 -68139 -42198
rect -67511 -42204 -67139 -42198
rect -66511 -42204 -66139 -42198
rect -65511 -42204 -65139 -42198
rect -64511 -42204 -64139 -42198
rect -63511 -42204 -63139 -42198
rect -62511 -42204 -62139 -42198
rect -61511 -42204 -61139 -42198
rect -60511 -42204 -60139 -42198
rect -59511 -42204 -59139 -42198
rect -58511 -42204 -58139 -42198
rect -57511 -42204 -57139 -42198
rect -56511 -42204 -56139 -42198
rect -55511 -42204 -55139 -42198
rect -54511 -42204 -54139 -42198
rect -53511 -42204 -53139 -42198
rect -52511 -42204 -52139 -42198
rect -51511 -42204 -51139 -42198
rect -50511 -42204 -50139 -42198
rect -49511 -42204 -49139 -42198
rect -48831 -42204 -48825 -41896
rect -74825 -42210 -48825 -42204
rect -74485 -42236 -74165 -42210
rect -74485 -42864 -74479 -42236
rect -74171 -42864 -74165 -42236
rect -74485 -42890 -74165 -42864
rect -73485 -42236 -73165 -42210
rect -73485 -42864 -73479 -42236
rect -73171 -42864 -73165 -42236
rect -73485 -42890 -73165 -42864
rect -72485 -42236 -72165 -42210
rect -72485 -42864 -72479 -42236
rect -72171 -42864 -72165 -42236
rect -72485 -42890 -72165 -42864
rect -71485 -42236 -71165 -42210
rect -71485 -42864 -71479 -42236
rect -71171 -42864 -71165 -42236
rect -71485 -42890 -71165 -42864
rect -70485 -42236 -70165 -42210
rect -70485 -42864 -70479 -42236
rect -70171 -42864 -70165 -42236
rect -70485 -42890 -70165 -42864
rect -69485 -42236 -69165 -42210
rect -69485 -42864 -69479 -42236
rect -69171 -42864 -69165 -42236
rect -69485 -42890 -69165 -42864
rect -68485 -42236 -68165 -42210
rect -68485 -42864 -68479 -42236
rect -68171 -42864 -68165 -42236
rect -68485 -42890 -68165 -42864
rect -67485 -42236 -67165 -42210
rect -67485 -42864 -67479 -42236
rect -67171 -42864 -67165 -42236
rect -67485 -42890 -67165 -42864
rect -66485 -42236 -66165 -42210
rect -66485 -42864 -66479 -42236
rect -66171 -42864 -66165 -42236
rect -66485 -42890 -66165 -42864
rect -65485 -42236 -65165 -42210
rect -65485 -42864 -65479 -42236
rect -65171 -42864 -65165 -42236
rect -65485 -42890 -65165 -42864
rect -64485 -42236 -64165 -42210
rect -64485 -42864 -64479 -42236
rect -64171 -42864 -64165 -42236
rect -64485 -42890 -64165 -42864
rect -63485 -42236 -63165 -42210
rect -63485 -42864 -63479 -42236
rect -63171 -42864 -63165 -42236
rect -63485 -42890 -63165 -42864
rect -62485 -42236 -62165 -42210
rect -62485 -42864 -62479 -42236
rect -62171 -42864 -62165 -42236
rect -62485 -42890 -62165 -42864
rect -61485 -42236 -61165 -42210
rect -61485 -42864 -61479 -42236
rect -61171 -42864 -61165 -42236
rect -61485 -42890 -61165 -42864
rect -60485 -42236 -60165 -42210
rect -60485 -42864 -60479 -42236
rect -60171 -42864 -60165 -42236
rect -60485 -42890 -60165 -42864
rect -59485 -42236 -59165 -42210
rect -59485 -42864 -59479 -42236
rect -59171 -42864 -59165 -42236
rect -59485 -42890 -59165 -42864
rect -58485 -42236 -58165 -42210
rect -58485 -42864 -58479 -42236
rect -58171 -42864 -58165 -42236
rect -58485 -42890 -58165 -42864
rect -57485 -42236 -57165 -42210
rect -57485 -42864 -57479 -42236
rect -57171 -42864 -57165 -42236
rect -57485 -42890 -57165 -42864
rect -56485 -42236 -56165 -42210
rect -56485 -42864 -56479 -42236
rect -56171 -42864 -56165 -42236
rect -56485 -42890 -56165 -42864
rect -55485 -42236 -55165 -42210
rect -55485 -42864 -55479 -42236
rect -55171 -42864 -55165 -42236
rect -55485 -42890 -55165 -42864
rect -54485 -42236 -54165 -42210
rect -54485 -42864 -54479 -42236
rect -54171 -42864 -54165 -42236
rect -54485 -42890 -54165 -42864
rect -53485 -42236 -53165 -42210
rect -53485 -42864 -53479 -42236
rect -53171 -42864 -53165 -42236
rect -53485 -42890 -53165 -42864
rect -52485 -42236 -52165 -42210
rect -52485 -42864 -52479 -42236
rect -52171 -42864 -52165 -42236
rect -52485 -42890 -52165 -42864
rect -51485 -42236 -51165 -42210
rect -51485 -42864 -51479 -42236
rect -51171 -42864 -51165 -42236
rect -51485 -42890 -51165 -42864
rect -50485 -42236 -50165 -42210
rect -50485 -42864 -50479 -42236
rect -50171 -42864 -50165 -42236
rect -50485 -42890 -50165 -42864
rect -49485 -42236 -49165 -42210
rect -49485 -42864 -49479 -42236
rect -49171 -42864 -49165 -42236
rect -49485 -42890 -49165 -42864
rect -74825 -42896 -48825 -42890
rect -74825 -43204 -74819 -42896
rect -74511 -42902 -74139 -42896
rect -73511 -42902 -73139 -42896
rect -72511 -42902 -72139 -42896
rect -71511 -42902 -71139 -42896
rect -70511 -42902 -70139 -42896
rect -69511 -42902 -69139 -42896
rect -68511 -42902 -68139 -42896
rect -67511 -42902 -67139 -42896
rect -66511 -42902 -66139 -42896
rect -65511 -42902 -65139 -42896
rect -64511 -42902 -64139 -42896
rect -63511 -42902 -63139 -42896
rect -62511 -42902 -62139 -42896
rect -61511 -42902 -61139 -42896
rect -60511 -42902 -60139 -42896
rect -59511 -42902 -59139 -42896
rect -58511 -42902 -58139 -42896
rect -57511 -42902 -57139 -42896
rect -56511 -42902 -56139 -42896
rect -55511 -42902 -55139 -42896
rect -54511 -42902 -54139 -42896
rect -53511 -42902 -53139 -42896
rect -52511 -42902 -52139 -42896
rect -51511 -42902 -51139 -42896
rect -50511 -42902 -50139 -42896
rect -49511 -42902 -49139 -42896
rect -74511 -43198 -74473 -42902
rect -74177 -43198 -74139 -42902
rect -73511 -43198 -73473 -42902
rect -73177 -43198 -73139 -42902
rect -72511 -43198 -72473 -42902
rect -72177 -43198 -72139 -42902
rect -71511 -43198 -71473 -42902
rect -71177 -43198 -71139 -42902
rect -70511 -43198 -70473 -42902
rect -70177 -43198 -70139 -42902
rect -69511 -43198 -69473 -42902
rect -69177 -43198 -69139 -42902
rect -68511 -43198 -68473 -42902
rect -68177 -43198 -68139 -42902
rect -67511 -43198 -67473 -42902
rect -67177 -43198 -67139 -42902
rect -66511 -43198 -66473 -42902
rect -66177 -43198 -66139 -42902
rect -65511 -43198 -65473 -42902
rect -65177 -43198 -65139 -42902
rect -64511 -43198 -64473 -42902
rect -64177 -43198 -64139 -42902
rect -63511 -43198 -63473 -42902
rect -63177 -43198 -63139 -42902
rect -62511 -43198 -62473 -42902
rect -62177 -43198 -62139 -42902
rect -61511 -43198 -61473 -42902
rect -61177 -43198 -61139 -42902
rect -60511 -43198 -60473 -42902
rect -60177 -43198 -60139 -42902
rect -59511 -43198 -59473 -42902
rect -59177 -43198 -59139 -42902
rect -58511 -43198 -58473 -42902
rect -58177 -43198 -58139 -42902
rect -57511 -43198 -57473 -42902
rect -57177 -43198 -57139 -42902
rect -56511 -43198 -56473 -42902
rect -56177 -43198 -56139 -42902
rect -55511 -43198 -55473 -42902
rect -55177 -43198 -55139 -42902
rect -54511 -43198 -54473 -42902
rect -54177 -43198 -54139 -42902
rect -53511 -43198 -53473 -42902
rect -53177 -43198 -53139 -42902
rect -52511 -43198 -52473 -42902
rect -52177 -43198 -52139 -42902
rect -51511 -43198 -51473 -42902
rect -51177 -43198 -51139 -42902
rect -50511 -43198 -50473 -42902
rect -50177 -43198 -50139 -42902
rect -49511 -43198 -49473 -42902
rect -49177 -43198 -49139 -42902
rect -74511 -43204 -74139 -43198
rect -73511 -43204 -73139 -43198
rect -72511 -43204 -72139 -43198
rect -71511 -43204 -71139 -43198
rect -70511 -43204 -70139 -43198
rect -69511 -43204 -69139 -43198
rect -68511 -43204 -68139 -43198
rect -67511 -43204 -67139 -43198
rect -66511 -43204 -66139 -43198
rect -65511 -43204 -65139 -43198
rect -64511 -43204 -64139 -43198
rect -63511 -43204 -63139 -43198
rect -62511 -43204 -62139 -43198
rect -61511 -43204 -61139 -43198
rect -60511 -43204 -60139 -43198
rect -59511 -43204 -59139 -43198
rect -58511 -43204 -58139 -43198
rect -57511 -43204 -57139 -43198
rect -56511 -43204 -56139 -43198
rect -55511 -43204 -55139 -43198
rect -54511 -43204 -54139 -43198
rect -53511 -43204 -53139 -43198
rect -52511 -43204 -52139 -43198
rect -51511 -43204 -51139 -43198
rect -50511 -43204 -50139 -43198
rect -49511 -43204 -49139 -43198
rect -48831 -43204 -48825 -42896
rect -74825 -43210 -48825 -43204
rect -74485 -43236 -74165 -43210
rect -74485 -43864 -74479 -43236
rect -74171 -43864 -74165 -43236
rect -74485 -43890 -74165 -43864
rect -73485 -43236 -73165 -43210
rect -73485 -43864 -73479 -43236
rect -73171 -43864 -73165 -43236
rect -73485 -43890 -73165 -43864
rect -72485 -43236 -72165 -43210
rect -72485 -43864 -72479 -43236
rect -72171 -43864 -72165 -43236
rect -72485 -43890 -72165 -43864
rect -71485 -43236 -71165 -43210
rect -71485 -43864 -71479 -43236
rect -71171 -43864 -71165 -43236
rect -71485 -43890 -71165 -43864
rect -70485 -43236 -70165 -43210
rect -70485 -43864 -70479 -43236
rect -70171 -43864 -70165 -43236
rect -70485 -43890 -70165 -43864
rect -69485 -43236 -69165 -43210
rect -69485 -43864 -69479 -43236
rect -69171 -43864 -69165 -43236
rect -69485 -43890 -69165 -43864
rect -68485 -43236 -68165 -43210
rect -68485 -43864 -68479 -43236
rect -68171 -43864 -68165 -43236
rect -68485 -43890 -68165 -43864
rect -67485 -43236 -67165 -43210
rect -67485 -43864 -67479 -43236
rect -67171 -43864 -67165 -43236
rect -67485 -43890 -67165 -43864
rect -66485 -43236 -66165 -43210
rect -66485 -43864 -66479 -43236
rect -66171 -43864 -66165 -43236
rect -66485 -43890 -66165 -43864
rect -65485 -43236 -65165 -43210
rect -65485 -43864 -65479 -43236
rect -65171 -43864 -65165 -43236
rect -65485 -43890 -65165 -43864
rect -64485 -43236 -64165 -43210
rect -64485 -43864 -64479 -43236
rect -64171 -43864 -64165 -43236
rect -64485 -43890 -64165 -43864
rect -63485 -43236 -63165 -43210
rect -63485 -43864 -63479 -43236
rect -63171 -43864 -63165 -43236
rect -63485 -43890 -63165 -43864
rect -62485 -43236 -62165 -43210
rect -62485 -43864 -62479 -43236
rect -62171 -43864 -62165 -43236
rect -62485 -43890 -62165 -43864
rect -61485 -43236 -61165 -43210
rect -61485 -43864 -61479 -43236
rect -61171 -43864 -61165 -43236
rect -61485 -43890 -61165 -43864
rect -60485 -43236 -60165 -43210
rect -60485 -43864 -60479 -43236
rect -60171 -43864 -60165 -43236
rect -60485 -43890 -60165 -43864
rect -59485 -43236 -59165 -43210
rect -59485 -43864 -59479 -43236
rect -59171 -43864 -59165 -43236
rect -59485 -43890 -59165 -43864
rect -58485 -43236 -58165 -43210
rect -58485 -43864 -58479 -43236
rect -58171 -43864 -58165 -43236
rect -58485 -43890 -58165 -43864
rect -57485 -43236 -57165 -43210
rect -57485 -43864 -57479 -43236
rect -57171 -43864 -57165 -43236
rect -57485 -43890 -57165 -43864
rect -56485 -43236 -56165 -43210
rect -56485 -43864 -56479 -43236
rect -56171 -43864 -56165 -43236
rect -56485 -43890 -56165 -43864
rect -55485 -43236 -55165 -43210
rect -55485 -43864 -55479 -43236
rect -55171 -43864 -55165 -43236
rect -55485 -43890 -55165 -43864
rect -54485 -43236 -54165 -43210
rect -54485 -43864 -54479 -43236
rect -54171 -43864 -54165 -43236
rect -54485 -43890 -54165 -43864
rect -53485 -43236 -53165 -43210
rect -53485 -43864 -53479 -43236
rect -53171 -43864 -53165 -43236
rect -53485 -43890 -53165 -43864
rect -52485 -43236 -52165 -43210
rect -52485 -43864 -52479 -43236
rect -52171 -43864 -52165 -43236
rect -52485 -43890 -52165 -43864
rect -51485 -43236 -51165 -43210
rect -51485 -43864 -51479 -43236
rect -51171 -43864 -51165 -43236
rect -51485 -43890 -51165 -43864
rect -50485 -43236 -50165 -43210
rect -50485 -43864 -50479 -43236
rect -50171 -43864 -50165 -43236
rect -50485 -43890 -50165 -43864
rect -49485 -43236 -49165 -43210
rect -49485 -43864 -49479 -43236
rect -49171 -43864 -49165 -43236
rect -49485 -43890 -49165 -43864
rect -74825 -43896 -48825 -43890
rect -74825 -44204 -74819 -43896
rect -74511 -43902 -74139 -43896
rect -73511 -43902 -73139 -43896
rect -72511 -43902 -72139 -43896
rect -71511 -43902 -71139 -43896
rect -70511 -43902 -70139 -43896
rect -69511 -43902 -69139 -43896
rect -68511 -43902 -68139 -43896
rect -67511 -43902 -67139 -43896
rect -66511 -43902 -66139 -43896
rect -65511 -43902 -65139 -43896
rect -64511 -43902 -64139 -43896
rect -63511 -43902 -63139 -43896
rect -62511 -43902 -62139 -43896
rect -61511 -43902 -61139 -43896
rect -60511 -43902 -60139 -43896
rect -59511 -43902 -59139 -43896
rect -58511 -43902 -58139 -43896
rect -57511 -43902 -57139 -43896
rect -56511 -43902 -56139 -43896
rect -55511 -43902 -55139 -43896
rect -54511 -43902 -54139 -43896
rect -53511 -43902 -53139 -43896
rect -52511 -43902 -52139 -43896
rect -51511 -43902 -51139 -43896
rect -50511 -43902 -50139 -43896
rect -49511 -43902 -49139 -43896
rect -74511 -44198 -74473 -43902
rect -74177 -44198 -74139 -43902
rect -73511 -44198 -73473 -43902
rect -73177 -44198 -73139 -43902
rect -72511 -44198 -72473 -43902
rect -72177 -44198 -72139 -43902
rect -71511 -44198 -71473 -43902
rect -71177 -44198 -71139 -43902
rect -70511 -44198 -70473 -43902
rect -70177 -44198 -70139 -43902
rect -69511 -44198 -69473 -43902
rect -69177 -44198 -69139 -43902
rect -68511 -44198 -68473 -43902
rect -68177 -44198 -68139 -43902
rect -67511 -44198 -67473 -43902
rect -67177 -44198 -67139 -43902
rect -66511 -44198 -66473 -43902
rect -66177 -44198 -66139 -43902
rect -65511 -44198 -65473 -43902
rect -65177 -44198 -65139 -43902
rect -64511 -44198 -64473 -43902
rect -64177 -44198 -64139 -43902
rect -63511 -44198 -63473 -43902
rect -63177 -44198 -63139 -43902
rect -62511 -44198 -62473 -43902
rect -62177 -44198 -62139 -43902
rect -61511 -44198 -61473 -43902
rect -61177 -44198 -61139 -43902
rect -60511 -44198 -60473 -43902
rect -60177 -44198 -60139 -43902
rect -59511 -44198 -59473 -43902
rect -59177 -44198 -59139 -43902
rect -58511 -44198 -58473 -43902
rect -58177 -44198 -58139 -43902
rect -57511 -44198 -57473 -43902
rect -57177 -44198 -57139 -43902
rect -56511 -44198 -56473 -43902
rect -56177 -44198 -56139 -43902
rect -55511 -44198 -55473 -43902
rect -55177 -44198 -55139 -43902
rect -54511 -44198 -54473 -43902
rect -54177 -44198 -54139 -43902
rect -53511 -44198 -53473 -43902
rect -53177 -44198 -53139 -43902
rect -52511 -44198 -52473 -43902
rect -52177 -44198 -52139 -43902
rect -51511 -44198 -51473 -43902
rect -51177 -44198 -51139 -43902
rect -50511 -44198 -50473 -43902
rect -50177 -44198 -50139 -43902
rect -49511 -44198 -49473 -43902
rect -49177 -44198 -49139 -43902
rect -74511 -44204 -74139 -44198
rect -73511 -44204 -73139 -44198
rect -72511 -44204 -72139 -44198
rect -71511 -44204 -71139 -44198
rect -70511 -44204 -70139 -44198
rect -69511 -44204 -69139 -44198
rect -68511 -44204 -68139 -44198
rect -67511 -44204 -67139 -44198
rect -66511 -44204 -66139 -44198
rect -65511 -44204 -65139 -44198
rect -64511 -44204 -64139 -44198
rect -63511 -44204 -63139 -44198
rect -62511 -44204 -62139 -44198
rect -61511 -44204 -61139 -44198
rect -60511 -44204 -60139 -44198
rect -59511 -44204 -59139 -44198
rect -58511 -44204 -58139 -44198
rect -57511 -44204 -57139 -44198
rect -56511 -44204 -56139 -44198
rect -55511 -44204 -55139 -44198
rect -54511 -44204 -54139 -44198
rect -53511 -44204 -53139 -44198
rect -52511 -44204 -52139 -44198
rect -51511 -44204 -51139 -44198
rect -50511 -44204 -50139 -44198
rect -49511 -44204 -49139 -44198
rect -48831 -44204 -48825 -43896
rect -74825 -44210 -48825 -44204
rect -74485 -44236 -74165 -44210
rect -74485 -44864 -74479 -44236
rect -74171 -44864 -74165 -44236
rect -74485 -44890 -74165 -44864
rect -73485 -44236 -73165 -44210
rect -73485 -44864 -73479 -44236
rect -73171 -44864 -73165 -44236
rect -73485 -44890 -73165 -44864
rect -72485 -44236 -72165 -44210
rect -72485 -44864 -72479 -44236
rect -72171 -44864 -72165 -44236
rect -72485 -44890 -72165 -44864
rect -71485 -44236 -71165 -44210
rect -71485 -44864 -71479 -44236
rect -71171 -44864 -71165 -44236
rect -71485 -44890 -71165 -44864
rect -70485 -44236 -70165 -44210
rect -70485 -44864 -70479 -44236
rect -70171 -44864 -70165 -44236
rect -70485 -44890 -70165 -44864
rect -69485 -44236 -69165 -44210
rect -69485 -44864 -69479 -44236
rect -69171 -44864 -69165 -44236
rect -69485 -44890 -69165 -44864
rect -68485 -44236 -68165 -44210
rect -68485 -44864 -68479 -44236
rect -68171 -44864 -68165 -44236
rect -68485 -44890 -68165 -44864
rect -67485 -44236 -67165 -44210
rect -67485 -44864 -67479 -44236
rect -67171 -44864 -67165 -44236
rect -67485 -44890 -67165 -44864
rect -66485 -44236 -66165 -44210
rect -66485 -44864 -66479 -44236
rect -66171 -44864 -66165 -44236
rect -66485 -44890 -66165 -44864
rect -65485 -44236 -65165 -44210
rect -65485 -44864 -65479 -44236
rect -65171 -44864 -65165 -44236
rect -65485 -44890 -65165 -44864
rect -64485 -44236 -64165 -44210
rect -64485 -44864 -64479 -44236
rect -64171 -44864 -64165 -44236
rect -64485 -44890 -64165 -44864
rect -63485 -44236 -63165 -44210
rect -63485 -44864 -63479 -44236
rect -63171 -44864 -63165 -44236
rect -63485 -44890 -63165 -44864
rect -62485 -44236 -62165 -44210
rect -62485 -44864 -62479 -44236
rect -62171 -44864 -62165 -44236
rect -62485 -44890 -62165 -44864
rect -61485 -44236 -61165 -44210
rect -61485 -44864 -61479 -44236
rect -61171 -44864 -61165 -44236
rect -61485 -44890 -61165 -44864
rect -60485 -44236 -60165 -44210
rect -60485 -44864 -60479 -44236
rect -60171 -44864 -60165 -44236
rect -60485 -44890 -60165 -44864
rect -59485 -44236 -59165 -44210
rect -59485 -44864 -59479 -44236
rect -59171 -44864 -59165 -44236
rect -59485 -44890 -59165 -44864
rect -58485 -44236 -58165 -44210
rect -58485 -44864 -58479 -44236
rect -58171 -44864 -58165 -44236
rect -58485 -44890 -58165 -44864
rect -57485 -44236 -57165 -44210
rect -57485 -44864 -57479 -44236
rect -57171 -44864 -57165 -44236
rect -57485 -44890 -57165 -44864
rect -56485 -44236 -56165 -44210
rect -56485 -44864 -56479 -44236
rect -56171 -44864 -56165 -44236
rect -56485 -44890 -56165 -44864
rect -55485 -44236 -55165 -44210
rect -55485 -44864 -55479 -44236
rect -55171 -44864 -55165 -44236
rect -55485 -44890 -55165 -44864
rect -54485 -44236 -54165 -44210
rect -54485 -44864 -54479 -44236
rect -54171 -44864 -54165 -44236
rect -54485 -44890 -54165 -44864
rect -53485 -44236 -53165 -44210
rect -53485 -44864 -53479 -44236
rect -53171 -44864 -53165 -44236
rect -53485 -44890 -53165 -44864
rect -52485 -44236 -52165 -44210
rect -52485 -44864 -52479 -44236
rect -52171 -44864 -52165 -44236
rect -52485 -44890 -52165 -44864
rect -51485 -44236 -51165 -44210
rect -51485 -44864 -51479 -44236
rect -51171 -44864 -51165 -44236
rect -51485 -44890 -51165 -44864
rect -50485 -44236 -50165 -44210
rect -50485 -44864 -50479 -44236
rect -50171 -44864 -50165 -44236
rect -50485 -44890 -50165 -44864
rect -49485 -44236 -49165 -44210
rect -49485 -44864 -49479 -44236
rect -49171 -44864 -49165 -44236
rect -46275 -44496 -46234 -32604
rect -36326 -44496 -36275 -32604
rect -46275 -44498 -46228 -44496
rect -36332 -44498 -36275 -44496
rect -46275 -44550 -36275 -44498
rect -4275 -32602 5725 -32550
rect -4275 -32604 -4228 -32602
rect 5668 -32604 5725 -32602
rect -4275 -44496 -4234 -32604
rect 5674 -44496 5725 -32604
rect 8615 -32864 8621 -32236
rect 8929 -32864 8935 -32236
rect 8615 -32890 8935 -32864
rect 9615 -32236 9935 -32210
rect 9615 -32864 9621 -32236
rect 9929 -32864 9935 -32236
rect 9615 -32890 9935 -32864
rect 10615 -32236 10935 -32210
rect 10615 -32864 10621 -32236
rect 10929 -32864 10935 -32236
rect 10615 -32890 10935 -32864
rect 11615 -32236 11935 -32210
rect 11615 -32864 11621 -32236
rect 11929 -32864 11935 -32236
rect 11615 -32890 11935 -32864
rect 12615 -32236 12935 -32210
rect 12615 -32864 12621 -32236
rect 12929 -32864 12935 -32236
rect 12615 -32890 12935 -32864
rect 13615 -32236 13935 -32210
rect 13615 -32864 13621 -32236
rect 13929 -32864 13935 -32236
rect 13615 -32890 13935 -32864
rect 14615 -32236 14935 -32210
rect 14615 -32864 14621 -32236
rect 14929 -32864 14935 -32236
rect 14615 -32890 14935 -32864
rect 15615 -32236 15935 -32210
rect 15615 -32864 15621 -32236
rect 15929 -32864 15935 -32236
rect 15615 -32890 15935 -32864
rect 16615 -32236 16935 -32210
rect 16615 -32864 16621 -32236
rect 16929 -32864 16935 -32236
rect 16615 -32890 16935 -32864
rect 17615 -32236 17935 -32210
rect 17615 -32864 17621 -32236
rect 17929 -32864 17935 -32236
rect 17615 -32890 17935 -32864
rect 18615 -32236 18935 -32210
rect 18615 -32864 18621 -32236
rect 18929 -32864 18935 -32236
rect 18615 -32890 18935 -32864
rect 19615 -32236 19935 -32210
rect 19615 -32864 19621 -32236
rect 19929 -32864 19935 -32236
rect 19615 -32890 19935 -32864
rect 20615 -32236 20935 -32210
rect 20615 -32864 20621 -32236
rect 20929 -32864 20935 -32236
rect 20615 -32890 20935 -32864
rect 21615 -32236 21935 -32210
rect 21615 -32864 21621 -32236
rect 21929 -32864 21935 -32236
rect 21615 -32890 21935 -32864
rect 22615 -32236 22935 -32210
rect 22615 -32864 22621 -32236
rect 22929 -32864 22935 -32236
rect 22615 -32890 22935 -32864
rect 23615 -32236 23935 -32210
rect 23615 -32864 23621 -32236
rect 23929 -32864 23935 -32236
rect 23615 -32890 23935 -32864
rect 24615 -32236 24935 -32210
rect 24615 -32864 24621 -32236
rect 24929 -32864 24935 -32236
rect 24615 -32890 24935 -32864
rect 25615 -32236 25935 -32210
rect 25615 -32864 25621 -32236
rect 25929 -32864 25935 -32236
rect 25615 -32890 25935 -32864
rect 26615 -32236 26935 -32210
rect 26615 -32864 26621 -32236
rect 26929 -32864 26935 -32236
rect 26615 -32890 26935 -32864
rect 27615 -32236 27935 -32210
rect 27615 -32864 27621 -32236
rect 27929 -32864 27935 -32236
rect 27615 -32890 27935 -32864
rect 28615 -32236 28935 -32210
rect 28615 -32864 28621 -32236
rect 28929 -32864 28935 -32236
rect 28615 -32890 28935 -32864
rect 29615 -32236 29935 -32210
rect 29615 -32864 29621 -32236
rect 29929 -32864 29935 -32236
rect 29615 -32890 29935 -32864
rect 30615 -32236 30935 -32210
rect 30615 -32864 30621 -32236
rect 30929 -32864 30935 -32236
rect 30615 -32890 30935 -32864
rect 31615 -32236 31935 -32210
rect 31615 -32864 31621 -32236
rect 31929 -32864 31935 -32236
rect 31615 -32890 31935 -32864
rect 32615 -32236 32935 -32210
rect 32615 -32864 32621 -32236
rect 32929 -32864 32935 -32236
rect 32615 -32890 32935 -32864
rect 33615 -32236 33935 -32210
rect 33615 -32864 33621 -32236
rect 33929 -32864 33935 -32236
rect 33615 -32890 33935 -32864
rect 8275 -32896 34275 -32890
rect 8275 -33204 8281 -32896
rect 8589 -32902 8961 -32896
rect 9589 -32902 9961 -32896
rect 10589 -32902 10961 -32896
rect 11589 -32902 11961 -32896
rect 12589 -32902 12961 -32896
rect 13589 -32902 13961 -32896
rect 14589 -32902 14961 -32896
rect 15589 -32902 15961 -32896
rect 16589 -32902 16961 -32896
rect 17589 -32902 17961 -32896
rect 18589 -32902 18961 -32896
rect 19589 -32902 19961 -32896
rect 20589 -32902 20961 -32896
rect 21589 -32902 21961 -32896
rect 22589 -32902 22961 -32896
rect 23589 -32902 23961 -32896
rect 24589 -32902 24961 -32896
rect 25589 -32902 25961 -32896
rect 26589 -32902 26961 -32896
rect 27589 -32902 27961 -32896
rect 28589 -32902 28961 -32896
rect 29589 -32902 29961 -32896
rect 30589 -32902 30961 -32896
rect 31589 -32902 31961 -32896
rect 32589 -32902 32961 -32896
rect 33589 -32902 33961 -32896
rect 8589 -33198 8627 -32902
rect 8923 -33198 8961 -32902
rect 9589 -33198 9627 -32902
rect 9923 -33198 9961 -32902
rect 10589 -33198 10627 -32902
rect 10923 -33198 10961 -32902
rect 11589 -33198 11627 -32902
rect 11923 -33198 11961 -32902
rect 12589 -33198 12627 -32902
rect 12923 -33198 12961 -32902
rect 13589 -33198 13627 -32902
rect 13923 -33198 13961 -32902
rect 14589 -33198 14627 -32902
rect 14923 -33198 14961 -32902
rect 15589 -33198 15627 -32902
rect 15923 -33198 15961 -32902
rect 16589 -33198 16627 -32902
rect 16923 -33198 16961 -32902
rect 17589 -33198 17627 -32902
rect 17923 -33198 17961 -32902
rect 18589 -33198 18627 -32902
rect 18923 -33198 18961 -32902
rect 19589 -33198 19627 -32902
rect 19923 -33198 19961 -32902
rect 20589 -33198 20627 -32902
rect 20923 -33198 20961 -32902
rect 21589 -33198 21627 -32902
rect 21923 -33198 21961 -32902
rect 22589 -33198 22627 -32902
rect 22923 -33198 22961 -32902
rect 23589 -33198 23627 -32902
rect 23923 -33198 23961 -32902
rect 24589 -33198 24627 -32902
rect 24923 -33198 24961 -32902
rect 25589 -33198 25627 -32902
rect 25923 -33198 25961 -32902
rect 26589 -33198 26627 -32902
rect 26923 -33198 26961 -32902
rect 27589 -33198 27627 -32902
rect 27923 -33198 27961 -32902
rect 28589 -33198 28627 -32902
rect 28923 -33198 28961 -32902
rect 29589 -33198 29627 -32902
rect 29923 -33198 29961 -32902
rect 30589 -33198 30627 -32902
rect 30923 -33198 30961 -32902
rect 31589 -33198 31627 -32902
rect 31923 -33198 31961 -32902
rect 32589 -33198 32627 -32902
rect 32923 -33198 32961 -32902
rect 33589 -33198 33627 -32902
rect 33923 -33198 33961 -32902
rect 8589 -33204 8961 -33198
rect 9589 -33204 9961 -33198
rect 10589 -33204 10961 -33198
rect 11589 -33204 11961 -33198
rect 12589 -33204 12961 -33198
rect 13589 -33204 13961 -33198
rect 14589 -33204 14961 -33198
rect 15589 -33204 15961 -33198
rect 16589 -33204 16961 -33198
rect 17589 -33204 17961 -33198
rect 18589 -33204 18961 -33198
rect 19589 -33204 19961 -33198
rect 20589 -33204 20961 -33198
rect 21589 -33204 21961 -33198
rect 22589 -33204 22961 -33198
rect 23589 -33204 23961 -33198
rect 24589 -33204 24961 -33198
rect 25589 -33204 25961 -33198
rect 26589 -33204 26961 -33198
rect 27589 -33204 27961 -33198
rect 28589 -33204 28961 -33198
rect 29589 -33204 29961 -33198
rect 30589 -33204 30961 -33198
rect 31589 -33204 31961 -33198
rect 32589 -33204 32961 -33198
rect 33589 -33204 33961 -33198
rect 34269 -33204 34275 -32896
rect 8275 -33210 34275 -33204
rect 8615 -33236 8935 -33210
rect 8615 -33864 8621 -33236
rect 8929 -33864 8935 -33236
rect 8615 -33890 8935 -33864
rect 9615 -33236 9935 -33210
rect 9615 -33864 9621 -33236
rect 9929 -33864 9935 -33236
rect 9615 -33890 9935 -33864
rect 10615 -33236 10935 -33210
rect 10615 -33864 10621 -33236
rect 10929 -33864 10935 -33236
rect 10615 -33890 10935 -33864
rect 11615 -33236 11935 -33210
rect 11615 -33864 11621 -33236
rect 11929 -33864 11935 -33236
rect 11615 -33890 11935 -33864
rect 12615 -33236 12935 -33210
rect 12615 -33864 12621 -33236
rect 12929 -33864 12935 -33236
rect 12615 -33890 12935 -33864
rect 13615 -33236 13935 -33210
rect 13615 -33864 13621 -33236
rect 13929 -33864 13935 -33236
rect 13615 -33890 13935 -33864
rect 14615 -33236 14935 -33210
rect 14615 -33864 14621 -33236
rect 14929 -33864 14935 -33236
rect 14615 -33890 14935 -33864
rect 15615 -33236 15935 -33210
rect 15615 -33864 15621 -33236
rect 15929 -33864 15935 -33236
rect 15615 -33890 15935 -33864
rect 16615 -33236 16935 -33210
rect 16615 -33864 16621 -33236
rect 16929 -33864 16935 -33236
rect 16615 -33890 16935 -33864
rect 17615 -33236 17935 -33210
rect 17615 -33864 17621 -33236
rect 17929 -33864 17935 -33236
rect 17615 -33890 17935 -33864
rect 18615 -33236 18935 -33210
rect 18615 -33864 18621 -33236
rect 18929 -33864 18935 -33236
rect 18615 -33890 18935 -33864
rect 19615 -33236 19935 -33210
rect 19615 -33864 19621 -33236
rect 19929 -33864 19935 -33236
rect 19615 -33890 19935 -33864
rect 20615 -33236 20935 -33210
rect 20615 -33864 20621 -33236
rect 20929 -33864 20935 -33236
rect 20615 -33890 20935 -33864
rect 21615 -33236 21935 -33210
rect 21615 -33864 21621 -33236
rect 21929 -33864 21935 -33236
rect 21615 -33890 21935 -33864
rect 22615 -33236 22935 -33210
rect 22615 -33864 22621 -33236
rect 22929 -33864 22935 -33236
rect 22615 -33890 22935 -33864
rect 23615 -33236 23935 -33210
rect 23615 -33864 23621 -33236
rect 23929 -33864 23935 -33236
rect 23615 -33890 23935 -33864
rect 24615 -33236 24935 -33210
rect 24615 -33864 24621 -33236
rect 24929 -33864 24935 -33236
rect 24615 -33890 24935 -33864
rect 25615 -33236 25935 -33210
rect 25615 -33864 25621 -33236
rect 25929 -33864 25935 -33236
rect 25615 -33890 25935 -33864
rect 26615 -33236 26935 -33210
rect 26615 -33864 26621 -33236
rect 26929 -33864 26935 -33236
rect 26615 -33890 26935 -33864
rect 27615 -33236 27935 -33210
rect 27615 -33864 27621 -33236
rect 27929 -33864 27935 -33236
rect 27615 -33890 27935 -33864
rect 28615 -33236 28935 -33210
rect 28615 -33864 28621 -33236
rect 28929 -33864 28935 -33236
rect 28615 -33890 28935 -33864
rect 29615 -33236 29935 -33210
rect 29615 -33864 29621 -33236
rect 29929 -33864 29935 -33236
rect 29615 -33890 29935 -33864
rect 30615 -33236 30935 -33210
rect 30615 -33864 30621 -33236
rect 30929 -33864 30935 -33236
rect 30615 -33890 30935 -33864
rect 31615 -33236 31935 -33210
rect 31615 -33864 31621 -33236
rect 31929 -33864 31935 -33236
rect 31615 -33890 31935 -33864
rect 32615 -33236 32935 -33210
rect 32615 -33864 32621 -33236
rect 32929 -33864 32935 -33236
rect 32615 -33890 32935 -33864
rect 33615 -33236 33935 -33210
rect 33615 -33864 33621 -33236
rect 33929 -33864 33935 -33236
rect 33615 -33890 33935 -33864
rect 8275 -33896 34275 -33890
rect 8275 -34204 8281 -33896
rect 8589 -33902 8961 -33896
rect 9589 -33902 9961 -33896
rect 10589 -33902 10961 -33896
rect 11589 -33902 11961 -33896
rect 12589 -33902 12961 -33896
rect 13589 -33902 13961 -33896
rect 14589 -33902 14961 -33896
rect 15589 -33902 15961 -33896
rect 16589 -33902 16961 -33896
rect 17589 -33902 17961 -33896
rect 18589 -33902 18961 -33896
rect 19589 -33902 19961 -33896
rect 20589 -33902 20961 -33896
rect 21589 -33902 21961 -33896
rect 22589 -33902 22961 -33896
rect 23589 -33902 23961 -33896
rect 24589 -33902 24961 -33896
rect 25589 -33902 25961 -33896
rect 26589 -33902 26961 -33896
rect 27589 -33902 27961 -33896
rect 28589 -33902 28961 -33896
rect 29589 -33902 29961 -33896
rect 30589 -33902 30961 -33896
rect 31589 -33902 31961 -33896
rect 32589 -33902 32961 -33896
rect 33589 -33902 33961 -33896
rect 8589 -34198 8627 -33902
rect 8923 -34198 8961 -33902
rect 9589 -34198 9627 -33902
rect 9923 -34198 9961 -33902
rect 10589 -34198 10627 -33902
rect 10923 -34198 10961 -33902
rect 11589 -34198 11627 -33902
rect 11923 -34198 11961 -33902
rect 12589 -34198 12627 -33902
rect 12923 -34198 12961 -33902
rect 13589 -34198 13627 -33902
rect 13923 -34198 13961 -33902
rect 14589 -34198 14627 -33902
rect 14923 -34198 14961 -33902
rect 15589 -34198 15627 -33902
rect 15923 -34198 15961 -33902
rect 16589 -34198 16627 -33902
rect 16923 -34198 16961 -33902
rect 17589 -34198 17627 -33902
rect 17923 -34198 17961 -33902
rect 18589 -34198 18627 -33902
rect 18923 -34198 18961 -33902
rect 19589 -34198 19627 -33902
rect 19923 -34198 19961 -33902
rect 20589 -34198 20627 -33902
rect 20923 -34198 20961 -33902
rect 21589 -34198 21627 -33902
rect 21923 -34198 21961 -33902
rect 22589 -34198 22627 -33902
rect 22923 -34198 22961 -33902
rect 23589 -34198 23627 -33902
rect 23923 -34198 23961 -33902
rect 24589 -34198 24627 -33902
rect 24923 -34198 24961 -33902
rect 25589 -34198 25627 -33902
rect 25923 -34198 25961 -33902
rect 26589 -34198 26627 -33902
rect 26923 -34198 26961 -33902
rect 27589 -34198 27627 -33902
rect 27923 -34198 27961 -33902
rect 28589 -34198 28627 -33902
rect 28923 -34198 28961 -33902
rect 29589 -34198 29627 -33902
rect 29923 -34198 29961 -33902
rect 30589 -34198 30627 -33902
rect 30923 -34198 30961 -33902
rect 31589 -34198 31627 -33902
rect 31923 -34198 31961 -33902
rect 32589 -34198 32627 -33902
rect 32923 -34198 32961 -33902
rect 33589 -34198 33627 -33902
rect 33923 -34198 33961 -33902
rect 8589 -34204 8961 -34198
rect 9589 -34204 9961 -34198
rect 10589 -34204 10961 -34198
rect 11589 -34204 11961 -34198
rect 12589 -34204 12961 -34198
rect 13589 -34204 13961 -34198
rect 14589 -34204 14961 -34198
rect 15589 -34204 15961 -34198
rect 16589 -34204 16961 -34198
rect 17589 -34204 17961 -34198
rect 18589 -34204 18961 -34198
rect 19589 -34204 19961 -34198
rect 20589 -34204 20961 -34198
rect 21589 -34204 21961 -34198
rect 22589 -34204 22961 -34198
rect 23589 -34204 23961 -34198
rect 24589 -34204 24961 -34198
rect 25589 -34204 25961 -34198
rect 26589 -34204 26961 -34198
rect 27589 -34204 27961 -34198
rect 28589 -34204 28961 -34198
rect 29589 -34204 29961 -34198
rect 30589 -34204 30961 -34198
rect 31589 -34204 31961 -34198
rect 32589 -34204 32961 -34198
rect 33589 -34204 33961 -34198
rect 34269 -34204 34275 -33896
rect 8275 -34210 34275 -34204
rect 8615 -34236 8935 -34210
rect 8615 -34864 8621 -34236
rect 8929 -34864 8935 -34236
rect 8615 -34890 8935 -34864
rect 9615 -34236 9935 -34210
rect 9615 -34864 9621 -34236
rect 9929 -34864 9935 -34236
rect 9615 -34890 9935 -34864
rect 10615 -34236 10935 -34210
rect 10615 -34864 10621 -34236
rect 10929 -34864 10935 -34236
rect 10615 -34890 10935 -34864
rect 11615 -34236 11935 -34210
rect 11615 -34864 11621 -34236
rect 11929 -34864 11935 -34236
rect 11615 -34890 11935 -34864
rect 12615 -34236 12935 -34210
rect 12615 -34864 12621 -34236
rect 12929 -34864 12935 -34236
rect 12615 -34890 12935 -34864
rect 13615 -34236 13935 -34210
rect 13615 -34864 13621 -34236
rect 13929 -34864 13935 -34236
rect 13615 -34890 13935 -34864
rect 14615 -34236 14935 -34210
rect 14615 -34864 14621 -34236
rect 14929 -34864 14935 -34236
rect 14615 -34890 14935 -34864
rect 15615 -34236 15935 -34210
rect 15615 -34864 15621 -34236
rect 15929 -34864 15935 -34236
rect 15615 -34890 15935 -34864
rect 16615 -34236 16935 -34210
rect 16615 -34864 16621 -34236
rect 16929 -34864 16935 -34236
rect 16615 -34890 16935 -34864
rect 17615 -34236 17935 -34210
rect 17615 -34864 17621 -34236
rect 17929 -34864 17935 -34236
rect 17615 -34890 17935 -34864
rect 18615 -34236 18935 -34210
rect 18615 -34864 18621 -34236
rect 18929 -34864 18935 -34236
rect 18615 -34890 18935 -34864
rect 19615 -34236 19935 -34210
rect 19615 -34864 19621 -34236
rect 19929 -34864 19935 -34236
rect 19615 -34890 19935 -34864
rect 20615 -34236 20935 -34210
rect 20615 -34864 20621 -34236
rect 20929 -34864 20935 -34236
rect 20615 -34890 20935 -34864
rect 21615 -34236 21935 -34210
rect 21615 -34864 21621 -34236
rect 21929 -34864 21935 -34236
rect 21615 -34890 21935 -34864
rect 22615 -34236 22935 -34210
rect 22615 -34864 22621 -34236
rect 22929 -34864 22935 -34236
rect 22615 -34890 22935 -34864
rect 23615 -34236 23935 -34210
rect 23615 -34864 23621 -34236
rect 23929 -34864 23935 -34236
rect 23615 -34890 23935 -34864
rect 24615 -34236 24935 -34210
rect 24615 -34864 24621 -34236
rect 24929 -34864 24935 -34236
rect 24615 -34890 24935 -34864
rect 25615 -34236 25935 -34210
rect 25615 -34864 25621 -34236
rect 25929 -34864 25935 -34236
rect 25615 -34890 25935 -34864
rect 26615 -34236 26935 -34210
rect 26615 -34864 26621 -34236
rect 26929 -34864 26935 -34236
rect 26615 -34890 26935 -34864
rect 27615 -34236 27935 -34210
rect 27615 -34864 27621 -34236
rect 27929 -34864 27935 -34236
rect 27615 -34890 27935 -34864
rect 28615 -34236 28935 -34210
rect 28615 -34864 28621 -34236
rect 28929 -34864 28935 -34236
rect 28615 -34890 28935 -34864
rect 29615 -34236 29935 -34210
rect 29615 -34864 29621 -34236
rect 29929 -34864 29935 -34236
rect 29615 -34890 29935 -34864
rect 30615 -34236 30935 -34210
rect 30615 -34864 30621 -34236
rect 30929 -34864 30935 -34236
rect 30615 -34890 30935 -34864
rect 31615 -34236 31935 -34210
rect 31615 -34864 31621 -34236
rect 31929 -34864 31935 -34236
rect 31615 -34890 31935 -34864
rect 32615 -34236 32935 -34210
rect 32615 -34864 32621 -34236
rect 32929 -34864 32935 -34236
rect 32615 -34890 32935 -34864
rect 33615 -34236 33935 -34210
rect 33615 -34864 33621 -34236
rect 33929 -34864 33935 -34236
rect 33615 -34890 33935 -34864
rect 8275 -34896 34275 -34890
rect 8275 -35204 8281 -34896
rect 8589 -34902 8961 -34896
rect 9589 -34902 9961 -34896
rect 10589 -34902 10961 -34896
rect 11589 -34902 11961 -34896
rect 12589 -34902 12961 -34896
rect 13589 -34902 13961 -34896
rect 14589 -34902 14961 -34896
rect 15589 -34902 15961 -34896
rect 16589 -34902 16961 -34896
rect 17589 -34902 17961 -34896
rect 18589 -34902 18961 -34896
rect 19589 -34902 19961 -34896
rect 20589 -34902 20961 -34896
rect 21589 -34902 21961 -34896
rect 22589 -34902 22961 -34896
rect 23589 -34902 23961 -34896
rect 24589 -34902 24961 -34896
rect 25589 -34902 25961 -34896
rect 26589 -34902 26961 -34896
rect 27589 -34902 27961 -34896
rect 28589 -34902 28961 -34896
rect 29589 -34902 29961 -34896
rect 30589 -34902 30961 -34896
rect 31589 -34902 31961 -34896
rect 32589 -34902 32961 -34896
rect 33589 -34902 33961 -34896
rect 8589 -35198 8627 -34902
rect 8923 -35198 8961 -34902
rect 9589 -35198 9627 -34902
rect 9923 -35198 9961 -34902
rect 10589 -35198 10627 -34902
rect 10923 -35198 10961 -34902
rect 11589 -35198 11627 -34902
rect 11923 -35198 11961 -34902
rect 12589 -35198 12627 -34902
rect 12923 -35198 12961 -34902
rect 13589 -35198 13627 -34902
rect 13923 -35198 13961 -34902
rect 14589 -35198 14627 -34902
rect 14923 -35198 14961 -34902
rect 15589 -35198 15627 -34902
rect 15923 -35198 15961 -34902
rect 16589 -35198 16627 -34902
rect 16923 -35198 16961 -34902
rect 17589 -35198 17627 -34902
rect 17923 -35198 17961 -34902
rect 18589 -35198 18627 -34902
rect 18923 -35198 18961 -34902
rect 19589 -35198 19627 -34902
rect 19923 -35198 19961 -34902
rect 20589 -35198 20627 -34902
rect 20923 -35198 20961 -34902
rect 21589 -35198 21627 -34902
rect 21923 -35198 21961 -34902
rect 22589 -35198 22627 -34902
rect 22923 -35198 22961 -34902
rect 23589 -35198 23627 -34902
rect 23923 -35198 23961 -34902
rect 24589 -35198 24627 -34902
rect 24923 -35198 24961 -34902
rect 25589 -35198 25627 -34902
rect 25923 -35198 25961 -34902
rect 26589 -35198 26627 -34902
rect 26923 -35198 26961 -34902
rect 27589 -35198 27627 -34902
rect 27923 -35198 27961 -34902
rect 28589 -35198 28627 -34902
rect 28923 -35198 28961 -34902
rect 29589 -35198 29627 -34902
rect 29923 -35198 29961 -34902
rect 30589 -35198 30627 -34902
rect 30923 -35198 30961 -34902
rect 31589 -35198 31627 -34902
rect 31923 -35198 31961 -34902
rect 32589 -35198 32627 -34902
rect 32923 -35198 32961 -34902
rect 33589 -35198 33627 -34902
rect 33923 -35198 33961 -34902
rect 8589 -35204 8961 -35198
rect 9589 -35204 9961 -35198
rect 10589 -35204 10961 -35198
rect 11589 -35204 11961 -35198
rect 12589 -35204 12961 -35198
rect 13589 -35204 13961 -35198
rect 14589 -35204 14961 -35198
rect 15589 -35204 15961 -35198
rect 16589 -35204 16961 -35198
rect 17589 -35204 17961 -35198
rect 18589 -35204 18961 -35198
rect 19589 -35204 19961 -35198
rect 20589 -35204 20961 -35198
rect 21589 -35204 21961 -35198
rect 22589 -35204 22961 -35198
rect 23589 -35204 23961 -35198
rect 24589 -35204 24961 -35198
rect 25589 -35204 25961 -35198
rect 26589 -35204 26961 -35198
rect 27589 -35204 27961 -35198
rect 28589 -35204 28961 -35198
rect 29589 -35204 29961 -35198
rect 30589 -35204 30961 -35198
rect 31589 -35204 31961 -35198
rect 32589 -35204 32961 -35198
rect 33589 -35204 33961 -35198
rect 34269 -35204 34275 -34896
rect 8275 -35210 34275 -35204
rect 8615 -35236 8935 -35210
rect 8615 -35864 8621 -35236
rect 8929 -35864 8935 -35236
rect 8615 -35890 8935 -35864
rect 9615 -35236 9935 -35210
rect 9615 -35864 9621 -35236
rect 9929 -35864 9935 -35236
rect 9615 -35890 9935 -35864
rect 10615 -35236 10935 -35210
rect 10615 -35864 10621 -35236
rect 10929 -35864 10935 -35236
rect 10615 -35890 10935 -35864
rect 11615 -35236 11935 -35210
rect 11615 -35864 11621 -35236
rect 11929 -35864 11935 -35236
rect 11615 -35890 11935 -35864
rect 12615 -35236 12935 -35210
rect 12615 -35864 12621 -35236
rect 12929 -35864 12935 -35236
rect 12615 -35890 12935 -35864
rect 13615 -35236 13935 -35210
rect 13615 -35864 13621 -35236
rect 13929 -35864 13935 -35236
rect 13615 -35890 13935 -35864
rect 14615 -35236 14935 -35210
rect 14615 -35864 14621 -35236
rect 14929 -35864 14935 -35236
rect 14615 -35890 14935 -35864
rect 15615 -35236 15935 -35210
rect 15615 -35864 15621 -35236
rect 15929 -35864 15935 -35236
rect 15615 -35890 15935 -35864
rect 16615 -35236 16935 -35210
rect 16615 -35864 16621 -35236
rect 16929 -35864 16935 -35236
rect 16615 -35890 16935 -35864
rect 17615 -35236 17935 -35210
rect 17615 -35864 17621 -35236
rect 17929 -35864 17935 -35236
rect 17615 -35890 17935 -35864
rect 18615 -35236 18935 -35210
rect 18615 -35864 18621 -35236
rect 18929 -35864 18935 -35236
rect 18615 -35890 18935 -35864
rect 19615 -35236 19935 -35210
rect 19615 -35864 19621 -35236
rect 19929 -35864 19935 -35236
rect 19615 -35890 19935 -35864
rect 20615 -35236 20935 -35210
rect 20615 -35864 20621 -35236
rect 20929 -35864 20935 -35236
rect 20615 -35890 20935 -35864
rect 21615 -35236 21935 -35210
rect 21615 -35864 21621 -35236
rect 21929 -35864 21935 -35236
rect 21615 -35890 21935 -35864
rect 22615 -35236 22935 -35210
rect 22615 -35864 22621 -35236
rect 22929 -35864 22935 -35236
rect 22615 -35890 22935 -35864
rect 23615 -35236 23935 -35210
rect 23615 -35864 23621 -35236
rect 23929 -35864 23935 -35236
rect 23615 -35890 23935 -35864
rect 24615 -35236 24935 -35210
rect 24615 -35864 24621 -35236
rect 24929 -35864 24935 -35236
rect 24615 -35890 24935 -35864
rect 25615 -35236 25935 -35210
rect 25615 -35864 25621 -35236
rect 25929 -35864 25935 -35236
rect 25615 -35890 25935 -35864
rect 26615 -35236 26935 -35210
rect 26615 -35864 26621 -35236
rect 26929 -35864 26935 -35236
rect 26615 -35890 26935 -35864
rect 27615 -35236 27935 -35210
rect 27615 -35864 27621 -35236
rect 27929 -35864 27935 -35236
rect 27615 -35890 27935 -35864
rect 28615 -35236 28935 -35210
rect 28615 -35864 28621 -35236
rect 28929 -35864 28935 -35236
rect 28615 -35890 28935 -35864
rect 29615 -35236 29935 -35210
rect 29615 -35864 29621 -35236
rect 29929 -35864 29935 -35236
rect 29615 -35890 29935 -35864
rect 30615 -35236 30935 -35210
rect 30615 -35864 30621 -35236
rect 30929 -35864 30935 -35236
rect 30615 -35890 30935 -35864
rect 31615 -35236 31935 -35210
rect 31615 -35864 31621 -35236
rect 31929 -35864 31935 -35236
rect 31615 -35890 31935 -35864
rect 32615 -35236 32935 -35210
rect 32615 -35864 32621 -35236
rect 32929 -35864 32935 -35236
rect 32615 -35890 32935 -35864
rect 33615 -35236 33935 -35210
rect 33615 -35864 33621 -35236
rect 33929 -35864 33935 -35236
rect 33615 -35890 33935 -35864
rect 8275 -35896 34275 -35890
rect 8275 -36204 8281 -35896
rect 8589 -35902 8961 -35896
rect 9589 -35902 9961 -35896
rect 10589 -35902 10961 -35896
rect 11589 -35902 11961 -35896
rect 12589 -35902 12961 -35896
rect 13589 -35902 13961 -35896
rect 14589 -35902 14961 -35896
rect 15589 -35902 15961 -35896
rect 16589 -35902 16961 -35896
rect 17589 -35902 17961 -35896
rect 18589 -35902 18961 -35896
rect 19589 -35902 19961 -35896
rect 20589 -35902 20961 -35896
rect 21589 -35902 21961 -35896
rect 22589 -35902 22961 -35896
rect 23589 -35902 23961 -35896
rect 24589 -35902 24961 -35896
rect 25589 -35902 25961 -35896
rect 26589 -35902 26961 -35896
rect 27589 -35902 27961 -35896
rect 28589 -35902 28961 -35896
rect 29589 -35902 29961 -35896
rect 30589 -35902 30961 -35896
rect 31589 -35902 31961 -35896
rect 32589 -35902 32961 -35896
rect 33589 -35902 33961 -35896
rect 8589 -36198 8627 -35902
rect 8923 -36198 8961 -35902
rect 9589 -36198 9627 -35902
rect 9923 -36198 9961 -35902
rect 10589 -36198 10627 -35902
rect 10923 -36198 10961 -35902
rect 11589 -36198 11627 -35902
rect 11923 -36198 11961 -35902
rect 12589 -36198 12627 -35902
rect 12923 -36198 12961 -35902
rect 13589 -36198 13627 -35902
rect 13923 -36198 13961 -35902
rect 14589 -36198 14627 -35902
rect 14923 -36198 14961 -35902
rect 15589 -36198 15627 -35902
rect 15923 -36198 15961 -35902
rect 16589 -36198 16627 -35902
rect 16923 -36198 16961 -35902
rect 17589 -36198 17627 -35902
rect 17923 -36198 17961 -35902
rect 18589 -36198 18627 -35902
rect 18923 -36198 18961 -35902
rect 19589 -36198 19627 -35902
rect 19923 -36198 19961 -35902
rect 20589 -36198 20627 -35902
rect 20923 -36198 20961 -35902
rect 21589 -36198 21627 -35902
rect 21923 -36198 21961 -35902
rect 22589 -36198 22627 -35902
rect 22923 -36198 22961 -35902
rect 23589 -36198 23627 -35902
rect 23923 -36198 23961 -35902
rect 24589 -36198 24627 -35902
rect 24923 -36198 24961 -35902
rect 25589 -36198 25627 -35902
rect 25923 -36198 25961 -35902
rect 26589 -36198 26627 -35902
rect 26923 -36198 26961 -35902
rect 27589 -36198 27627 -35902
rect 27923 -36198 27961 -35902
rect 28589 -36198 28627 -35902
rect 28923 -36198 28961 -35902
rect 29589 -36198 29627 -35902
rect 29923 -36198 29961 -35902
rect 30589 -36198 30627 -35902
rect 30923 -36198 30961 -35902
rect 31589 -36198 31627 -35902
rect 31923 -36198 31961 -35902
rect 32589 -36198 32627 -35902
rect 32923 -36198 32961 -35902
rect 33589 -36198 33627 -35902
rect 33923 -36198 33961 -35902
rect 8589 -36204 8961 -36198
rect 9589 -36204 9961 -36198
rect 10589 -36204 10961 -36198
rect 11589 -36204 11961 -36198
rect 12589 -36204 12961 -36198
rect 13589 -36204 13961 -36198
rect 14589 -36204 14961 -36198
rect 15589 -36204 15961 -36198
rect 16589 -36204 16961 -36198
rect 17589 -36204 17961 -36198
rect 18589 -36204 18961 -36198
rect 19589 -36204 19961 -36198
rect 20589 -36204 20961 -36198
rect 21589 -36204 21961 -36198
rect 22589 -36204 22961 -36198
rect 23589 -36204 23961 -36198
rect 24589 -36204 24961 -36198
rect 25589 -36204 25961 -36198
rect 26589 -36204 26961 -36198
rect 27589 -36204 27961 -36198
rect 28589 -36204 28961 -36198
rect 29589 -36204 29961 -36198
rect 30589 -36204 30961 -36198
rect 31589 -36204 31961 -36198
rect 32589 -36204 32961 -36198
rect 33589 -36204 33961 -36198
rect 34269 -36204 34275 -35896
rect 8275 -36210 34275 -36204
rect 8615 -36236 8935 -36210
rect 8615 -36864 8621 -36236
rect 8929 -36864 8935 -36236
rect 8615 -36890 8935 -36864
rect 9615 -36236 9935 -36210
rect 9615 -36864 9621 -36236
rect 9929 -36864 9935 -36236
rect 9615 -36890 9935 -36864
rect 10615 -36236 10935 -36210
rect 10615 -36864 10621 -36236
rect 10929 -36864 10935 -36236
rect 10615 -36890 10935 -36864
rect 11615 -36236 11935 -36210
rect 11615 -36864 11621 -36236
rect 11929 -36864 11935 -36236
rect 11615 -36890 11935 -36864
rect 12615 -36236 12935 -36210
rect 12615 -36864 12621 -36236
rect 12929 -36864 12935 -36236
rect 12615 -36890 12935 -36864
rect 13615 -36236 13935 -36210
rect 13615 -36864 13621 -36236
rect 13929 -36864 13935 -36236
rect 13615 -36890 13935 -36864
rect 14615 -36236 14935 -36210
rect 14615 -36864 14621 -36236
rect 14929 -36864 14935 -36236
rect 14615 -36890 14935 -36864
rect 15615 -36236 15935 -36210
rect 15615 -36864 15621 -36236
rect 15929 -36864 15935 -36236
rect 15615 -36890 15935 -36864
rect 16615 -36236 16935 -36210
rect 16615 -36864 16621 -36236
rect 16929 -36864 16935 -36236
rect 16615 -36890 16935 -36864
rect 17615 -36236 17935 -36210
rect 17615 -36864 17621 -36236
rect 17929 -36864 17935 -36236
rect 17615 -36890 17935 -36864
rect 18615 -36236 18935 -36210
rect 18615 -36864 18621 -36236
rect 18929 -36864 18935 -36236
rect 18615 -36890 18935 -36864
rect 19615 -36236 19935 -36210
rect 19615 -36864 19621 -36236
rect 19929 -36864 19935 -36236
rect 19615 -36890 19935 -36864
rect 20615 -36236 20935 -36210
rect 20615 -36864 20621 -36236
rect 20929 -36864 20935 -36236
rect 20615 -36890 20935 -36864
rect 21615 -36236 21935 -36210
rect 21615 -36864 21621 -36236
rect 21929 -36864 21935 -36236
rect 21615 -36890 21935 -36864
rect 22615 -36236 22935 -36210
rect 22615 -36864 22621 -36236
rect 22929 -36864 22935 -36236
rect 22615 -36890 22935 -36864
rect 23615 -36236 23935 -36210
rect 23615 -36864 23621 -36236
rect 23929 -36864 23935 -36236
rect 23615 -36890 23935 -36864
rect 24615 -36236 24935 -36210
rect 24615 -36864 24621 -36236
rect 24929 -36864 24935 -36236
rect 24615 -36890 24935 -36864
rect 25615 -36236 25935 -36210
rect 25615 -36864 25621 -36236
rect 25929 -36864 25935 -36236
rect 25615 -36890 25935 -36864
rect 26615 -36236 26935 -36210
rect 26615 -36864 26621 -36236
rect 26929 -36864 26935 -36236
rect 26615 -36890 26935 -36864
rect 27615 -36236 27935 -36210
rect 27615 -36864 27621 -36236
rect 27929 -36864 27935 -36236
rect 27615 -36890 27935 -36864
rect 28615 -36236 28935 -36210
rect 28615 -36864 28621 -36236
rect 28929 -36864 28935 -36236
rect 28615 -36890 28935 -36864
rect 29615 -36236 29935 -36210
rect 29615 -36864 29621 -36236
rect 29929 -36864 29935 -36236
rect 29615 -36890 29935 -36864
rect 30615 -36236 30935 -36210
rect 30615 -36864 30621 -36236
rect 30929 -36864 30935 -36236
rect 30615 -36890 30935 -36864
rect 31615 -36236 31935 -36210
rect 31615 -36864 31621 -36236
rect 31929 -36864 31935 -36236
rect 31615 -36890 31935 -36864
rect 32615 -36236 32935 -36210
rect 32615 -36864 32621 -36236
rect 32929 -36864 32935 -36236
rect 32615 -36890 32935 -36864
rect 33615 -36236 33935 -36210
rect 33615 -36864 33621 -36236
rect 33929 -36864 33935 -36236
rect 33615 -36890 33935 -36864
rect 8275 -36896 34275 -36890
rect 8275 -37204 8281 -36896
rect 8589 -36902 8961 -36896
rect 9589 -36902 9961 -36896
rect 10589 -36902 10961 -36896
rect 11589 -36902 11961 -36896
rect 12589 -36902 12961 -36896
rect 13589 -36902 13961 -36896
rect 14589 -36902 14961 -36896
rect 15589 -36902 15961 -36896
rect 16589 -36902 16961 -36896
rect 17589 -36902 17961 -36896
rect 18589 -36902 18961 -36896
rect 19589 -36902 19961 -36896
rect 20589 -36902 20961 -36896
rect 21589 -36902 21961 -36896
rect 22589 -36902 22961 -36896
rect 23589 -36902 23961 -36896
rect 24589 -36902 24961 -36896
rect 25589 -36902 25961 -36896
rect 26589 -36902 26961 -36896
rect 27589 -36902 27961 -36896
rect 28589 -36902 28961 -36896
rect 29589 -36902 29961 -36896
rect 30589 -36902 30961 -36896
rect 31589 -36902 31961 -36896
rect 32589 -36902 32961 -36896
rect 33589 -36902 33961 -36896
rect 8589 -37198 8627 -36902
rect 8923 -37198 8961 -36902
rect 9589 -37198 9627 -36902
rect 9923 -37198 9961 -36902
rect 10589 -37198 10627 -36902
rect 10923 -37198 10961 -36902
rect 11589 -37198 11627 -36902
rect 11923 -37198 11961 -36902
rect 12589 -37198 12627 -36902
rect 12923 -37198 12961 -36902
rect 13589 -37198 13627 -36902
rect 13923 -37198 13961 -36902
rect 14589 -37198 14627 -36902
rect 14923 -37198 14961 -36902
rect 15589 -37198 15627 -36902
rect 15923 -37198 15961 -36902
rect 16589 -37198 16627 -36902
rect 16923 -37198 16961 -36902
rect 17589 -37198 17627 -36902
rect 17923 -37198 17961 -36902
rect 18589 -37198 18627 -36902
rect 18923 -37198 18961 -36902
rect 19589 -37198 19627 -36902
rect 19923 -37198 19961 -36902
rect 20589 -37198 20627 -36902
rect 20923 -37198 20961 -36902
rect 21589 -37198 21627 -36902
rect 21923 -37198 21961 -36902
rect 22589 -37198 22627 -36902
rect 22923 -37198 22961 -36902
rect 23589 -37198 23627 -36902
rect 23923 -37198 23961 -36902
rect 24589 -37198 24627 -36902
rect 24923 -37198 24961 -36902
rect 25589 -37198 25627 -36902
rect 25923 -37198 25961 -36902
rect 26589 -37198 26627 -36902
rect 26923 -37198 26961 -36902
rect 27589 -37198 27627 -36902
rect 27923 -37198 27961 -36902
rect 28589 -37198 28627 -36902
rect 28923 -37198 28961 -36902
rect 29589 -37198 29627 -36902
rect 29923 -37198 29961 -36902
rect 30589 -37198 30627 -36902
rect 30923 -37198 30961 -36902
rect 31589 -37198 31627 -36902
rect 31923 -37198 31961 -36902
rect 32589 -37198 32627 -36902
rect 32923 -37198 32961 -36902
rect 33589 -37198 33627 -36902
rect 33923 -37198 33961 -36902
rect 8589 -37204 8961 -37198
rect 9589 -37204 9961 -37198
rect 10589 -37204 10961 -37198
rect 11589 -37204 11961 -37198
rect 12589 -37204 12961 -37198
rect 13589 -37204 13961 -37198
rect 14589 -37204 14961 -37198
rect 15589 -37204 15961 -37198
rect 16589 -37204 16961 -37198
rect 17589 -37204 17961 -37198
rect 18589 -37204 18961 -37198
rect 19589 -37204 19961 -37198
rect 20589 -37204 20961 -37198
rect 21589 -37204 21961 -37198
rect 22589 -37204 22961 -37198
rect 23589 -37204 23961 -37198
rect 24589 -37204 24961 -37198
rect 25589 -37204 25961 -37198
rect 26589 -37204 26961 -37198
rect 27589 -37204 27961 -37198
rect 28589 -37204 28961 -37198
rect 29589 -37204 29961 -37198
rect 30589 -37204 30961 -37198
rect 31589 -37204 31961 -37198
rect 32589 -37204 32961 -37198
rect 33589 -37204 33961 -37198
rect 34269 -37204 34275 -36896
rect 8275 -37210 34275 -37204
rect 8615 -37236 8935 -37210
rect 8615 -37864 8621 -37236
rect 8929 -37864 8935 -37236
rect 8615 -37890 8935 -37864
rect 9615 -37236 9935 -37210
rect 9615 -37864 9621 -37236
rect 9929 -37864 9935 -37236
rect 9615 -37890 9935 -37864
rect 10615 -37236 10935 -37210
rect 10615 -37864 10621 -37236
rect 10929 -37864 10935 -37236
rect 10615 -37890 10935 -37864
rect 11615 -37236 11935 -37210
rect 11615 -37864 11621 -37236
rect 11929 -37864 11935 -37236
rect 11615 -37890 11935 -37864
rect 12615 -37236 12935 -37210
rect 12615 -37864 12621 -37236
rect 12929 -37864 12935 -37236
rect 12615 -37890 12935 -37864
rect 13615 -37236 13935 -37210
rect 13615 -37864 13621 -37236
rect 13929 -37864 13935 -37236
rect 13615 -37890 13935 -37864
rect 14615 -37236 14935 -37210
rect 14615 -37864 14621 -37236
rect 14929 -37864 14935 -37236
rect 14615 -37890 14935 -37864
rect 15615 -37236 15935 -37210
rect 15615 -37864 15621 -37236
rect 15929 -37864 15935 -37236
rect 15615 -37890 15935 -37864
rect 16615 -37236 16935 -37210
rect 16615 -37864 16621 -37236
rect 16929 -37864 16935 -37236
rect 16615 -37890 16935 -37864
rect 17615 -37236 17935 -37210
rect 17615 -37864 17621 -37236
rect 17929 -37864 17935 -37236
rect 17615 -37890 17935 -37864
rect 18615 -37236 18935 -37210
rect 18615 -37864 18621 -37236
rect 18929 -37864 18935 -37236
rect 18615 -37890 18935 -37864
rect 19615 -37236 19935 -37210
rect 19615 -37864 19621 -37236
rect 19929 -37864 19935 -37236
rect 19615 -37890 19935 -37864
rect 20615 -37236 20935 -37210
rect 20615 -37864 20621 -37236
rect 20929 -37864 20935 -37236
rect 20615 -37890 20935 -37864
rect 21615 -37236 21935 -37210
rect 21615 -37864 21621 -37236
rect 21929 -37864 21935 -37236
rect 21615 -37890 21935 -37864
rect 22615 -37236 22935 -37210
rect 22615 -37864 22621 -37236
rect 22929 -37864 22935 -37236
rect 22615 -37890 22935 -37864
rect 23615 -37236 23935 -37210
rect 23615 -37864 23621 -37236
rect 23929 -37864 23935 -37236
rect 23615 -37890 23935 -37864
rect 24615 -37236 24935 -37210
rect 24615 -37864 24621 -37236
rect 24929 -37864 24935 -37236
rect 24615 -37890 24935 -37864
rect 25615 -37236 25935 -37210
rect 25615 -37864 25621 -37236
rect 25929 -37864 25935 -37236
rect 25615 -37890 25935 -37864
rect 26615 -37236 26935 -37210
rect 26615 -37864 26621 -37236
rect 26929 -37864 26935 -37236
rect 26615 -37890 26935 -37864
rect 27615 -37236 27935 -37210
rect 27615 -37864 27621 -37236
rect 27929 -37864 27935 -37236
rect 27615 -37890 27935 -37864
rect 28615 -37236 28935 -37210
rect 28615 -37864 28621 -37236
rect 28929 -37864 28935 -37236
rect 28615 -37890 28935 -37864
rect 29615 -37236 29935 -37210
rect 29615 -37864 29621 -37236
rect 29929 -37864 29935 -37236
rect 29615 -37890 29935 -37864
rect 30615 -37236 30935 -37210
rect 30615 -37864 30621 -37236
rect 30929 -37864 30935 -37236
rect 30615 -37890 30935 -37864
rect 31615 -37236 31935 -37210
rect 31615 -37864 31621 -37236
rect 31929 -37864 31935 -37236
rect 31615 -37890 31935 -37864
rect 32615 -37236 32935 -37210
rect 32615 -37864 32621 -37236
rect 32929 -37864 32935 -37236
rect 32615 -37890 32935 -37864
rect 33615 -37236 33935 -37210
rect 33615 -37864 33621 -37236
rect 33929 -37864 33935 -37236
rect 33615 -37890 33935 -37864
rect 8275 -37896 34275 -37890
rect 8275 -38204 8281 -37896
rect 8589 -37902 8961 -37896
rect 9589 -37902 9961 -37896
rect 10589 -37902 10961 -37896
rect 11589 -37902 11961 -37896
rect 12589 -37902 12961 -37896
rect 13589 -37902 13961 -37896
rect 14589 -37902 14961 -37896
rect 15589 -37902 15961 -37896
rect 16589 -37902 16961 -37896
rect 17589 -37902 17961 -37896
rect 18589 -37902 18961 -37896
rect 19589 -37902 19961 -37896
rect 20589 -37902 20961 -37896
rect 21589 -37902 21961 -37896
rect 22589 -37902 22961 -37896
rect 23589 -37902 23961 -37896
rect 24589 -37902 24961 -37896
rect 25589 -37902 25961 -37896
rect 26589 -37902 26961 -37896
rect 27589 -37902 27961 -37896
rect 28589 -37902 28961 -37896
rect 29589 -37902 29961 -37896
rect 30589 -37902 30961 -37896
rect 31589 -37902 31961 -37896
rect 32589 -37902 32961 -37896
rect 33589 -37902 33961 -37896
rect 8589 -38198 8627 -37902
rect 8923 -38198 8961 -37902
rect 9589 -38198 9627 -37902
rect 9923 -38198 9961 -37902
rect 10589 -38198 10627 -37902
rect 10923 -38198 10961 -37902
rect 11589 -38198 11627 -37902
rect 11923 -38198 11961 -37902
rect 12589 -38198 12627 -37902
rect 12923 -38198 12961 -37902
rect 13589 -38198 13627 -37902
rect 13923 -38198 13961 -37902
rect 14589 -38198 14627 -37902
rect 14923 -38198 14961 -37902
rect 15589 -38198 15627 -37902
rect 15923 -38198 15961 -37902
rect 16589 -38198 16627 -37902
rect 16923 -38198 16961 -37902
rect 17589 -38198 17627 -37902
rect 17923 -38198 17961 -37902
rect 18589 -38198 18627 -37902
rect 18923 -38198 18961 -37902
rect 19589 -38198 19627 -37902
rect 19923 -38198 19961 -37902
rect 20589 -38198 20627 -37902
rect 20923 -38198 20961 -37902
rect 21589 -38198 21627 -37902
rect 21923 -38198 21961 -37902
rect 22589 -38198 22627 -37902
rect 22923 -38198 22961 -37902
rect 23589 -38198 23627 -37902
rect 23923 -38198 23961 -37902
rect 24589 -38198 24627 -37902
rect 24923 -38198 24961 -37902
rect 25589 -38198 25627 -37902
rect 25923 -38198 25961 -37902
rect 26589 -38198 26627 -37902
rect 26923 -38198 26961 -37902
rect 27589 -38198 27627 -37902
rect 27923 -38198 27961 -37902
rect 28589 -38198 28627 -37902
rect 28923 -38198 28961 -37902
rect 29589 -38198 29627 -37902
rect 29923 -38198 29961 -37902
rect 30589 -38198 30627 -37902
rect 30923 -38198 30961 -37902
rect 31589 -38198 31627 -37902
rect 31923 -38198 31961 -37902
rect 32589 -38198 32627 -37902
rect 32923 -38198 32961 -37902
rect 33589 -38198 33627 -37902
rect 33923 -38198 33961 -37902
rect 8589 -38204 8961 -38198
rect 9589 -38204 9961 -38198
rect 10589 -38204 10961 -38198
rect 11589 -38204 11961 -38198
rect 12589 -38204 12961 -38198
rect 13589 -38204 13961 -38198
rect 14589 -38204 14961 -38198
rect 15589 -38204 15961 -38198
rect 16589 -38204 16961 -38198
rect 17589 -38204 17961 -38198
rect 18589 -38204 18961 -38198
rect 19589 -38204 19961 -38198
rect 20589 -38204 20961 -38198
rect 21589 -38204 21961 -38198
rect 22589 -38204 22961 -38198
rect 23589 -38204 23961 -38198
rect 24589 -38204 24961 -38198
rect 25589 -38204 25961 -38198
rect 26589 -38204 26961 -38198
rect 27589 -38204 27961 -38198
rect 28589 -38204 28961 -38198
rect 29589 -38204 29961 -38198
rect 30589 -38204 30961 -38198
rect 31589 -38204 31961 -38198
rect 32589 -38204 32961 -38198
rect 33589 -38204 33961 -38198
rect 34269 -38204 34275 -37896
rect 8275 -38210 34275 -38204
rect 8615 -38236 8935 -38210
rect 8615 -38864 8621 -38236
rect 8929 -38864 8935 -38236
rect 8615 -38890 8935 -38864
rect 9615 -38236 9935 -38210
rect 9615 -38864 9621 -38236
rect 9929 -38864 9935 -38236
rect 9615 -38890 9935 -38864
rect 10615 -38236 10935 -38210
rect 10615 -38864 10621 -38236
rect 10929 -38864 10935 -38236
rect 10615 -38890 10935 -38864
rect 11615 -38236 11935 -38210
rect 11615 -38864 11621 -38236
rect 11929 -38864 11935 -38236
rect 11615 -38890 11935 -38864
rect 12615 -38236 12935 -38210
rect 12615 -38864 12621 -38236
rect 12929 -38864 12935 -38236
rect 12615 -38890 12935 -38864
rect 13615 -38236 13935 -38210
rect 13615 -38864 13621 -38236
rect 13929 -38864 13935 -38236
rect 13615 -38890 13935 -38864
rect 14615 -38236 14935 -38210
rect 14615 -38864 14621 -38236
rect 14929 -38864 14935 -38236
rect 14615 -38890 14935 -38864
rect 15615 -38236 15935 -38210
rect 15615 -38864 15621 -38236
rect 15929 -38864 15935 -38236
rect 15615 -38890 15935 -38864
rect 16615 -38236 16935 -38210
rect 16615 -38864 16621 -38236
rect 16929 -38864 16935 -38236
rect 16615 -38890 16935 -38864
rect 17615 -38236 17935 -38210
rect 17615 -38864 17621 -38236
rect 17929 -38864 17935 -38236
rect 17615 -38890 17935 -38864
rect 18615 -38236 18935 -38210
rect 18615 -38864 18621 -38236
rect 18929 -38864 18935 -38236
rect 18615 -38890 18935 -38864
rect 19615 -38236 19935 -38210
rect 19615 -38864 19621 -38236
rect 19929 -38864 19935 -38236
rect 19615 -38890 19935 -38864
rect 20615 -38236 20935 -38210
rect 20615 -38864 20621 -38236
rect 20929 -38864 20935 -38236
rect 20615 -38890 20935 -38864
rect 21615 -38236 21935 -38210
rect 21615 -38864 21621 -38236
rect 21929 -38864 21935 -38236
rect 21615 -38890 21935 -38864
rect 22615 -38236 22935 -38210
rect 22615 -38864 22621 -38236
rect 22929 -38864 22935 -38236
rect 22615 -38890 22935 -38864
rect 23615 -38236 23935 -38210
rect 23615 -38864 23621 -38236
rect 23929 -38864 23935 -38236
rect 23615 -38890 23935 -38864
rect 24615 -38236 24935 -38210
rect 24615 -38864 24621 -38236
rect 24929 -38864 24935 -38236
rect 24615 -38890 24935 -38864
rect 25615 -38236 25935 -38210
rect 25615 -38864 25621 -38236
rect 25929 -38864 25935 -38236
rect 25615 -38890 25935 -38864
rect 26615 -38236 26935 -38210
rect 26615 -38864 26621 -38236
rect 26929 -38864 26935 -38236
rect 26615 -38890 26935 -38864
rect 27615 -38236 27935 -38210
rect 27615 -38864 27621 -38236
rect 27929 -38864 27935 -38236
rect 27615 -38890 27935 -38864
rect 28615 -38236 28935 -38210
rect 28615 -38864 28621 -38236
rect 28929 -38864 28935 -38236
rect 28615 -38890 28935 -38864
rect 29615 -38236 29935 -38210
rect 29615 -38864 29621 -38236
rect 29929 -38864 29935 -38236
rect 29615 -38890 29935 -38864
rect 30615 -38236 30935 -38210
rect 30615 -38864 30621 -38236
rect 30929 -38864 30935 -38236
rect 30615 -38890 30935 -38864
rect 31615 -38236 31935 -38210
rect 31615 -38864 31621 -38236
rect 31929 -38864 31935 -38236
rect 31615 -38890 31935 -38864
rect 32615 -38236 32935 -38210
rect 32615 -38864 32621 -38236
rect 32929 -38864 32935 -38236
rect 32615 -38890 32935 -38864
rect 33615 -38236 33935 -38210
rect 33615 -38864 33621 -38236
rect 33929 -38864 33935 -38236
rect 33615 -38890 33935 -38864
rect 8275 -38896 34275 -38890
rect 8275 -39204 8281 -38896
rect 8589 -38902 8961 -38896
rect 9589 -38902 9961 -38896
rect 10589 -38902 10961 -38896
rect 11589 -38902 11961 -38896
rect 12589 -38902 12961 -38896
rect 13589 -38902 13961 -38896
rect 14589 -38902 14961 -38896
rect 15589 -38902 15961 -38896
rect 16589 -38902 16961 -38896
rect 17589 -38902 17961 -38896
rect 18589 -38902 18961 -38896
rect 19589 -38902 19961 -38896
rect 20589 -38902 20961 -38896
rect 21589 -38902 21961 -38896
rect 22589 -38902 22961 -38896
rect 23589 -38902 23961 -38896
rect 24589 -38902 24961 -38896
rect 25589 -38902 25961 -38896
rect 26589 -38902 26961 -38896
rect 27589 -38902 27961 -38896
rect 28589 -38902 28961 -38896
rect 29589 -38902 29961 -38896
rect 30589 -38902 30961 -38896
rect 31589 -38902 31961 -38896
rect 32589 -38902 32961 -38896
rect 33589 -38902 33961 -38896
rect 8589 -39198 8627 -38902
rect 8923 -39198 8961 -38902
rect 9589 -39198 9627 -38902
rect 9923 -39198 9961 -38902
rect 10589 -39198 10627 -38902
rect 10923 -39198 10961 -38902
rect 11589 -39198 11627 -38902
rect 11923 -39198 11961 -38902
rect 12589 -39198 12627 -38902
rect 12923 -39198 12961 -38902
rect 13589 -39198 13627 -38902
rect 13923 -39198 13961 -38902
rect 14589 -39198 14627 -38902
rect 14923 -39198 14961 -38902
rect 15589 -39198 15627 -38902
rect 15923 -39198 15961 -38902
rect 16589 -39198 16627 -38902
rect 16923 -39198 16961 -38902
rect 17589 -39198 17627 -38902
rect 17923 -39198 17961 -38902
rect 18589 -39198 18627 -38902
rect 18923 -39198 18961 -38902
rect 19589 -39198 19627 -38902
rect 19923 -39198 19961 -38902
rect 20589 -39198 20627 -38902
rect 20923 -39198 20961 -38902
rect 21589 -39198 21627 -38902
rect 21923 -39198 21961 -38902
rect 22589 -39198 22627 -38902
rect 22923 -39198 22961 -38902
rect 23589 -39198 23627 -38902
rect 23923 -39198 23961 -38902
rect 24589 -39198 24627 -38902
rect 24923 -39198 24961 -38902
rect 25589 -39198 25627 -38902
rect 25923 -39198 25961 -38902
rect 26589 -39198 26627 -38902
rect 26923 -39198 26961 -38902
rect 27589 -39198 27627 -38902
rect 27923 -39198 27961 -38902
rect 28589 -39198 28627 -38902
rect 28923 -39198 28961 -38902
rect 29589 -39198 29627 -38902
rect 29923 -39198 29961 -38902
rect 30589 -39198 30627 -38902
rect 30923 -39198 30961 -38902
rect 31589 -39198 31627 -38902
rect 31923 -39198 31961 -38902
rect 32589 -39198 32627 -38902
rect 32923 -39198 32961 -38902
rect 33589 -39198 33627 -38902
rect 33923 -39198 33961 -38902
rect 8589 -39204 8961 -39198
rect 9589 -39204 9961 -39198
rect 10589 -39204 10961 -39198
rect 11589 -39204 11961 -39198
rect 12589 -39204 12961 -39198
rect 13589 -39204 13961 -39198
rect 14589 -39204 14961 -39198
rect 15589 -39204 15961 -39198
rect 16589 -39204 16961 -39198
rect 17589 -39204 17961 -39198
rect 18589 -39204 18961 -39198
rect 19589 -39204 19961 -39198
rect 20589 -39204 20961 -39198
rect 21589 -39204 21961 -39198
rect 22589 -39204 22961 -39198
rect 23589 -39204 23961 -39198
rect 24589 -39204 24961 -39198
rect 25589 -39204 25961 -39198
rect 26589 -39204 26961 -39198
rect 27589 -39204 27961 -39198
rect 28589 -39204 28961 -39198
rect 29589 -39204 29961 -39198
rect 30589 -39204 30961 -39198
rect 31589 -39204 31961 -39198
rect 32589 -39204 32961 -39198
rect 33589 -39204 33961 -39198
rect 34269 -39204 34275 -38896
rect 8275 -39210 34275 -39204
rect 8615 -39236 8935 -39210
rect 8615 -39864 8621 -39236
rect 8929 -39864 8935 -39236
rect 8615 -39890 8935 -39864
rect 9615 -39236 9935 -39210
rect 9615 -39864 9621 -39236
rect 9929 -39864 9935 -39236
rect 9615 -39890 9935 -39864
rect 10615 -39236 10935 -39210
rect 10615 -39864 10621 -39236
rect 10929 -39864 10935 -39236
rect 10615 -39890 10935 -39864
rect 11615 -39236 11935 -39210
rect 11615 -39864 11621 -39236
rect 11929 -39864 11935 -39236
rect 11615 -39890 11935 -39864
rect 12615 -39236 12935 -39210
rect 12615 -39864 12621 -39236
rect 12929 -39864 12935 -39236
rect 12615 -39890 12935 -39864
rect 13615 -39236 13935 -39210
rect 13615 -39864 13621 -39236
rect 13929 -39864 13935 -39236
rect 13615 -39890 13935 -39864
rect 14615 -39236 14935 -39210
rect 14615 -39864 14621 -39236
rect 14929 -39864 14935 -39236
rect 14615 -39890 14935 -39864
rect 15615 -39236 15935 -39210
rect 15615 -39864 15621 -39236
rect 15929 -39864 15935 -39236
rect 15615 -39890 15935 -39864
rect 16615 -39236 16935 -39210
rect 16615 -39864 16621 -39236
rect 16929 -39864 16935 -39236
rect 16615 -39890 16935 -39864
rect 17615 -39236 17935 -39210
rect 17615 -39864 17621 -39236
rect 17929 -39864 17935 -39236
rect 17615 -39890 17935 -39864
rect 18615 -39236 18935 -39210
rect 18615 -39864 18621 -39236
rect 18929 -39864 18935 -39236
rect 18615 -39890 18935 -39864
rect 19615 -39236 19935 -39210
rect 19615 -39864 19621 -39236
rect 19929 -39864 19935 -39236
rect 19615 -39890 19935 -39864
rect 20615 -39236 20935 -39210
rect 20615 -39864 20621 -39236
rect 20929 -39864 20935 -39236
rect 20615 -39890 20935 -39864
rect 21615 -39236 21935 -39210
rect 21615 -39864 21621 -39236
rect 21929 -39864 21935 -39236
rect 21615 -39890 21935 -39864
rect 22615 -39236 22935 -39210
rect 22615 -39864 22621 -39236
rect 22929 -39864 22935 -39236
rect 22615 -39890 22935 -39864
rect 23615 -39236 23935 -39210
rect 23615 -39864 23621 -39236
rect 23929 -39864 23935 -39236
rect 23615 -39890 23935 -39864
rect 24615 -39236 24935 -39210
rect 24615 -39864 24621 -39236
rect 24929 -39864 24935 -39236
rect 24615 -39890 24935 -39864
rect 25615 -39236 25935 -39210
rect 25615 -39864 25621 -39236
rect 25929 -39864 25935 -39236
rect 25615 -39890 25935 -39864
rect 26615 -39236 26935 -39210
rect 26615 -39864 26621 -39236
rect 26929 -39864 26935 -39236
rect 26615 -39890 26935 -39864
rect 27615 -39236 27935 -39210
rect 27615 -39864 27621 -39236
rect 27929 -39864 27935 -39236
rect 27615 -39890 27935 -39864
rect 28615 -39236 28935 -39210
rect 28615 -39864 28621 -39236
rect 28929 -39864 28935 -39236
rect 28615 -39890 28935 -39864
rect 29615 -39236 29935 -39210
rect 29615 -39864 29621 -39236
rect 29929 -39864 29935 -39236
rect 29615 -39890 29935 -39864
rect 30615 -39236 30935 -39210
rect 30615 -39864 30621 -39236
rect 30929 -39864 30935 -39236
rect 30615 -39890 30935 -39864
rect 31615 -39236 31935 -39210
rect 31615 -39864 31621 -39236
rect 31929 -39864 31935 -39236
rect 31615 -39890 31935 -39864
rect 32615 -39236 32935 -39210
rect 32615 -39864 32621 -39236
rect 32929 -39864 32935 -39236
rect 32615 -39890 32935 -39864
rect 33615 -39236 33935 -39210
rect 33615 -39864 33621 -39236
rect 33929 -39864 33935 -39236
rect 33615 -39890 33935 -39864
rect 8275 -39896 34275 -39890
rect 8275 -40204 8281 -39896
rect 8589 -39902 8961 -39896
rect 9589 -39902 9961 -39896
rect 10589 -39902 10961 -39896
rect 11589 -39902 11961 -39896
rect 12589 -39902 12961 -39896
rect 13589 -39902 13961 -39896
rect 14589 -39902 14961 -39896
rect 15589 -39902 15961 -39896
rect 16589 -39902 16961 -39896
rect 17589 -39902 17961 -39896
rect 18589 -39902 18961 -39896
rect 19589 -39902 19961 -39896
rect 20589 -39902 20961 -39896
rect 21589 -39902 21961 -39896
rect 22589 -39902 22961 -39896
rect 23589 -39902 23961 -39896
rect 24589 -39902 24961 -39896
rect 25589 -39902 25961 -39896
rect 26589 -39902 26961 -39896
rect 27589 -39902 27961 -39896
rect 28589 -39902 28961 -39896
rect 29589 -39902 29961 -39896
rect 30589 -39902 30961 -39896
rect 31589 -39902 31961 -39896
rect 32589 -39902 32961 -39896
rect 33589 -39902 33961 -39896
rect 8589 -40198 8627 -39902
rect 8923 -40198 8961 -39902
rect 9589 -40198 9627 -39902
rect 9923 -40198 9961 -39902
rect 10589 -40198 10627 -39902
rect 10923 -40198 10961 -39902
rect 11589 -40198 11627 -39902
rect 11923 -40198 11961 -39902
rect 12589 -40198 12627 -39902
rect 12923 -40198 12961 -39902
rect 13589 -40198 13627 -39902
rect 13923 -40198 13961 -39902
rect 14589 -40198 14627 -39902
rect 14923 -40198 14961 -39902
rect 15589 -40198 15627 -39902
rect 15923 -40198 15961 -39902
rect 16589 -40198 16627 -39902
rect 16923 -40198 16961 -39902
rect 17589 -40198 17627 -39902
rect 17923 -40198 17961 -39902
rect 18589 -40198 18627 -39902
rect 18923 -40198 18961 -39902
rect 19589 -40198 19627 -39902
rect 19923 -40198 19961 -39902
rect 20589 -40198 20627 -39902
rect 20923 -40198 20961 -39902
rect 21589 -40198 21627 -39902
rect 21923 -40198 21961 -39902
rect 22589 -40198 22627 -39902
rect 22923 -40198 22961 -39902
rect 23589 -40198 23627 -39902
rect 23923 -40198 23961 -39902
rect 24589 -40198 24627 -39902
rect 24923 -40198 24961 -39902
rect 25589 -40198 25627 -39902
rect 25923 -40198 25961 -39902
rect 26589 -40198 26627 -39902
rect 26923 -40198 26961 -39902
rect 27589 -40198 27627 -39902
rect 27923 -40198 27961 -39902
rect 28589 -40198 28627 -39902
rect 28923 -40198 28961 -39902
rect 29589 -40198 29627 -39902
rect 29923 -40198 29961 -39902
rect 30589 -40198 30627 -39902
rect 30923 -40198 30961 -39902
rect 31589 -40198 31627 -39902
rect 31923 -40198 31961 -39902
rect 32589 -40198 32627 -39902
rect 32923 -40198 32961 -39902
rect 33589 -40198 33627 -39902
rect 33923 -40198 33961 -39902
rect 8589 -40204 8961 -40198
rect 9589 -40204 9961 -40198
rect 10589 -40204 10961 -40198
rect 11589 -40204 11961 -40198
rect 12589 -40204 12961 -40198
rect 13589 -40204 13961 -40198
rect 14589 -40204 14961 -40198
rect 15589 -40204 15961 -40198
rect 16589 -40204 16961 -40198
rect 17589 -40204 17961 -40198
rect 18589 -40204 18961 -40198
rect 19589 -40204 19961 -40198
rect 20589 -40204 20961 -40198
rect 21589 -40204 21961 -40198
rect 22589 -40204 22961 -40198
rect 23589 -40204 23961 -40198
rect 24589 -40204 24961 -40198
rect 25589 -40204 25961 -40198
rect 26589 -40204 26961 -40198
rect 27589 -40204 27961 -40198
rect 28589 -40204 28961 -40198
rect 29589 -40204 29961 -40198
rect 30589 -40204 30961 -40198
rect 31589 -40204 31961 -40198
rect 32589 -40204 32961 -40198
rect 33589 -40204 33961 -40198
rect 34269 -40204 34275 -39896
rect 8275 -40210 34275 -40204
rect 8615 -40236 8935 -40210
rect 8615 -40864 8621 -40236
rect 8929 -40864 8935 -40236
rect 8615 -40890 8935 -40864
rect 9615 -40236 9935 -40210
rect 9615 -40864 9621 -40236
rect 9929 -40864 9935 -40236
rect 9615 -40890 9935 -40864
rect 10615 -40236 10935 -40210
rect 10615 -40864 10621 -40236
rect 10929 -40864 10935 -40236
rect 10615 -40890 10935 -40864
rect 11615 -40236 11935 -40210
rect 11615 -40864 11621 -40236
rect 11929 -40864 11935 -40236
rect 11615 -40890 11935 -40864
rect 12615 -40236 12935 -40210
rect 12615 -40864 12621 -40236
rect 12929 -40864 12935 -40236
rect 12615 -40890 12935 -40864
rect 13615 -40236 13935 -40210
rect 13615 -40864 13621 -40236
rect 13929 -40864 13935 -40236
rect 13615 -40890 13935 -40864
rect 14615 -40236 14935 -40210
rect 14615 -40864 14621 -40236
rect 14929 -40864 14935 -40236
rect 14615 -40890 14935 -40864
rect 15615 -40236 15935 -40210
rect 15615 -40864 15621 -40236
rect 15929 -40864 15935 -40236
rect 15615 -40890 15935 -40864
rect 16615 -40236 16935 -40210
rect 16615 -40864 16621 -40236
rect 16929 -40864 16935 -40236
rect 16615 -40890 16935 -40864
rect 17615 -40236 17935 -40210
rect 17615 -40864 17621 -40236
rect 17929 -40864 17935 -40236
rect 17615 -40890 17935 -40864
rect 18615 -40236 18935 -40210
rect 18615 -40864 18621 -40236
rect 18929 -40864 18935 -40236
rect 18615 -40890 18935 -40864
rect 19615 -40236 19935 -40210
rect 19615 -40864 19621 -40236
rect 19929 -40864 19935 -40236
rect 19615 -40890 19935 -40864
rect 20615 -40236 20935 -40210
rect 20615 -40864 20621 -40236
rect 20929 -40864 20935 -40236
rect 20615 -40890 20935 -40864
rect 21615 -40236 21935 -40210
rect 21615 -40864 21621 -40236
rect 21929 -40864 21935 -40236
rect 21615 -40890 21935 -40864
rect 22615 -40236 22935 -40210
rect 22615 -40864 22621 -40236
rect 22929 -40864 22935 -40236
rect 22615 -40890 22935 -40864
rect 23615 -40236 23935 -40210
rect 23615 -40864 23621 -40236
rect 23929 -40864 23935 -40236
rect 23615 -40890 23935 -40864
rect 24615 -40236 24935 -40210
rect 24615 -40864 24621 -40236
rect 24929 -40864 24935 -40236
rect 24615 -40890 24935 -40864
rect 25615 -40236 25935 -40210
rect 25615 -40864 25621 -40236
rect 25929 -40864 25935 -40236
rect 25615 -40890 25935 -40864
rect 26615 -40236 26935 -40210
rect 26615 -40864 26621 -40236
rect 26929 -40864 26935 -40236
rect 26615 -40890 26935 -40864
rect 27615 -40236 27935 -40210
rect 27615 -40864 27621 -40236
rect 27929 -40864 27935 -40236
rect 27615 -40890 27935 -40864
rect 28615 -40236 28935 -40210
rect 28615 -40864 28621 -40236
rect 28929 -40864 28935 -40236
rect 28615 -40890 28935 -40864
rect 29615 -40236 29935 -40210
rect 29615 -40864 29621 -40236
rect 29929 -40864 29935 -40236
rect 29615 -40890 29935 -40864
rect 30615 -40236 30935 -40210
rect 30615 -40864 30621 -40236
rect 30929 -40864 30935 -40236
rect 30615 -40890 30935 -40864
rect 31615 -40236 31935 -40210
rect 31615 -40864 31621 -40236
rect 31929 -40864 31935 -40236
rect 31615 -40890 31935 -40864
rect 32615 -40236 32935 -40210
rect 32615 -40864 32621 -40236
rect 32929 -40864 32935 -40236
rect 32615 -40890 32935 -40864
rect 33615 -40236 33935 -40210
rect 33615 -40864 33621 -40236
rect 33929 -40864 33935 -40236
rect 33615 -40890 33935 -40864
rect 8275 -40896 34275 -40890
rect 8275 -41204 8281 -40896
rect 8589 -40902 8961 -40896
rect 9589 -40902 9961 -40896
rect 10589 -40902 10961 -40896
rect 11589 -40902 11961 -40896
rect 12589 -40902 12961 -40896
rect 13589 -40902 13961 -40896
rect 14589 -40902 14961 -40896
rect 15589 -40902 15961 -40896
rect 16589 -40902 16961 -40896
rect 17589 -40902 17961 -40896
rect 18589 -40902 18961 -40896
rect 19589 -40902 19961 -40896
rect 20589 -40902 20961 -40896
rect 21589 -40902 21961 -40896
rect 22589 -40902 22961 -40896
rect 23589 -40902 23961 -40896
rect 24589 -40902 24961 -40896
rect 25589 -40902 25961 -40896
rect 26589 -40902 26961 -40896
rect 27589 -40902 27961 -40896
rect 28589 -40902 28961 -40896
rect 29589 -40902 29961 -40896
rect 30589 -40902 30961 -40896
rect 31589 -40902 31961 -40896
rect 32589 -40902 32961 -40896
rect 33589 -40902 33961 -40896
rect 8589 -41198 8627 -40902
rect 8923 -41198 8961 -40902
rect 9589 -41198 9627 -40902
rect 9923 -41198 9961 -40902
rect 10589 -41198 10627 -40902
rect 10923 -41198 10961 -40902
rect 11589 -41198 11627 -40902
rect 11923 -41198 11961 -40902
rect 12589 -41198 12627 -40902
rect 12923 -41198 12961 -40902
rect 13589 -41198 13627 -40902
rect 13923 -41198 13961 -40902
rect 14589 -41198 14627 -40902
rect 14923 -41198 14961 -40902
rect 15589 -41198 15627 -40902
rect 15923 -41198 15961 -40902
rect 16589 -41198 16627 -40902
rect 16923 -41198 16961 -40902
rect 17589 -41198 17627 -40902
rect 17923 -41198 17961 -40902
rect 18589 -41198 18627 -40902
rect 18923 -41198 18961 -40902
rect 19589 -41198 19627 -40902
rect 19923 -41198 19961 -40902
rect 20589 -41198 20627 -40902
rect 20923 -41198 20961 -40902
rect 21589 -41198 21627 -40902
rect 21923 -41198 21961 -40902
rect 22589 -41198 22627 -40902
rect 22923 -41198 22961 -40902
rect 23589 -41198 23627 -40902
rect 23923 -41198 23961 -40902
rect 24589 -41198 24627 -40902
rect 24923 -41198 24961 -40902
rect 25589 -41198 25627 -40902
rect 25923 -41198 25961 -40902
rect 26589 -41198 26627 -40902
rect 26923 -41198 26961 -40902
rect 27589 -41198 27627 -40902
rect 27923 -41198 27961 -40902
rect 28589 -41198 28627 -40902
rect 28923 -41198 28961 -40902
rect 29589 -41198 29627 -40902
rect 29923 -41198 29961 -40902
rect 30589 -41198 30627 -40902
rect 30923 -41198 30961 -40902
rect 31589 -41198 31627 -40902
rect 31923 -41198 31961 -40902
rect 32589 -41198 32627 -40902
rect 32923 -41198 32961 -40902
rect 33589 -41198 33627 -40902
rect 33923 -41198 33961 -40902
rect 8589 -41204 8961 -41198
rect 9589 -41204 9961 -41198
rect 10589 -41204 10961 -41198
rect 11589 -41204 11961 -41198
rect 12589 -41204 12961 -41198
rect 13589 -41204 13961 -41198
rect 14589 -41204 14961 -41198
rect 15589 -41204 15961 -41198
rect 16589 -41204 16961 -41198
rect 17589 -41204 17961 -41198
rect 18589 -41204 18961 -41198
rect 19589 -41204 19961 -41198
rect 20589 -41204 20961 -41198
rect 21589 -41204 21961 -41198
rect 22589 -41204 22961 -41198
rect 23589 -41204 23961 -41198
rect 24589 -41204 24961 -41198
rect 25589 -41204 25961 -41198
rect 26589 -41204 26961 -41198
rect 27589 -41204 27961 -41198
rect 28589 -41204 28961 -41198
rect 29589 -41204 29961 -41198
rect 30589 -41204 30961 -41198
rect 31589 -41204 31961 -41198
rect 32589 -41204 32961 -41198
rect 33589 -41204 33961 -41198
rect 34269 -41204 34275 -40896
rect 8275 -41210 34275 -41204
rect 8615 -41236 8935 -41210
rect 8615 -41864 8621 -41236
rect 8929 -41864 8935 -41236
rect 8615 -41890 8935 -41864
rect 9615 -41236 9935 -41210
rect 9615 -41864 9621 -41236
rect 9929 -41864 9935 -41236
rect 9615 -41890 9935 -41864
rect 10615 -41236 10935 -41210
rect 10615 -41864 10621 -41236
rect 10929 -41864 10935 -41236
rect 10615 -41890 10935 -41864
rect 11615 -41236 11935 -41210
rect 11615 -41864 11621 -41236
rect 11929 -41864 11935 -41236
rect 11615 -41890 11935 -41864
rect 12615 -41236 12935 -41210
rect 12615 -41864 12621 -41236
rect 12929 -41864 12935 -41236
rect 12615 -41890 12935 -41864
rect 13615 -41236 13935 -41210
rect 13615 -41864 13621 -41236
rect 13929 -41864 13935 -41236
rect 13615 -41890 13935 -41864
rect 14615 -41236 14935 -41210
rect 14615 -41864 14621 -41236
rect 14929 -41864 14935 -41236
rect 14615 -41890 14935 -41864
rect 15615 -41236 15935 -41210
rect 15615 -41864 15621 -41236
rect 15929 -41864 15935 -41236
rect 15615 -41890 15935 -41864
rect 16615 -41236 16935 -41210
rect 16615 -41864 16621 -41236
rect 16929 -41864 16935 -41236
rect 16615 -41890 16935 -41864
rect 17615 -41236 17935 -41210
rect 17615 -41864 17621 -41236
rect 17929 -41864 17935 -41236
rect 17615 -41890 17935 -41864
rect 18615 -41236 18935 -41210
rect 18615 -41864 18621 -41236
rect 18929 -41864 18935 -41236
rect 18615 -41890 18935 -41864
rect 19615 -41236 19935 -41210
rect 19615 -41864 19621 -41236
rect 19929 -41864 19935 -41236
rect 19615 -41890 19935 -41864
rect 20615 -41236 20935 -41210
rect 20615 -41864 20621 -41236
rect 20929 -41864 20935 -41236
rect 20615 -41890 20935 -41864
rect 21615 -41236 21935 -41210
rect 21615 -41864 21621 -41236
rect 21929 -41864 21935 -41236
rect 21615 -41890 21935 -41864
rect 22615 -41236 22935 -41210
rect 22615 -41864 22621 -41236
rect 22929 -41864 22935 -41236
rect 22615 -41890 22935 -41864
rect 23615 -41236 23935 -41210
rect 23615 -41864 23621 -41236
rect 23929 -41864 23935 -41236
rect 23615 -41890 23935 -41864
rect 24615 -41236 24935 -41210
rect 24615 -41864 24621 -41236
rect 24929 -41864 24935 -41236
rect 24615 -41890 24935 -41864
rect 25615 -41236 25935 -41210
rect 25615 -41864 25621 -41236
rect 25929 -41864 25935 -41236
rect 25615 -41890 25935 -41864
rect 26615 -41236 26935 -41210
rect 26615 -41864 26621 -41236
rect 26929 -41864 26935 -41236
rect 26615 -41890 26935 -41864
rect 27615 -41236 27935 -41210
rect 27615 -41864 27621 -41236
rect 27929 -41864 27935 -41236
rect 27615 -41890 27935 -41864
rect 28615 -41236 28935 -41210
rect 28615 -41864 28621 -41236
rect 28929 -41864 28935 -41236
rect 28615 -41890 28935 -41864
rect 29615 -41236 29935 -41210
rect 29615 -41864 29621 -41236
rect 29929 -41864 29935 -41236
rect 29615 -41890 29935 -41864
rect 30615 -41236 30935 -41210
rect 30615 -41864 30621 -41236
rect 30929 -41864 30935 -41236
rect 30615 -41890 30935 -41864
rect 31615 -41236 31935 -41210
rect 31615 -41864 31621 -41236
rect 31929 -41864 31935 -41236
rect 31615 -41890 31935 -41864
rect 32615 -41236 32935 -41210
rect 32615 -41864 32621 -41236
rect 32929 -41864 32935 -41236
rect 32615 -41890 32935 -41864
rect 33615 -41236 33935 -41210
rect 33615 -41864 33621 -41236
rect 33929 -41864 33935 -41236
rect 33615 -41890 33935 -41864
rect 8275 -41896 34275 -41890
rect 8275 -42204 8281 -41896
rect 8589 -41902 8961 -41896
rect 9589 -41902 9961 -41896
rect 10589 -41902 10961 -41896
rect 11589 -41902 11961 -41896
rect 12589 -41902 12961 -41896
rect 13589 -41902 13961 -41896
rect 14589 -41902 14961 -41896
rect 15589 -41902 15961 -41896
rect 16589 -41902 16961 -41896
rect 17589 -41902 17961 -41896
rect 18589 -41902 18961 -41896
rect 19589 -41902 19961 -41896
rect 20589 -41902 20961 -41896
rect 21589 -41902 21961 -41896
rect 22589 -41902 22961 -41896
rect 23589 -41902 23961 -41896
rect 24589 -41902 24961 -41896
rect 25589 -41902 25961 -41896
rect 26589 -41902 26961 -41896
rect 27589 -41902 27961 -41896
rect 28589 -41902 28961 -41896
rect 29589 -41902 29961 -41896
rect 30589 -41902 30961 -41896
rect 31589 -41902 31961 -41896
rect 32589 -41902 32961 -41896
rect 33589 -41902 33961 -41896
rect 8589 -42198 8627 -41902
rect 8923 -42198 8961 -41902
rect 9589 -42198 9627 -41902
rect 9923 -42198 9961 -41902
rect 10589 -42198 10627 -41902
rect 10923 -42198 10961 -41902
rect 11589 -42198 11627 -41902
rect 11923 -42198 11961 -41902
rect 12589 -42198 12627 -41902
rect 12923 -42198 12961 -41902
rect 13589 -42198 13627 -41902
rect 13923 -42198 13961 -41902
rect 14589 -42198 14627 -41902
rect 14923 -42198 14961 -41902
rect 15589 -42198 15627 -41902
rect 15923 -42198 15961 -41902
rect 16589 -42198 16627 -41902
rect 16923 -42198 16961 -41902
rect 17589 -42198 17627 -41902
rect 17923 -42198 17961 -41902
rect 18589 -42198 18627 -41902
rect 18923 -42198 18961 -41902
rect 19589 -42198 19627 -41902
rect 19923 -42198 19961 -41902
rect 20589 -42198 20627 -41902
rect 20923 -42198 20961 -41902
rect 21589 -42198 21627 -41902
rect 21923 -42198 21961 -41902
rect 22589 -42198 22627 -41902
rect 22923 -42198 22961 -41902
rect 23589 -42198 23627 -41902
rect 23923 -42198 23961 -41902
rect 24589 -42198 24627 -41902
rect 24923 -42198 24961 -41902
rect 25589 -42198 25627 -41902
rect 25923 -42198 25961 -41902
rect 26589 -42198 26627 -41902
rect 26923 -42198 26961 -41902
rect 27589 -42198 27627 -41902
rect 27923 -42198 27961 -41902
rect 28589 -42198 28627 -41902
rect 28923 -42198 28961 -41902
rect 29589 -42198 29627 -41902
rect 29923 -42198 29961 -41902
rect 30589 -42198 30627 -41902
rect 30923 -42198 30961 -41902
rect 31589 -42198 31627 -41902
rect 31923 -42198 31961 -41902
rect 32589 -42198 32627 -41902
rect 32923 -42198 32961 -41902
rect 33589 -42198 33627 -41902
rect 33923 -42198 33961 -41902
rect 8589 -42204 8961 -42198
rect 9589 -42204 9961 -42198
rect 10589 -42204 10961 -42198
rect 11589 -42204 11961 -42198
rect 12589 -42204 12961 -42198
rect 13589 -42204 13961 -42198
rect 14589 -42204 14961 -42198
rect 15589 -42204 15961 -42198
rect 16589 -42204 16961 -42198
rect 17589 -42204 17961 -42198
rect 18589 -42204 18961 -42198
rect 19589 -42204 19961 -42198
rect 20589 -42204 20961 -42198
rect 21589 -42204 21961 -42198
rect 22589 -42204 22961 -42198
rect 23589 -42204 23961 -42198
rect 24589 -42204 24961 -42198
rect 25589 -42204 25961 -42198
rect 26589 -42204 26961 -42198
rect 27589 -42204 27961 -42198
rect 28589 -42204 28961 -42198
rect 29589 -42204 29961 -42198
rect 30589 -42204 30961 -42198
rect 31589 -42204 31961 -42198
rect 32589 -42204 32961 -42198
rect 33589 -42204 33961 -42198
rect 34269 -42204 34275 -41896
rect 8275 -42210 34275 -42204
rect 8615 -42236 8935 -42210
rect 8615 -42864 8621 -42236
rect 8929 -42864 8935 -42236
rect 8615 -42890 8935 -42864
rect 9615 -42236 9935 -42210
rect 9615 -42864 9621 -42236
rect 9929 -42864 9935 -42236
rect 9615 -42890 9935 -42864
rect 10615 -42236 10935 -42210
rect 10615 -42864 10621 -42236
rect 10929 -42864 10935 -42236
rect 10615 -42890 10935 -42864
rect 11615 -42236 11935 -42210
rect 11615 -42864 11621 -42236
rect 11929 -42864 11935 -42236
rect 11615 -42890 11935 -42864
rect 12615 -42236 12935 -42210
rect 12615 -42864 12621 -42236
rect 12929 -42864 12935 -42236
rect 12615 -42890 12935 -42864
rect 13615 -42236 13935 -42210
rect 13615 -42864 13621 -42236
rect 13929 -42864 13935 -42236
rect 13615 -42890 13935 -42864
rect 14615 -42236 14935 -42210
rect 14615 -42864 14621 -42236
rect 14929 -42864 14935 -42236
rect 14615 -42890 14935 -42864
rect 15615 -42236 15935 -42210
rect 15615 -42864 15621 -42236
rect 15929 -42864 15935 -42236
rect 15615 -42890 15935 -42864
rect 16615 -42236 16935 -42210
rect 16615 -42864 16621 -42236
rect 16929 -42864 16935 -42236
rect 16615 -42890 16935 -42864
rect 17615 -42236 17935 -42210
rect 17615 -42864 17621 -42236
rect 17929 -42864 17935 -42236
rect 17615 -42890 17935 -42864
rect 18615 -42236 18935 -42210
rect 18615 -42864 18621 -42236
rect 18929 -42864 18935 -42236
rect 18615 -42890 18935 -42864
rect 19615 -42236 19935 -42210
rect 19615 -42864 19621 -42236
rect 19929 -42864 19935 -42236
rect 19615 -42890 19935 -42864
rect 20615 -42236 20935 -42210
rect 20615 -42864 20621 -42236
rect 20929 -42864 20935 -42236
rect 20615 -42890 20935 -42864
rect 21615 -42236 21935 -42210
rect 21615 -42864 21621 -42236
rect 21929 -42864 21935 -42236
rect 21615 -42890 21935 -42864
rect 22615 -42236 22935 -42210
rect 22615 -42864 22621 -42236
rect 22929 -42864 22935 -42236
rect 22615 -42890 22935 -42864
rect 23615 -42236 23935 -42210
rect 23615 -42864 23621 -42236
rect 23929 -42864 23935 -42236
rect 23615 -42890 23935 -42864
rect 24615 -42236 24935 -42210
rect 24615 -42864 24621 -42236
rect 24929 -42864 24935 -42236
rect 24615 -42890 24935 -42864
rect 25615 -42236 25935 -42210
rect 25615 -42864 25621 -42236
rect 25929 -42864 25935 -42236
rect 25615 -42890 25935 -42864
rect 26615 -42236 26935 -42210
rect 26615 -42864 26621 -42236
rect 26929 -42864 26935 -42236
rect 26615 -42890 26935 -42864
rect 27615 -42236 27935 -42210
rect 27615 -42864 27621 -42236
rect 27929 -42864 27935 -42236
rect 27615 -42890 27935 -42864
rect 28615 -42236 28935 -42210
rect 28615 -42864 28621 -42236
rect 28929 -42864 28935 -42236
rect 28615 -42890 28935 -42864
rect 29615 -42236 29935 -42210
rect 29615 -42864 29621 -42236
rect 29929 -42864 29935 -42236
rect 29615 -42890 29935 -42864
rect 30615 -42236 30935 -42210
rect 30615 -42864 30621 -42236
rect 30929 -42864 30935 -42236
rect 30615 -42890 30935 -42864
rect 31615 -42236 31935 -42210
rect 31615 -42864 31621 -42236
rect 31929 -42864 31935 -42236
rect 31615 -42890 31935 -42864
rect 32615 -42236 32935 -42210
rect 32615 -42864 32621 -42236
rect 32929 -42864 32935 -42236
rect 32615 -42890 32935 -42864
rect 33615 -42236 33935 -42210
rect 33615 -42864 33621 -42236
rect 33929 -42864 33935 -42236
rect 33615 -42890 33935 -42864
rect 8275 -42896 34275 -42890
rect 8275 -43204 8281 -42896
rect 8589 -42902 8961 -42896
rect 9589 -42902 9961 -42896
rect 10589 -42902 10961 -42896
rect 11589 -42902 11961 -42896
rect 12589 -42902 12961 -42896
rect 13589 -42902 13961 -42896
rect 14589 -42902 14961 -42896
rect 15589 -42902 15961 -42896
rect 16589 -42902 16961 -42896
rect 17589 -42902 17961 -42896
rect 18589 -42902 18961 -42896
rect 19589 -42902 19961 -42896
rect 20589 -42902 20961 -42896
rect 21589 -42902 21961 -42896
rect 22589 -42902 22961 -42896
rect 23589 -42902 23961 -42896
rect 24589 -42902 24961 -42896
rect 25589 -42902 25961 -42896
rect 26589 -42902 26961 -42896
rect 27589 -42902 27961 -42896
rect 28589 -42902 28961 -42896
rect 29589 -42902 29961 -42896
rect 30589 -42902 30961 -42896
rect 31589 -42902 31961 -42896
rect 32589 -42902 32961 -42896
rect 33589 -42902 33961 -42896
rect 8589 -43198 8627 -42902
rect 8923 -43198 8961 -42902
rect 9589 -43198 9627 -42902
rect 9923 -43198 9961 -42902
rect 10589 -43198 10627 -42902
rect 10923 -43198 10961 -42902
rect 11589 -43198 11627 -42902
rect 11923 -43198 11961 -42902
rect 12589 -43198 12627 -42902
rect 12923 -43198 12961 -42902
rect 13589 -43198 13627 -42902
rect 13923 -43198 13961 -42902
rect 14589 -43198 14627 -42902
rect 14923 -43198 14961 -42902
rect 15589 -43198 15627 -42902
rect 15923 -43198 15961 -42902
rect 16589 -43198 16627 -42902
rect 16923 -43198 16961 -42902
rect 17589 -43198 17627 -42902
rect 17923 -43198 17961 -42902
rect 18589 -43198 18627 -42902
rect 18923 -43198 18961 -42902
rect 19589 -43198 19627 -42902
rect 19923 -43198 19961 -42902
rect 20589 -43198 20627 -42902
rect 20923 -43198 20961 -42902
rect 21589 -43198 21627 -42902
rect 21923 -43198 21961 -42902
rect 22589 -43198 22627 -42902
rect 22923 -43198 22961 -42902
rect 23589 -43198 23627 -42902
rect 23923 -43198 23961 -42902
rect 24589 -43198 24627 -42902
rect 24923 -43198 24961 -42902
rect 25589 -43198 25627 -42902
rect 25923 -43198 25961 -42902
rect 26589 -43198 26627 -42902
rect 26923 -43198 26961 -42902
rect 27589 -43198 27627 -42902
rect 27923 -43198 27961 -42902
rect 28589 -43198 28627 -42902
rect 28923 -43198 28961 -42902
rect 29589 -43198 29627 -42902
rect 29923 -43198 29961 -42902
rect 30589 -43198 30627 -42902
rect 30923 -43198 30961 -42902
rect 31589 -43198 31627 -42902
rect 31923 -43198 31961 -42902
rect 32589 -43198 32627 -42902
rect 32923 -43198 32961 -42902
rect 33589 -43198 33627 -42902
rect 33923 -43198 33961 -42902
rect 8589 -43204 8961 -43198
rect 9589 -43204 9961 -43198
rect 10589 -43204 10961 -43198
rect 11589 -43204 11961 -43198
rect 12589 -43204 12961 -43198
rect 13589 -43204 13961 -43198
rect 14589 -43204 14961 -43198
rect 15589 -43204 15961 -43198
rect 16589 -43204 16961 -43198
rect 17589 -43204 17961 -43198
rect 18589 -43204 18961 -43198
rect 19589 -43204 19961 -43198
rect 20589 -43204 20961 -43198
rect 21589 -43204 21961 -43198
rect 22589 -43204 22961 -43198
rect 23589 -43204 23961 -43198
rect 24589 -43204 24961 -43198
rect 25589 -43204 25961 -43198
rect 26589 -43204 26961 -43198
rect 27589 -43204 27961 -43198
rect 28589 -43204 28961 -43198
rect 29589 -43204 29961 -43198
rect 30589 -43204 30961 -43198
rect 31589 -43204 31961 -43198
rect 32589 -43204 32961 -43198
rect 33589 -43204 33961 -43198
rect 34269 -43204 34275 -42896
rect 8275 -43210 34275 -43204
rect 8615 -43236 8935 -43210
rect 8615 -43864 8621 -43236
rect 8929 -43864 8935 -43236
rect 8615 -43890 8935 -43864
rect 9615 -43236 9935 -43210
rect 9615 -43864 9621 -43236
rect 9929 -43864 9935 -43236
rect 9615 -43890 9935 -43864
rect 10615 -43236 10935 -43210
rect 10615 -43864 10621 -43236
rect 10929 -43864 10935 -43236
rect 10615 -43890 10935 -43864
rect 11615 -43236 11935 -43210
rect 11615 -43864 11621 -43236
rect 11929 -43864 11935 -43236
rect 11615 -43890 11935 -43864
rect 12615 -43236 12935 -43210
rect 12615 -43864 12621 -43236
rect 12929 -43864 12935 -43236
rect 12615 -43890 12935 -43864
rect 13615 -43236 13935 -43210
rect 13615 -43864 13621 -43236
rect 13929 -43864 13935 -43236
rect 13615 -43890 13935 -43864
rect 14615 -43236 14935 -43210
rect 14615 -43864 14621 -43236
rect 14929 -43864 14935 -43236
rect 14615 -43890 14935 -43864
rect 15615 -43236 15935 -43210
rect 15615 -43864 15621 -43236
rect 15929 -43864 15935 -43236
rect 15615 -43890 15935 -43864
rect 16615 -43236 16935 -43210
rect 16615 -43864 16621 -43236
rect 16929 -43864 16935 -43236
rect 16615 -43890 16935 -43864
rect 17615 -43236 17935 -43210
rect 17615 -43864 17621 -43236
rect 17929 -43864 17935 -43236
rect 17615 -43890 17935 -43864
rect 18615 -43236 18935 -43210
rect 18615 -43864 18621 -43236
rect 18929 -43864 18935 -43236
rect 18615 -43890 18935 -43864
rect 19615 -43236 19935 -43210
rect 19615 -43864 19621 -43236
rect 19929 -43864 19935 -43236
rect 19615 -43890 19935 -43864
rect 20615 -43236 20935 -43210
rect 20615 -43864 20621 -43236
rect 20929 -43864 20935 -43236
rect 20615 -43890 20935 -43864
rect 21615 -43236 21935 -43210
rect 21615 -43864 21621 -43236
rect 21929 -43864 21935 -43236
rect 21615 -43890 21935 -43864
rect 22615 -43236 22935 -43210
rect 22615 -43864 22621 -43236
rect 22929 -43864 22935 -43236
rect 22615 -43890 22935 -43864
rect 23615 -43236 23935 -43210
rect 23615 -43864 23621 -43236
rect 23929 -43864 23935 -43236
rect 23615 -43890 23935 -43864
rect 24615 -43236 24935 -43210
rect 24615 -43864 24621 -43236
rect 24929 -43864 24935 -43236
rect 24615 -43890 24935 -43864
rect 25615 -43236 25935 -43210
rect 25615 -43864 25621 -43236
rect 25929 -43864 25935 -43236
rect 25615 -43890 25935 -43864
rect 26615 -43236 26935 -43210
rect 26615 -43864 26621 -43236
rect 26929 -43864 26935 -43236
rect 26615 -43890 26935 -43864
rect 27615 -43236 27935 -43210
rect 27615 -43864 27621 -43236
rect 27929 -43864 27935 -43236
rect 27615 -43890 27935 -43864
rect 28615 -43236 28935 -43210
rect 28615 -43864 28621 -43236
rect 28929 -43864 28935 -43236
rect 28615 -43890 28935 -43864
rect 29615 -43236 29935 -43210
rect 29615 -43864 29621 -43236
rect 29929 -43864 29935 -43236
rect 29615 -43890 29935 -43864
rect 30615 -43236 30935 -43210
rect 30615 -43864 30621 -43236
rect 30929 -43864 30935 -43236
rect 30615 -43890 30935 -43864
rect 31615 -43236 31935 -43210
rect 31615 -43864 31621 -43236
rect 31929 -43864 31935 -43236
rect 31615 -43890 31935 -43864
rect 32615 -43236 32935 -43210
rect 32615 -43864 32621 -43236
rect 32929 -43864 32935 -43236
rect 32615 -43890 32935 -43864
rect 33615 -43236 33935 -43210
rect 33615 -43864 33621 -43236
rect 33929 -43864 33935 -43236
rect 33615 -43890 33935 -43864
rect 8275 -43896 34275 -43890
rect 8275 -44204 8281 -43896
rect 8589 -43902 8961 -43896
rect 9589 -43902 9961 -43896
rect 10589 -43902 10961 -43896
rect 11589 -43902 11961 -43896
rect 12589 -43902 12961 -43896
rect 13589 -43902 13961 -43896
rect 14589 -43902 14961 -43896
rect 15589 -43902 15961 -43896
rect 16589 -43902 16961 -43896
rect 17589 -43902 17961 -43896
rect 18589 -43902 18961 -43896
rect 19589 -43902 19961 -43896
rect 20589 -43902 20961 -43896
rect 21589 -43902 21961 -43896
rect 22589 -43902 22961 -43896
rect 23589 -43902 23961 -43896
rect 24589 -43902 24961 -43896
rect 25589 -43902 25961 -43896
rect 26589 -43902 26961 -43896
rect 27589 -43902 27961 -43896
rect 28589 -43902 28961 -43896
rect 29589 -43902 29961 -43896
rect 30589 -43902 30961 -43896
rect 31589 -43902 31961 -43896
rect 32589 -43902 32961 -43896
rect 33589 -43902 33961 -43896
rect 8589 -44198 8627 -43902
rect 8923 -44198 8961 -43902
rect 9589 -44198 9627 -43902
rect 9923 -44198 9961 -43902
rect 10589 -44198 10627 -43902
rect 10923 -44198 10961 -43902
rect 11589 -44198 11627 -43902
rect 11923 -44198 11961 -43902
rect 12589 -44198 12627 -43902
rect 12923 -44198 12961 -43902
rect 13589 -44198 13627 -43902
rect 13923 -44198 13961 -43902
rect 14589 -44198 14627 -43902
rect 14923 -44198 14961 -43902
rect 15589 -44198 15627 -43902
rect 15923 -44198 15961 -43902
rect 16589 -44198 16627 -43902
rect 16923 -44198 16961 -43902
rect 17589 -44198 17627 -43902
rect 17923 -44198 17961 -43902
rect 18589 -44198 18627 -43902
rect 18923 -44198 18961 -43902
rect 19589 -44198 19627 -43902
rect 19923 -44198 19961 -43902
rect 20589 -44198 20627 -43902
rect 20923 -44198 20961 -43902
rect 21589 -44198 21627 -43902
rect 21923 -44198 21961 -43902
rect 22589 -44198 22627 -43902
rect 22923 -44198 22961 -43902
rect 23589 -44198 23627 -43902
rect 23923 -44198 23961 -43902
rect 24589 -44198 24627 -43902
rect 24923 -44198 24961 -43902
rect 25589 -44198 25627 -43902
rect 25923 -44198 25961 -43902
rect 26589 -44198 26627 -43902
rect 26923 -44198 26961 -43902
rect 27589 -44198 27627 -43902
rect 27923 -44198 27961 -43902
rect 28589 -44198 28627 -43902
rect 28923 -44198 28961 -43902
rect 29589 -44198 29627 -43902
rect 29923 -44198 29961 -43902
rect 30589 -44198 30627 -43902
rect 30923 -44198 30961 -43902
rect 31589 -44198 31627 -43902
rect 31923 -44198 31961 -43902
rect 32589 -44198 32627 -43902
rect 32923 -44198 32961 -43902
rect 33589 -44198 33627 -43902
rect 33923 -44198 33961 -43902
rect 8589 -44204 8961 -44198
rect 9589 -44204 9961 -44198
rect 10589 -44204 10961 -44198
rect 11589 -44204 11961 -44198
rect 12589 -44204 12961 -44198
rect 13589 -44204 13961 -44198
rect 14589 -44204 14961 -44198
rect 15589 -44204 15961 -44198
rect 16589 -44204 16961 -44198
rect 17589 -44204 17961 -44198
rect 18589 -44204 18961 -44198
rect 19589 -44204 19961 -44198
rect 20589 -44204 20961 -44198
rect 21589 -44204 21961 -44198
rect 22589 -44204 22961 -44198
rect 23589 -44204 23961 -44198
rect 24589 -44204 24961 -44198
rect 25589 -44204 25961 -44198
rect 26589 -44204 26961 -44198
rect 27589 -44204 27961 -44198
rect 28589 -44204 28961 -44198
rect 29589 -44204 29961 -44198
rect 30589 -44204 30961 -44198
rect 31589 -44204 31961 -44198
rect 32589 -44204 32961 -44198
rect 33589 -44204 33961 -44198
rect 34269 -44204 34275 -43896
rect 8275 -44210 34275 -44204
rect -4275 -44498 -4228 -44496
rect 5668 -44498 5725 -44496
rect -4275 -44550 5725 -44498
rect 8615 -44236 8935 -44210
rect -49485 -44890 -49165 -44864
rect 8615 -44864 8621 -44236
rect 8929 -44864 8935 -44236
rect 8615 -44890 8935 -44864
rect 9615 -44236 9935 -44210
rect 9615 -44864 9621 -44236
rect 9929 -44864 9935 -44236
rect 9615 -44890 9935 -44864
rect 10615 -44236 10935 -44210
rect 10615 -44864 10621 -44236
rect 10929 -44864 10935 -44236
rect 10615 -44890 10935 -44864
rect 11615 -44236 11935 -44210
rect 11615 -44864 11621 -44236
rect 11929 -44864 11935 -44236
rect 11615 -44890 11935 -44864
rect 12615 -44236 12935 -44210
rect 12615 -44864 12621 -44236
rect 12929 -44864 12935 -44236
rect 12615 -44890 12935 -44864
rect 13615 -44236 13935 -44210
rect 13615 -44864 13621 -44236
rect 13929 -44864 13935 -44236
rect 13615 -44890 13935 -44864
rect 14615 -44236 14935 -44210
rect 14615 -44864 14621 -44236
rect 14929 -44864 14935 -44236
rect 14615 -44890 14935 -44864
rect 15615 -44236 15935 -44210
rect 15615 -44864 15621 -44236
rect 15929 -44864 15935 -44236
rect 15615 -44890 15935 -44864
rect 16615 -44236 16935 -44210
rect 16615 -44864 16621 -44236
rect 16929 -44864 16935 -44236
rect 16615 -44890 16935 -44864
rect 17615 -44236 17935 -44210
rect 17615 -44864 17621 -44236
rect 17929 -44864 17935 -44236
rect 17615 -44890 17935 -44864
rect 18615 -44236 18935 -44210
rect 18615 -44864 18621 -44236
rect 18929 -44864 18935 -44236
rect 18615 -44890 18935 -44864
rect 19615 -44236 19935 -44210
rect 19615 -44864 19621 -44236
rect 19929 -44864 19935 -44236
rect 19615 -44890 19935 -44864
rect 20615 -44236 20935 -44210
rect 20615 -44864 20621 -44236
rect 20929 -44864 20935 -44236
rect 20615 -44890 20935 -44864
rect 21615 -44236 21935 -44210
rect 21615 -44864 21621 -44236
rect 21929 -44864 21935 -44236
rect 21615 -44890 21935 -44864
rect 22615 -44236 22935 -44210
rect 22615 -44864 22621 -44236
rect 22929 -44864 22935 -44236
rect 22615 -44890 22935 -44864
rect 23615 -44236 23935 -44210
rect 23615 -44864 23621 -44236
rect 23929 -44864 23935 -44236
rect 23615 -44890 23935 -44864
rect 24615 -44236 24935 -44210
rect 24615 -44864 24621 -44236
rect 24929 -44864 24935 -44236
rect 24615 -44890 24935 -44864
rect 25615 -44236 25935 -44210
rect 25615 -44864 25621 -44236
rect 25929 -44864 25935 -44236
rect 25615 -44890 25935 -44864
rect 26615 -44236 26935 -44210
rect 26615 -44864 26621 -44236
rect 26929 -44864 26935 -44236
rect 26615 -44890 26935 -44864
rect 27615 -44236 27935 -44210
rect 27615 -44864 27621 -44236
rect 27929 -44864 27935 -44236
rect 27615 -44890 27935 -44864
rect 28615 -44236 28935 -44210
rect 28615 -44864 28621 -44236
rect 28929 -44864 28935 -44236
rect 28615 -44890 28935 -44864
rect 29615 -44236 29935 -44210
rect 29615 -44864 29621 -44236
rect 29929 -44864 29935 -44236
rect 29615 -44890 29935 -44864
rect 30615 -44236 30935 -44210
rect 30615 -44864 30621 -44236
rect 30929 -44864 30935 -44236
rect 30615 -44890 30935 -44864
rect 31615 -44236 31935 -44210
rect 31615 -44864 31621 -44236
rect 31929 -44864 31935 -44236
rect 31615 -44890 31935 -44864
rect 32615 -44236 32935 -44210
rect 32615 -44864 32621 -44236
rect 32929 -44864 32935 -44236
rect 32615 -44890 32935 -44864
rect 33615 -44236 33935 -44210
rect 33615 -44864 33621 -44236
rect 33929 -44864 33935 -44236
rect 33615 -44890 33935 -44864
rect -74825 -44896 -48825 -44890
rect -74825 -45204 -74819 -44896
rect -74511 -44902 -74139 -44896
rect -73511 -44902 -73139 -44896
rect -72511 -44902 -72139 -44896
rect -71511 -44902 -71139 -44896
rect -70511 -44902 -70139 -44896
rect -69511 -44902 -69139 -44896
rect -68511 -44902 -68139 -44896
rect -67511 -44902 -67139 -44896
rect -66511 -44902 -66139 -44896
rect -65511 -44902 -65139 -44896
rect -64511 -44902 -64139 -44896
rect -63511 -44902 -63139 -44896
rect -62511 -44902 -62139 -44896
rect -61511 -44902 -61139 -44896
rect -60511 -44902 -60139 -44896
rect -59511 -44902 -59139 -44896
rect -58511 -44902 -58139 -44896
rect -57511 -44902 -57139 -44896
rect -56511 -44902 -56139 -44896
rect -55511 -44902 -55139 -44896
rect -54511 -44902 -54139 -44896
rect -53511 -44902 -53139 -44896
rect -52511 -44902 -52139 -44896
rect -51511 -44902 -51139 -44896
rect -50511 -44902 -50139 -44896
rect -49511 -44902 -49139 -44896
rect -74511 -45198 -74473 -44902
rect -74177 -45198 -74139 -44902
rect -73511 -45198 -73473 -44902
rect -73177 -45198 -73139 -44902
rect -72511 -45198 -72473 -44902
rect -72177 -45198 -72139 -44902
rect -71511 -45198 -71473 -44902
rect -71177 -45198 -71139 -44902
rect -70511 -45198 -70473 -44902
rect -70177 -45198 -70139 -44902
rect -69511 -45198 -69473 -44902
rect -69177 -45198 -69139 -44902
rect -68511 -45198 -68473 -44902
rect -68177 -45198 -68139 -44902
rect -67511 -45198 -67473 -44902
rect -67177 -45198 -67139 -44902
rect -66511 -45198 -66473 -44902
rect -66177 -45198 -66139 -44902
rect -65511 -45198 -65473 -44902
rect -65177 -45198 -65139 -44902
rect -64511 -45198 -64473 -44902
rect -64177 -45198 -64139 -44902
rect -63511 -45198 -63473 -44902
rect -63177 -45198 -63139 -44902
rect -62511 -45198 -62473 -44902
rect -62177 -45198 -62139 -44902
rect -61511 -45198 -61473 -44902
rect -61177 -45198 -61139 -44902
rect -60511 -45198 -60473 -44902
rect -60177 -45198 -60139 -44902
rect -59511 -45198 -59473 -44902
rect -59177 -45198 -59139 -44902
rect -58511 -45198 -58473 -44902
rect -58177 -45198 -58139 -44902
rect -57511 -45198 -57473 -44902
rect -57177 -45198 -57139 -44902
rect -56511 -45198 -56473 -44902
rect -56177 -45198 -56139 -44902
rect -55511 -45198 -55473 -44902
rect -55177 -45198 -55139 -44902
rect -54511 -45198 -54473 -44902
rect -54177 -45198 -54139 -44902
rect -53511 -45198 -53473 -44902
rect -53177 -45198 -53139 -44902
rect -52511 -45198 -52473 -44902
rect -52177 -45198 -52139 -44902
rect -51511 -45198 -51473 -44902
rect -51177 -45198 -51139 -44902
rect -50511 -45198 -50473 -44902
rect -50177 -45198 -50139 -44902
rect -49511 -45198 -49473 -44902
rect -49177 -45198 -49139 -44902
rect -74511 -45204 -74139 -45198
rect -73511 -45204 -73139 -45198
rect -72511 -45204 -72139 -45198
rect -71511 -45204 -71139 -45198
rect -70511 -45204 -70139 -45198
rect -69511 -45204 -69139 -45198
rect -68511 -45204 -68139 -45198
rect -67511 -45204 -67139 -45198
rect -66511 -45204 -66139 -45198
rect -65511 -45204 -65139 -45198
rect -64511 -45204 -64139 -45198
rect -63511 -45204 -63139 -45198
rect -62511 -45204 -62139 -45198
rect -61511 -45204 -61139 -45198
rect -60511 -45204 -60139 -45198
rect -59511 -45204 -59139 -45198
rect -58511 -45204 -58139 -45198
rect -57511 -45204 -57139 -45198
rect -56511 -45204 -56139 -45198
rect -55511 -45204 -55139 -45198
rect -54511 -45204 -54139 -45198
rect -53511 -45204 -53139 -45198
rect -52511 -45204 -52139 -45198
rect -51511 -45204 -51139 -45198
rect -50511 -45204 -50139 -45198
rect -49511 -45204 -49139 -45198
rect -48831 -45204 -48825 -44896
rect -74825 -45210 -48825 -45204
rect 8275 -44896 34275 -44890
rect 8275 -45204 8281 -44896
rect 8589 -44902 8961 -44896
rect 9589 -44902 9961 -44896
rect 10589 -44902 10961 -44896
rect 11589 -44902 11961 -44896
rect 12589 -44902 12961 -44896
rect 13589 -44902 13961 -44896
rect 14589 -44902 14961 -44896
rect 15589 -44902 15961 -44896
rect 16589 -44902 16961 -44896
rect 17589 -44902 17961 -44896
rect 18589 -44902 18961 -44896
rect 19589 -44902 19961 -44896
rect 20589 -44902 20961 -44896
rect 21589 -44902 21961 -44896
rect 22589 -44902 22961 -44896
rect 23589 -44902 23961 -44896
rect 24589 -44902 24961 -44896
rect 25589 -44902 25961 -44896
rect 26589 -44902 26961 -44896
rect 27589 -44902 27961 -44896
rect 28589 -44902 28961 -44896
rect 29589 -44902 29961 -44896
rect 30589 -44902 30961 -44896
rect 31589 -44902 31961 -44896
rect 32589 -44902 32961 -44896
rect 33589 -44902 33961 -44896
rect 8589 -45198 8627 -44902
rect 8923 -45198 8961 -44902
rect 9589 -45198 9627 -44902
rect 9923 -45198 9961 -44902
rect 10589 -45198 10627 -44902
rect 10923 -45198 10961 -44902
rect 11589 -45198 11627 -44902
rect 11923 -45198 11961 -44902
rect 12589 -45198 12627 -44902
rect 12923 -45198 12961 -44902
rect 13589 -45198 13627 -44902
rect 13923 -45198 13961 -44902
rect 14589 -45198 14627 -44902
rect 14923 -45198 14961 -44902
rect 15589 -45198 15627 -44902
rect 15923 -45198 15961 -44902
rect 16589 -45198 16627 -44902
rect 16923 -45198 16961 -44902
rect 17589 -45198 17627 -44902
rect 17923 -45198 17961 -44902
rect 18589 -45198 18627 -44902
rect 18923 -45198 18961 -44902
rect 19589 -45198 19627 -44902
rect 19923 -45198 19961 -44902
rect 20589 -45198 20627 -44902
rect 20923 -45198 20961 -44902
rect 21589 -45198 21627 -44902
rect 21923 -45198 21961 -44902
rect 22589 -45198 22627 -44902
rect 22923 -45198 22961 -44902
rect 23589 -45198 23627 -44902
rect 23923 -45198 23961 -44902
rect 24589 -45198 24627 -44902
rect 24923 -45198 24961 -44902
rect 25589 -45198 25627 -44902
rect 25923 -45198 25961 -44902
rect 26589 -45198 26627 -44902
rect 26923 -45198 26961 -44902
rect 27589 -45198 27627 -44902
rect 27923 -45198 27961 -44902
rect 28589 -45198 28627 -44902
rect 28923 -45198 28961 -44902
rect 29589 -45198 29627 -44902
rect 29923 -45198 29961 -44902
rect 30589 -45198 30627 -44902
rect 30923 -45198 30961 -44902
rect 31589 -45198 31627 -44902
rect 31923 -45198 31961 -44902
rect 32589 -45198 32627 -44902
rect 32923 -45198 32961 -44902
rect 33589 -45198 33627 -44902
rect 33923 -45198 33961 -44902
rect 8589 -45204 8961 -45198
rect 9589 -45204 9961 -45198
rect 10589 -45204 10961 -45198
rect 11589 -45204 11961 -45198
rect 12589 -45204 12961 -45198
rect 13589 -45204 13961 -45198
rect 14589 -45204 14961 -45198
rect 15589 -45204 15961 -45198
rect 16589 -45204 16961 -45198
rect 17589 -45204 17961 -45198
rect 18589 -45204 18961 -45198
rect 19589 -45204 19961 -45198
rect 20589 -45204 20961 -45198
rect 21589 -45204 21961 -45198
rect 22589 -45204 22961 -45198
rect 23589 -45204 23961 -45198
rect 24589 -45204 24961 -45198
rect 25589 -45204 25961 -45198
rect 26589 -45204 26961 -45198
rect 27589 -45204 27961 -45198
rect 28589 -45204 28961 -45198
rect 29589 -45204 29961 -45198
rect 30589 -45204 30961 -45198
rect 31589 -45204 31961 -45198
rect 32589 -45204 32961 -45198
rect 33589 -45204 33961 -45198
rect 34269 -45204 34275 -44896
rect 8275 -45210 34275 -45204
rect -74485 -45236 -74165 -45210
rect -74485 -45864 -74479 -45236
rect -74171 -45864 -74165 -45236
rect -74485 -45890 -74165 -45864
rect -73485 -45236 -73165 -45210
rect -73485 -45864 -73479 -45236
rect -73171 -45864 -73165 -45236
rect -73485 -45890 -73165 -45864
rect -72485 -45236 -72165 -45210
rect -72485 -45864 -72479 -45236
rect -72171 -45864 -72165 -45236
rect -72485 -45890 -72165 -45864
rect -71485 -45236 -71165 -45210
rect -71485 -45864 -71479 -45236
rect -71171 -45864 -71165 -45236
rect -71485 -45890 -71165 -45864
rect -70485 -45236 -70165 -45210
rect -70485 -45864 -70479 -45236
rect -70171 -45864 -70165 -45236
rect -70485 -45890 -70165 -45864
rect -69485 -45236 -69165 -45210
rect -69485 -45864 -69479 -45236
rect -69171 -45864 -69165 -45236
rect -69485 -45890 -69165 -45864
rect -68485 -45236 -68165 -45210
rect -68485 -45864 -68479 -45236
rect -68171 -45864 -68165 -45236
rect -68485 -45890 -68165 -45864
rect -67485 -45236 -67165 -45210
rect -67485 -45864 -67479 -45236
rect -67171 -45864 -67165 -45236
rect -67485 -45890 -67165 -45864
rect -66485 -45236 -66165 -45210
rect -66485 -45864 -66479 -45236
rect -66171 -45864 -66165 -45236
rect -66485 -45890 -66165 -45864
rect -65485 -45236 -65165 -45210
rect -65485 -45864 -65479 -45236
rect -65171 -45864 -65165 -45236
rect -65485 -45890 -65165 -45864
rect -64485 -45236 -64165 -45210
rect -64485 -45864 -64479 -45236
rect -64171 -45864 -64165 -45236
rect -64485 -45890 -64165 -45864
rect -63485 -45236 -63165 -45210
rect -63485 -45864 -63479 -45236
rect -63171 -45864 -63165 -45236
rect -63485 -45890 -63165 -45864
rect -62485 -45236 -62165 -45210
rect -62485 -45864 -62479 -45236
rect -62171 -45864 -62165 -45236
rect -62485 -45890 -62165 -45864
rect -61485 -45236 -61165 -45210
rect -61485 -45864 -61479 -45236
rect -61171 -45864 -61165 -45236
rect -61485 -45890 -61165 -45864
rect -60485 -45236 -60165 -45210
rect -60485 -45864 -60479 -45236
rect -60171 -45864 -60165 -45236
rect -60485 -45890 -60165 -45864
rect -59485 -45236 -59165 -45210
rect -59485 -45864 -59479 -45236
rect -59171 -45864 -59165 -45236
rect -59485 -45890 -59165 -45864
rect -58485 -45236 -58165 -45210
rect -58485 -45864 -58479 -45236
rect -58171 -45864 -58165 -45236
rect -58485 -45890 -58165 -45864
rect -57485 -45236 -57165 -45210
rect -57485 -45864 -57479 -45236
rect -57171 -45864 -57165 -45236
rect -57485 -45890 -57165 -45864
rect -56485 -45236 -56165 -45210
rect -56485 -45864 -56479 -45236
rect -56171 -45864 -56165 -45236
rect -56485 -45890 -56165 -45864
rect -55485 -45236 -55165 -45210
rect -55485 -45864 -55479 -45236
rect -55171 -45864 -55165 -45236
rect -55485 -45890 -55165 -45864
rect -54485 -45236 -54165 -45210
rect -54485 -45864 -54479 -45236
rect -54171 -45864 -54165 -45236
rect -54485 -45890 -54165 -45864
rect -53485 -45236 -53165 -45210
rect -53485 -45864 -53479 -45236
rect -53171 -45864 -53165 -45236
rect -53485 -45890 -53165 -45864
rect -52485 -45236 -52165 -45210
rect -52485 -45864 -52479 -45236
rect -52171 -45864 -52165 -45236
rect -52485 -45890 -52165 -45864
rect -51485 -45236 -51165 -45210
rect -51485 -45864 -51479 -45236
rect -51171 -45864 -51165 -45236
rect -51485 -45890 -51165 -45864
rect -50485 -45236 -50165 -45210
rect -50485 -45864 -50479 -45236
rect -50171 -45864 -50165 -45236
rect -50485 -45890 -50165 -45864
rect -49485 -45236 -49165 -45210
rect -49485 -45864 -49479 -45236
rect -49171 -45864 -49165 -45236
rect -49485 -45890 -49165 -45864
rect 8615 -45236 8935 -45210
rect 8615 -45864 8621 -45236
rect 8929 -45864 8935 -45236
rect 8615 -45890 8935 -45864
rect 9615 -45236 9935 -45210
rect 9615 -45864 9621 -45236
rect 9929 -45864 9935 -45236
rect 9615 -45890 9935 -45864
rect 10615 -45236 10935 -45210
rect 10615 -45864 10621 -45236
rect 10929 -45864 10935 -45236
rect 10615 -45890 10935 -45864
rect 11615 -45236 11935 -45210
rect 11615 -45864 11621 -45236
rect 11929 -45864 11935 -45236
rect 11615 -45890 11935 -45864
rect 12615 -45236 12935 -45210
rect 12615 -45864 12621 -45236
rect 12929 -45864 12935 -45236
rect 12615 -45890 12935 -45864
rect 13615 -45236 13935 -45210
rect 13615 -45864 13621 -45236
rect 13929 -45864 13935 -45236
rect 13615 -45890 13935 -45864
rect 14615 -45236 14935 -45210
rect 14615 -45864 14621 -45236
rect 14929 -45864 14935 -45236
rect 14615 -45890 14935 -45864
rect 15615 -45236 15935 -45210
rect 15615 -45864 15621 -45236
rect 15929 -45864 15935 -45236
rect 15615 -45890 15935 -45864
rect 16615 -45236 16935 -45210
rect 16615 -45864 16621 -45236
rect 16929 -45864 16935 -45236
rect 16615 -45890 16935 -45864
rect 17615 -45236 17935 -45210
rect 17615 -45864 17621 -45236
rect 17929 -45864 17935 -45236
rect 17615 -45890 17935 -45864
rect 18615 -45236 18935 -45210
rect 18615 -45864 18621 -45236
rect 18929 -45864 18935 -45236
rect 18615 -45890 18935 -45864
rect 19615 -45236 19935 -45210
rect 19615 -45864 19621 -45236
rect 19929 -45864 19935 -45236
rect 19615 -45890 19935 -45864
rect 20615 -45236 20935 -45210
rect 20615 -45864 20621 -45236
rect 20929 -45864 20935 -45236
rect 20615 -45890 20935 -45864
rect 21615 -45236 21935 -45210
rect 21615 -45864 21621 -45236
rect 21929 -45864 21935 -45236
rect 21615 -45890 21935 -45864
rect 22615 -45236 22935 -45210
rect 22615 -45864 22621 -45236
rect 22929 -45864 22935 -45236
rect 22615 -45890 22935 -45864
rect 23615 -45236 23935 -45210
rect 23615 -45864 23621 -45236
rect 23929 -45864 23935 -45236
rect 23615 -45890 23935 -45864
rect 24615 -45236 24935 -45210
rect 24615 -45864 24621 -45236
rect 24929 -45864 24935 -45236
rect 24615 -45890 24935 -45864
rect 25615 -45236 25935 -45210
rect 25615 -45864 25621 -45236
rect 25929 -45864 25935 -45236
rect 25615 -45890 25935 -45864
rect 26615 -45236 26935 -45210
rect 26615 -45864 26621 -45236
rect 26929 -45864 26935 -45236
rect 26615 -45890 26935 -45864
rect 27615 -45236 27935 -45210
rect 27615 -45864 27621 -45236
rect 27929 -45864 27935 -45236
rect 27615 -45890 27935 -45864
rect 28615 -45236 28935 -45210
rect 28615 -45864 28621 -45236
rect 28929 -45864 28935 -45236
rect 28615 -45890 28935 -45864
rect 29615 -45236 29935 -45210
rect 29615 -45864 29621 -45236
rect 29929 -45864 29935 -45236
rect 29615 -45890 29935 -45864
rect 30615 -45236 30935 -45210
rect 30615 -45864 30621 -45236
rect 30929 -45864 30935 -45236
rect 30615 -45890 30935 -45864
rect 31615 -45236 31935 -45210
rect 31615 -45864 31621 -45236
rect 31929 -45864 31935 -45236
rect 31615 -45890 31935 -45864
rect 32615 -45236 32935 -45210
rect 32615 -45864 32621 -45236
rect 32929 -45864 32935 -45236
rect 32615 -45890 32935 -45864
rect 33615 -45236 33935 -45210
rect 33615 -45864 33621 -45236
rect 33929 -45864 33935 -45236
rect 33615 -45890 33935 -45864
rect -74825 -45896 -48825 -45890
rect -74825 -46204 -74819 -45896
rect -74511 -45902 -74139 -45896
rect -73511 -45902 -73139 -45896
rect -72511 -45902 -72139 -45896
rect -71511 -45902 -71139 -45896
rect -70511 -45902 -70139 -45896
rect -69511 -45902 -69139 -45896
rect -68511 -45902 -68139 -45896
rect -67511 -45902 -67139 -45896
rect -66511 -45902 -66139 -45896
rect -65511 -45902 -65139 -45896
rect -64511 -45902 -64139 -45896
rect -63511 -45902 -63139 -45896
rect -62511 -45902 -62139 -45896
rect -61511 -45902 -61139 -45896
rect -60511 -45902 -60139 -45896
rect -59511 -45902 -59139 -45896
rect -58511 -45902 -58139 -45896
rect -57511 -45902 -57139 -45896
rect -56511 -45902 -56139 -45896
rect -55511 -45902 -55139 -45896
rect -54511 -45902 -54139 -45896
rect -53511 -45902 -53139 -45896
rect -52511 -45902 -52139 -45896
rect -51511 -45902 -51139 -45896
rect -50511 -45902 -50139 -45896
rect -49511 -45902 -49139 -45896
rect -74511 -46198 -74473 -45902
rect -74177 -46198 -74139 -45902
rect -73511 -46198 -73473 -45902
rect -73177 -46198 -73139 -45902
rect -72511 -46198 -72473 -45902
rect -72177 -46198 -72139 -45902
rect -71511 -46198 -71473 -45902
rect -71177 -46198 -71139 -45902
rect -70511 -46198 -70473 -45902
rect -70177 -46198 -70139 -45902
rect -69511 -46198 -69473 -45902
rect -69177 -46198 -69139 -45902
rect -68511 -46198 -68473 -45902
rect -68177 -46198 -68139 -45902
rect -67511 -46198 -67473 -45902
rect -67177 -46198 -67139 -45902
rect -66511 -46198 -66473 -45902
rect -66177 -46198 -66139 -45902
rect -65511 -46198 -65473 -45902
rect -65177 -46198 -65139 -45902
rect -64511 -46198 -64473 -45902
rect -64177 -46198 -64139 -45902
rect -63511 -46198 -63473 -45902
rect -63177 -46198 -63139 -45902
rect -62511 -46198 -62473 -45902
rect -62177 -46198 -62139 -45902
rect -61511 -46198 -61473 -45902
rect -61177 -46198 -61139 -45902
rect -60511 -46198 -60473 -45902
rect -60177 -46198 -60139 -45902
rect -59511 -46198 -59473 -45902
rect -59177 -46198 -59139 -45902
rect -58511 -46198 -58473 -45902
rect -58177 -46198 -58139 -45902
rect -57511 -46198 -57473 -45902
rect -57177 -46198 -57139 -45902
rect -56511 -46198 -56473 -45902
rect -56177 -46198 -56139 -45902
rect -55511 -46198 -55473 -45902
rect -55177 -46198 -55139 -45902
rect -54511 -46198 -54473 -45902
rect -54177 -46198 -54139 -45902
rect -53511 -46198 -53473 -45902
rect -53177 -46198 -53139 -45902
rect -52511 -46198 -52473 -45902
rect -52177 -46198 -52139 -45902
rect -51511 -46198 -51473 -45902
rect -51177 -46198 -51139 -45902
rect -50511 -46198 -50473 -45902
rect -50177 -46198 -50139 -45902
rect -49511 -46198 -49473 -45902
rect -49177 -46198 -49139 -45902
rect -74511 -46204 -74139 -46198
rect -73511 -46204 -73139 -46198
rect -72511 -46204 -72139 -46198
rect -71511 -46204 -71139 -46198
rect -70511 -46204 -70139 -46198
rect -69511 -46204 -69139 -46198
rect -68511 -46204 -68139 -46198
rect -67511 -46204 -67139 -46198
rect -66511 -46204 -66139 -46198
rect -65511 -46204 -65139 -46198
rect -64511 -46204 -64139 -46198
rect -63511 -46204 -63139 -46198
rect -62511 -46204 -62139 -46198
rect -61511 -46204 -61139 -46198
rect -60511 -46204 -60139 -46198
rect -59511 -46204 -59139 -46198
rect -58511 -46204 -58139 -46198
rect -57511 -46204 -57139 -46198
rect -56511 -46204 -56139 -46198
rect -55511 -46204 -55139 -46198
rect -54511 -46204 -54139 -46198
rect -53511 -46204 -53139 -46198
rect -52511 -46204 -52139 -46198
rect -51511 -46204 -51139 -46198
rect -50511 -46204 -50139 -46198
rect -49511 -46204 -49139 -46198
rect -48831 -46204 -48825 -45896
rect -74825 -46210 -48825 -46204
rect 8275 -45896 34275 -45890
rect 8275 -46204 8281 -45896
rect 8589 -45902 8961 -45896
rect 9589 -45902 9961 -45896
rect 10589 -45902 10961 -45896
rect 11589 -45902 11961 -45896
rect 12589 -45902 12961 -45896
rect 13589 -45902 13961 -45896
rect 14589 -45902 14961 -45896
rect 15589 -45902 15961 -45896
rect 16589 -45902 16961 -45896
rect 17589 -45902 17961 -45896
rect 18589 -45902 18961 -45896
rect 19589 -45902 19961 -45896
rect 20589 -45902 20961 -45896
rect 21589 -45902 21961 -45896
rect 22589 -45902 22961 -45896
rect 23589 -45902 23961 -45896
rect 24589 -45902 24961 -45896
rect 25589 -45902 25961 -45896
rect 26589 -45902 26961 -45896
rect 27589 -45902 27961 -45896
rect 28589 -45902 28961 -45896
rect 29589 -45902 29961 -45896
rect 30589 -45902 30961 -45896
rect 31589 -45902 31961 -45896
rect 32589 -45902 32961 -45896
rect 33589 -45902 33961 -45896
rect 8589 -46198 8627 -45902
rect 8923 -46198 8961 -45902
rect 9589 -46198 9627 -45902
rect 9923 -46198 9961 -45902
rect 10589 -46198 10627 -45902
rect 10923 -46198 10961 -45902
rect 11589 -46198 11627 -45902
rect 11923 -46198 11961 -45902
rect 12589 -46198 12627 -45902
rect 12923 -46198 12961 -45902
rect 13589 -46198 13627 -45902
rect 13923 -46198 13961 -45902
rect 14589 -46198 14627 -45902
rect 14923 -46198 14961 -45902
rect 15589 -46198 15627 -45902
rect 15923 -46198 15961 -45902
rect 16589 -46198 16627 -45902
rect 16923 -46198 16961 -45902
rect 17589 -46198 17627 -45902
rect 17923 -46198 17961 -45902
rect 18589 -46198 18627 -45902
rect 18923 -46198 18961 -45902
rect 19589 -46198 19627 -45902
rect 19923 -46198 19961 -45902
rect 20589 -46198 20627 -45902
rect 20923 -46198 20961 -45902
rect 21589 -46198 21627 -45902
rect 21923 -46198 21961 -45902
rect 22589 -46198 22627 -45902
rect 22923 -46198 22961 -45902
rect 23589 -46198 23627 -45902
rect 23923 -46198 23961 -45902
rect 24589 -46198 24627 -45902
rect 24923 -46198 24961 -45902
rect 25589 -46198 25627 -45902
rect 25923 -46198 25961 -45902
rect 26589 -46198 26627 -45902
rect 26923 -46198 26961 -45902
rect 27589 -46198 27627 -45902
rect 27923 -46198 27961 -45902
rect 28589 -46198 28627 -45902
rect 28923 -46198 28961 -45902
rect 29589 -46198 29627 -45902
rect 29923 -46198 29961 -45902
rect 30589 -46198 30627 -45902
rect 30923 -46198 30961 -45902
rect 31589 -46198 31627 -45902
rect 31923 -46198 31961 -45902
rect 32589 -46198 32627 -45902
rect 32923 -46198 32961 -45902
rect 33589 -46198 33627 -45902
rect 33923 -46198 33961 -45902
rect 8589 -46204 8961 -46198
rect 9589 -46204 9961 -46198
rect 10589 -46204 10961 -46198
rect 11589 -46204 11961 -46198
rect 12589 -46204 12961 -46198
rect 13589 -46204 13961 -46198
rect 14589 -46204 14961 -46198
rect 15589 -46204 15961 -46198
rect 16589 -46204 16961 -46198
rect 17589 -46204 17961 -46198
rect 18589 -46204 18961 -46198
rect 19589 -46204 19961 -46198
rect 20589 -46204 20961 -46198
rect 21589 -46204 21961 -46198
rect 22589 -46204 22961 -46198
rect 23589 -46204 23961 -46198
rect 24589 -46204 24961 -46198
rect 25589 -46204 25961 -46198
rect 26589 -46204 26961 -46198
rect 27589 -46204 27961 -46198
rect 28589 -46204 28961 -46198
rect 29589 -46204 29961 -46198
rect 30589 -46204 30961 -46198
rect 31589 -46204 31961 -46198
rect 32589 -46204 32961 -46198
rect 33589 -46204 33961 -46198
rect 34269 -46204 34275 -45896
rect 8275 -46210 34275 -46204
rect -74485 -46236 -74165 -46210
rect -74485 -46544 -74479 -46236
rect -74171 -46544 -74165 -46236
rect -74485 -46550 -74165 -46544
rect -73485 -46236 -73165 -46210
rect -73485 -46544 -73479 -46236
rect -73171 -46544 -73165 -46236
rect -73485 -46550 -73165 -46544
rect -72485 -46236 -72165 -46210
rect -72485 -46544 -72479 -46236
rect -72171 -46544 -72165 -46236
rect -72485 -46550 -72165 -46544
rect -71485 -46236 -71165 -46210
rect -71485 -46544 -71479 -46236
rect -71171 -46544 -71165 -46236
rect -71485 -46550 -71165 -46544
rect -70485 -46236 -70165 -46210
rect -70485 -46544 -70479 -46236
rect -70171 -46544 -70165 -46236
rect -70485 -46550 -70165 -46544
rect -69485 -46236 -69165 -46210
rect -69485 -46544 -69479 -46236
rect -69171 -46544 -69165 -46236
rect -69485 -46550 -69165 -46544
rect -68485 -46236 -68165 -46210
rect -68485 -46544 -68479 -46236
rect -68171 -46544 -68165 -46236
rect -68485 -46550 -68165 -46544
rect -67485 -46236 -67165 -46210
rect -67485 -46544 -67479 -46236
rect -67171 -46544 -67165 -46236
rect -67485 -46550 -67165 -46544
rect -66485 -46236 -66165 -46210
rect -66485 -46544 -66479 -46236
rect -66171 -46544 -66165 -46236
rect -66485 -46550 -66165 -46544
rect -65485 -46236 -65165 -46210
rect -65485 -46544 -65479 -46236
rect -65171 -46544 -65165 -46236
rect -65485 -46550 -65165 -46544
rect -64485 -46236 -64165 -46210
rect -64485 -46544 -64479 -46236
rect -64171 -46544 -64165 -46236
rect -64485 -46550 -64165 -46544
rect -63485 -46236 -63165 -46210
rect -63485 -46544 -63479 -46236
rect -63171 -46544 -63165 -46236
rect -63485 -46550 -63165 -46544
rect -62485 -46236 -62165 -46210
rect -62485 -46544 -62479 -46236
rect -62171 -46544 -62165 -46236
rect -62485 -46550 -62165 -46544
rect -61485 -46236 -61165 -46210
rect -61485 -46544 -61479 -46236
rect -61171 -46544 -61165 -46236
rect -61485 -46550 -61165 -46544
rect -60485 -46236 -60165 -46210
rect -60485 -46544 -60479 -46236
rect -60171 -46544 -60165 -46236
rect -60485 -46550 -60165 -46544
rect -59485 -46236 -59165 -46210
rect -59485 -46544 -59479 -46236
rect -59171 -46544 -59165 -46236
rect -59485 -46550 -59165 -46544
rect -58485 -46236 -58165 -46210
rect -58485 -46544 -58479 -46236
rect -58171 -46544 -58165 -46236
rect -58485 -46550 -58165 -46544
rect -57485 -46236 -57165 -46210
rect -57485 -46544 -57479 -46236
rect -57171 -46544 -57165 -46236
rect -57485 -46550 -57165 -46544
rect -56485 -46236 -56165 -46210
rect -56485 -46544 -56479 -46236
rect -56171 -46544 -56165 -46236
rect -56485 -46550 -56165 -46544
rect -55485 -46236 -55165 -46210
rect -55485 -46544 -55479 -46236
rect -55171 -46544 -55165 -46236
rect -55485 -46550 -55165 -46544
rect -54485 -46236 -54165 -46210
rect -54485 -46544 -54479 -46236
rect -54171 -46544 -54165 -46236
rect -54485 -46550 -54165 -46544
rect -53485 -46236 -53165 -46210
rect -53485 -46544 -53479 -46236
rect -53171 -46544 -53165 -46236
rect -53485 -46550 -53165 -46544
rect -52485 -46236 -52165 -46210
rect -52485 -46544 -52479 -46236
rect -52171 -46544 -52165 -46236
rect -52485 -46550 -52165 -46544
rect -51485 -46236 -51165 -46210
rect -51485 -46544 -51479 -46236
rect -51171 -46544 -51165 -46236
rect -51485 -46550 -51165 -46544
rect -50485 -46236 -50165 -46210
rect -50485 -46544 -50479 -46236
rect -50171 -46544 -50165 -46236
rect -50485 -46550 -50165 -46544
rect -49485 -46236 -49165 -46210
rect -49485 -46544 -49479 -46236
rect -49171 -46544 -49165 -46236
rect -49485 -46550 -49165 -46544
rect 8615 -46236 8935 -46210
rect 8615 -46544 8621 -46236
rect 8929 -46544 8935 -46236
rect 8615 -46550 8935 -46544
rect 9615 -46236 9935 -46210
rect 9615 -46544 9621 -46236
rect 9929 -46544 9935 -46236
rect 9615 -46550 9935 -46544
rect 10615 -46236 10935 -46210
rect 10615 -46544 10621 -46236
rect 10929 -46544 10935 -46236
rect 10615 -46550 10935 -46544
rect 11615 -46236 11935 -46210
rect 11615 -46544 11621 -46236
rect 11929 -46544 11935 -46236
rect 11615 -46550 11935 -46544
rect 12615 -46236 12935 -46210
rect 12615 -46544 12621 -46236
rect 12929 -46544 12935 -46236
rect 12615 -46550 12935 -46544
rect 13615 -46236 13935 -46210
rect 13615 -46544 13621 -46236
rect 13929 -46544 13935 -46236
rect 13615 -46550 13935 -46544
rect 14615 -46236 14935 -46210
rect 14615 -46544 14621 -46236
rect 14929 -46544 14935 -46236
rect 14615 -46550 14935 -46544
rect 15615 -46236 15935 -46210
rect 15615 -46544 15621 -46236
rect 15929 -46544 15935 -46236
rect 15615 -46550 15935 -46544
rect 16615 -46236 16935 -46210
rect 16615 -46544 16621 -46236
rect 16929 -46544 16935 -46236
rect 16615 -46550 16935 -46544
rect 17615 -46236 17935 -46210
rect 17615 -46544 17621 -46236
rect 17929 -46544 17935 -46236
rect 17615 -46550 17935 -46544
rect 18615 -46236 18935 -46210
rect 18615 -46544 18621 -46236
rect 18929 -46544 18935 -46236
rect 18615 -46550 18935 -46544
rect 19615 -46236 19935 -46210
rect 19615 -46544 19621 -46236
rect 19929 -46544 19935 -46236
rect 19615 -46550 19935 -46544
rect 20615 -46236 20935 -46210
rect 20615 -46544 20621 -46236
rect 20929 -46544 20935 -46236
rect 20615 -46550 20935 -46544
rect 21615 -46236 21935 -46210
rect 21615 -46544 21621 -46236
rect 21929 -46544 21935 -46236
rect 21615 -46550 21935 -46544
rect 22615 -46236 22935 -46210
rect 22615 -46544 22621 -46236
rect 22929 -46544 22935 -46236
rect 22615 -46550 22935 -46544
rect 23615 -46236 23935 -46210
rect 23615 -46544 23621 -46236
rect 23929 -46544 23935 -46236
rect 23615 -46550 23935 -46544
rect 24615 -46236 24935 -46210
rect 24615 -46544 24621 -46236
rect 24929 -46544 24935 -46236
rect 24615 -46550 24935 -46544
rect 25615 -46236 25935 -46210
rect 25615 -46544 25621 -46236
rect 25929 -46544 25935 -46236
rect 25615 -46550 25935 -46544
rect 26615 -46236 26935 -46210
rect 26615 -46544 26621 -46236
rect 26929 -46544 26935 -46236
rect 26615 -46550 26935 -46544
rect 27615 -46236 27935 -46210
rect 27615 -46544 27621 -46236
rect 27929 -46544 27935 -46236
rect 27615 -46550 27935 -46544
rect 28615 -46236 28935 -46210
rect 28615 -46544 28621 -46236
rect 28929 -46544 28935 -46236
rect 28615 -46550 28935 -46544
rect 29615 -46236 29935 -46210
rect 29615 -46544 29621 -46236
rect 29929 -46544 29935 -46236
rect 29615 -46550 29935 -46544
rect 30615 -46236 30935 -46210
rect 30615 -46544 30621 -46236
rect 30929 -46544 30935 -46236
rect 30615 -46550 30935 -46544
rect 31615 -46236 31935 -46210
rect 31615 -46544 31621 -46236
rect 31929 -46544 31935 -46236
rect 31615 -46550 31935 -46544
rect 32615 -46236 32935 -46210
rect 32615 -46544 32621 -46236
rect 32929 -46544 32935 -46236
rect 32615 -46550 32935 -46544
rect 33615 -46236 33935 -46210
rect 33615 -46544 33621 -46236
rect 33929 -46544 33935 -46236
rect 33615 -46550 33935 -46544
<< via2 >>
rect -74473 38242 -74177 38538
rect -73473 38242 -73177 38538
rect -72473 38242 -72177 38538
rect -71473 38242 -71177 38538
rect -70473 38242 -70177 38538
rect -69473 38242 -69177 38538
rect -68473 38242 -68177 38538
rect -67473 38242 -67177 38538
rect -66473 38242 -66177 38538
rect -65473 38242 -65177 38538
rect -64473 38242 -64177 38538
rect -63473 38242 -63177 38538
rect -62473 38242 -62177 38538
rect -61473 38242 -61177 38538
rect -60473 38242 -60177 38538
rect -59473 38242 -59177 38538
rect 10006 38242 10302 38538
rect 11006 38242 11302 38538
rect 12006 38242 12302 38538
rect 13006 38242 13302 38538
rect 14006 38242 14302 38538
rect 15006 38242 15302 38538
rect 16006 38242 16302 38538
rect 17006 38242 17302 38538
rect 18006 38242 18302 38538
rect 19006 38242 19302 38538
rect 20006 38242 20302 38538
rect 21006 38242 21302 38538
rect 22006 38242 22302 38538
rect 23006 38242 23302 38538
rect 24006 38242 24302 38538
rect 25006 38242 25302 38538
rect 26006 38242 26302 38538
rect 27006 38242 27302 38538
rect 28006 38242 28302 38538
rect 29006 38242 29302 38538
rect 30006 38242 30302 38538
rect 31006 38242 31302 38538
rect 32006 38242 32302 38538
rect 33006 38242 33302 38538
rect 34006 38242 34302 38538
rect -74813 37902 -74517 38198
rect -74473 38172 -74177 38198
rect -74473 37928 -74447 38172
rect -74447 37928 -74203 38172
rect -74203 37928 -74177 38172
rect -74473 37902 -74177 37928
rect -74133 37902 -73517 38198
rect -73473 38172 -73177 38198
rect -73473 37928 -73447 38172
rect -73447 37928 -73203 38172
rect -73203 37928 -73177 38172
rect -73473 37902 -73177 37928
rect -73133 37902 -72517 38198
rect -72473 38172 -72177 38198
rect -72473 37928 -72447 38172
rect -72447 37928 -72203 38172
rect -72203 37928 -72177 38172
rect -72473 37902 -72177 37928
rect -72133 37902 -71517 38198
rect -71473 38172 -71177 38198
rect -71473 37928 -71447 38172
rect -71447 37928 -71203 38172
rect -71203 37928 -71177 38172
rect -71473 37902 -71177 37928
rect -71133 37902 -70517 38198
rect -70473 38172 -70177 38198
rect -70473 37928 -70447 38172
rect -70447 37928 -70203 38172
rect -70203 37928 -70177 38172
rect -70473 37902 -70177 37928
rect -70133 37902 -69517 38198
rect -69473 38172 -69177 38198
rect -69473 37928 -69447 38172
rect -69447 37928 -69203 38172
rect -69203 37928 -69177 38172
rect -69473 37902 -69177 37928
rect -69133 37902 -68517 38198
rect -68473 38172 -68177 38198
rect -68473 37928 -68447 38172
rect -68447 37928 -68203 38172
rect -68203 37928 -68177 38172
rect -68473 37902 -68177 37928
rect -68133 37902 -67517 38198
rect -67473 38172 -67177 38198
rect -67473 37928 -67447 38172
rect -67447 37928 -67203 38172
rect -67203 37928 -67177 38172
rect -67473 37902 -67177 37928
rect -67133 37902 -66517 38198
rect -66473 38172 -66177 38198
rect -66473 37928 -66447 38172
rect -66447 37928 -66203 38172
rect -66203 37928 -66177 38172
rect -66473 37902 -66177 37928
rect -66133 37902 -65517 38198
rect -65473 38172 -65177 38198
rect -65473 37928 -65447 38172
rect -65447 37928 -65203 38172
rect -65203 37928 -65177 38172
rect -65473 37902 -65177 37928
rect -65133 37902 -64517 38198
rect -64473 38172 -64177 38198
rect -64473 37928 -64447 38172
rect -64447 37928 -64203 38172
rect -64203 37928 -64177 38172
rect -64473 37902 -64177 37928
rect -64133 37902 -63517 38198
rect -63473 38172 -63177 38198
rect -63473 37928 -63447 38172
rect -63447 37928 -63203 38172
rect -63203 37928 -63177 38172
rect -63473 37902 -63177 37928
rect -63133 37902 -62517 38198
rect -62473 38172 -62177 38198
rect -62473 37928 -62447 38172
rect -62447 37928 -62203 38172
rect -62203 37928 -62177 38172
rect -62473 37902 -62177 37928
rect -62133 37902 -61517 38198
rect -61473 38172 -61177 38198
rect -61473 37928 -61447 38172
rect -61447 37928 -61203 38172
rect -61203 37928 -61177 38172
rect -61473 37902 -61177 37928
rect -61133 37902 -60517 38198
rect -60473 38172 -60177 38198
rect -60473 37928 -60447 38172
rect -60447 37928 -60203 38172
rect -60203 37928 -60177 38172
rect -60473 37902 -60177 37928
rect -60133 37902 -59517 38198
rect -59473 38172 -59177 38198
rect -59473 37928 -59447 38172
rect -59447 37928 -59203 38172
rect -59203 37928 -59177 38172
rect -59473 37902 -59177 37928
rect -59133 37902 -58837 38198
rect 9666 37902 9962 38198
rect 10006 38172 10302 38198
rect 10006 37928 10032 38172
rect 10032 37928 10276 38172
rect 10276 37928 10302 38172
rect 10006 37902 10302 37928
rect 10346 37902 10962 38198
rect 11006 38172 11302 38198
rect 11006 37928 11032 38172
rect 11032 37928 11276 38172
rect 11276 37928 11302 38172
rect 11006 37902 11302 37928
rect 11346 37902 11962 38198
rect 12006 38172 12302 38198
rect 12006 37928 12032 38172
rect 12032 37928 12276 38172
rect 12276 37928 12302 38172
rect 12006 37902 12302 37928
rect 12346 37902 12962 38198
rect 13006 38172 13302 38198
rect 13006 37928 13032 38172
rect 13032 37928 13276 38172
rect 13276 37928 13302 38172
rect 13006 37902 13302 37928
rect 13346 37902 13962 38198
rect 14006 38172 14302 38198
rect 14006 37928 14032 38172
rect 14032 37928 14276 38172
rect 14276 37928 14302 38172
rect 14006 37902 14302 37928
rect 14346 37902 14962 38198
rect 15006 38172 15302 38198
rect 15006 37928 15032 38172
rect 15032 37928 15276 38172
rect 15276 37928 15302 38172
rect 15006 37902 15302 37928
rect 15346 37902 15962 38198
rect 16006 38172 16302 38198
rect 16006 37928 16032 38172
rect 16032 37928 16276 38172
rect 16276 37928 16302 38172
rect 16006 37902 16302 37928
rect 16346 37902 16962 38198
rect 17006 38172 17302 38198
rect 17006 37928 17032 38172
rect 17032 37928 17276 38172
rect 17276 37928 17302 38172
rect 17006 37902 17302 37928
rect 17346 37902 17962 38198
rect 18006 38172 18302 38198
rect 18006 37928 18032 38172
rect 18032 37928 18276 38172
rect 18276 37928 18302 38172
rect 18006 37902 18302 37928
rect 18346 37902 18962 38198
rect 19006 38172 19302 38198
rect 19006 37928 19032 38172
rect 19032 37928 19276 38172
rect 19276 37928 19302 38172
rect 19006 37902 19302 37928
rect 19346 37902 19962 38198
rect 20006 38172 20302 38198
rect 20006 37928 20032 38172
rect 20032 37928 20276 38172
rect 20276 37928 20302 38172
rect 20006 37902 20302 37928
rect 20346 37902 20962 38198
rect 21006 38172 21302 38198
rect 21006 37928 21032 38172
rect 21032 37928 21276 38172
rect 21276 37928 21302 38172
rect 21006 37902 21302 37928
rect 21346 37902 21962 38198
rect 22006 38172 22302 38198
rect 22006 37928 22032 38172
rect 22032 37928 22276 38172
rect 22276 37928 22302 38172
rect 22006 37902 22302 37928
rect 22346 37902 22962 38198
rect 23006 38172 23302 38198
rect 23006 37928 23032 38172
rect 23032 37928 23276 38172
rect 23276 37928 23302 38172
rect 23006 37902 23302 37928
rect 23346 37902 23962 38198
rect 24006 38172 24302 38198
rect 24006 37928 24032 38172
rect 24032 37928 24276 38172
rect 24276 37928 24302 38172
rect 24006 37902 24302 37928
rect 24346 37902 24962 38198
rect 25006 38172 25302 38198
rect 25006 37928 25032 38172
rect 25032 37928 25276 38172
rect 25276 37928 25302 38172
rect 25006 37902 25302 37928
rect 25346 37902 25962 38198
rect 26006 38172 26302 38198
rect 26006 37928 26032 38172
rect 26032 37928 26276 38172
rect 26276 37928 26302 38172
rect 26006 37902 26302 37928
rect 26346 37902 26962 38198
rect 27006 38172 27302 38198
rect 27006 37928 27032 38172
rect 27032 37928 27276 38172
rect 27276 37928 27302 38172
rect 27006 37902 27302 37928
rect 27346 37902 27962 38198
rect 28006 38172 28302 38198
rect 28006 37928 28032 38172
rect 28032 37928 28276 38172
rect 28276 37928 28302 38172
rect 28006 37902 28302 37928
rect 28346 37902 28962 38198
rect 29006 38172 29302 38198
rect 29006 37928 29032 38172
rect 29032 37928 29276 38172
rect 29276 37928 29302 38172
rect 29006 37902 29302 37928
rect 29346 37902 29962 38198
rect 30006 38172 30302 38198
rect 30006 37928 30032 38172
rect 30032 37928 30276 38172
rect 30276 37928 30302 38172
rect 30006 37902 30302 37928
rect 30346 37902 30962 38198
rect 31006 38172 31302 38198
rect 31006 37928 31032 38172
rect 31032 37928 31276 38172
rect 31276 37928 31302 38172
rect 31006 37902 31302 37928
rect 31346 37902 31962 38198
rect 32006 38172 32302 38198
rect 32006 37928 32032 38172
rect 32032 37928 32276 38172
rect 32276 37928 32302 38172
rect 32006 37902 32302 37928
rect 32346 37902 32962 38198
rect 33006 38172 33302 38198
rect 33006 37928 33032 38172
rect 33032 37928 33276 38172
rect 33276 37928 33302 38172
rect 33006 37902 33302 37928
rect 33346 37902 33962 38198
rect 34006 38172 34302 38198
rect 34006 37928 34032 38172
rect 34032 37928 34276 38172
rect 34276 37928 34302 38172
rect 34006 37902 34302 37928
rect 34346 37902 34642 38198
rect -74473 37242 -74177 37858
rect -73473 37242 -73177 37858
rect -72473 37242 -72177 37858
rect -71473 37242 -71177 37858
rect -70473 37242 -70177 37858
rect -69473 37242 -69177 37858
rect -68473 37242 -68177 37858
rect -67473 37242 -67177 37858
rect -66473 37242 -66177 37858
rect -65473 37242 -65177 37858
rect -64473 37242 -64177 37858
rect -63473 37242 -63177 37858
rect -62473 37242 -62177 37858
rect -61473 37242 -61177 37858
rect -60473 37242 -60177 37858
rect -59473 37242 -59177 37858
rect 10006 37242 10302 37858
rect 11006 37242 11302 37858
rect 12006 37242 12302 37858
rect 13006 37242 13302 37858
rect 14006 37242 14302 37858
rect 15006 37242 15302 37858
rect 16006 37242 16302 37858
rect 17006 37242 17302 37858
rect 18006 37242 18302 37858
rect 19006 37242 19302 37858
rect 20006 37242 20302 37858
rect 21006 37242 21302 37858
rect 22006 37242 22302 37858
rect 23006 37242 23302 37858
rect 24006 37242 24302 37858
rect 25006 37242 25302 37858
rect 26006 37242 26302 37858
rect 27006 37242 27302 37858
rect 28006 37242 28302 37858
rect 29006 37242 29302 37858
rect 30006 37242 30302 37858
rect 31006 37242 31302 37858
rect 32006 37242 32302 37858
rect 33006 37242 33302 37858
rect 34006 37242 34302 37858
rect -74813 36902 -74517 37198
rect -74473 37172 -74177 37198
rect -74473 36928 -74447 37172
rect -74447 36928 -74203 37172
rect -74203 36928 -74177 37172
rect -74473 36902 -74177 36928
rect -74133 36902 -73517 37198
rect -73473 37172 -73177 37198
rect -73473 36928 -73447 37172
rect -73447 36928 -73203 37172
rect -73203 36928 -73177 37172
rect -73473 36902 -73177 36928
rect -73133 36902 -72517 37198
rect -72473 37172 -72177 37198
rect -72473 36928 -72447 37172
rect -72447 36928 -72203 37172
rect -72203 36928 -72177 37172
rect -72473 36902 -72177 36928
rect -72133 36902 -71517 37198
rect -71473 37172 -71177 37198
rect -71473 36928 -71447 37172
rect -71447 36928 -71203 37172
rect -71203 36928 -71177 37172
rect -71473 36902 -71177 36928
rect -71133 36902 -70517 37198
rect -70473 37172 -70177 37198
rect -70473 36928 -70447 37172
rect -70447 36928 -70203 37172
rect -70203 36928 -70177 37172
rect -70473 36902 -70177 36928
rect -70133 36902 -69517 37198
rect -69473 37172 -69177 37198
rect -69473 36928 -69447 37172
rect -69447 36928 -69203 37172
rect -69203 36928 -69177 37172
rect -69473 36902 -69177 36928
rect -69133 36902 -68517 37198
rect -68473 37172 -68177 37198
rect -68473 36928 -68447 37172
rect -68447 36928 -68203 37172
rect -68203 36928 -68177 37172
rect -68473 36902 -68177 36928
rect -68133 36902 -67517 37198
rect -67473 37172 -67177 37198
rect -67473 36928 -67447 37172
rect -67447 36928 -67203 37172
rect -67203 36928 -67177 37172
rect -67473 36902 -67177 36928
rect -67133 36902 -66517 37198
rect -66473 37172 -66177 37198
rect -66473 36928 -66447 37172
rect -66447 36928 -66203 37172
rect -66203 36928 -66177 37172
rect -66473 36902 -66177 36928
rect -66133 36902 -65517 37198
rect -65473 37172 -65177 37198
rect -65473 36928 -65447 37172
rect -65447 36928 -65203 37172
rect -65203 36928 -65177 37172
rect -65473 36902 -65177 36928
rect -65133 36902 -64517 37198
rect -64473 37172 -64177 37198
rect -64473 36928 -64447 37172
rect -64447 36928 -64203 37172
rect -64203 36928 -64177 37172
rect -64473 36902 -64177 36928
rect -64133 36902 -63517 37198
rect -63473 37172 -63177 37198
rect -63473 36928 -63447 37172
rect -63447 36928 -63203 37172
rect -63203 36928 -63177 37172
rect -63473 36902 -63177 36928
rect -63133 36902 -62517 37198
rect -62473 37172 -62177 37198
rect -62473 36928 -62447 37172
rect -62447 36928 -62203 37172
rect -62203 36928 -62177 37172
rect -62473 36902 -62177 36928
rect -62133 36902 -61517 37198
rect -61473 37172 -61177 37198
rect -61473 36928 -61447 37172
rect -61447 36928 -61203 37172
rect -61203 36928 -61177 37172
rect -61473 36902 -61177 36928
rect -61133 36902 -60517 37198
rect -60473 37172 -60177 37198
rect -60473 36928 -60447 37172
rect -60447 36928 -60203 37172
rect -60203 36928 -60177 37172
rect -60473 36902 -60177 36928
rect -60133 36902 -59517 37198
rect -59473 37172 -59177 37198
rect -59473 36928 -59447 37172
rect -59447 36928 -59203 37172
rect -59203 36928 -59177 37172
rect -59473 36902 -59177 36928
rect -59133 36902 -58837 37198
rect 9666 36902 9962 37198
rect 10006 37172 10302 37198
rect 10006 36928 10032 37172
rect 10032 36928 10276 37172
rect 10276 36928 10302 37172
rect 10006 36902 10302 36928
rect 10346 36902 10962 37198
rect 11006 37172 11302 37198
rect 11006 36928 11032 37172
rect 11032 36928 11276 37172
rect 11276 36928 11302 37172
rect 11006 36902 11302 36928
rect 11346 36902 11962 37198
rect 12006 37172 12302 37198
rect 12006 36928 12032 37172
rect 12032 36928 12276 37172
rect 12276 36928 12302 37172
rect 12006 36902 12302 36928
rect 12346 36902 12962 37198
rect 13006 37172 13302 37198
rect 13006 36928 13032 37172
rect 13032 36928 13276 37172
rect 13276 36928 13302 37172
rect 13006 36902 13302 36928
rect 13346 36902 13962 37198
rect 14006 37172 14302 37198
rect 14006 36928 14032 37172
rect 14032 36928 14276 37172
rect 14276 36928 14302 37172
rect 14006 36902 14302 36928
rect 14346 36902 14962 37198
rect 15006 37172 15302 37198
rect 15006 36928 15032 37172
rect 15032 36928 15276 37172
rect 15276 36928 15302 37172
rect 15006 36902 15302 36928
rect 15346 36902 15962 37198
rect 16006 37172 16302 37198
rect 16006 36928 16032 37172
rect 16032 36928 16276 37172
rect 16276 36928 16302 37172
rect 16006 36902 16302 36928
rect 16346 36902 16962 37198
rect 17006 37172 17302 37198
rect 17006 36928 17032 37172
rect 17032 36928 17276 37172
rect 17276 36928 17302 37172
rect 17006 36902 17302 36928
rect 17346 36902 17962 37198
rect 18006 37172 18302 37198
rect 18006 36928 18032 37172
rect 18032 36928 18276 37172
rect 18276 36928 18302 37172
rect 18006 36902 18302 36928
rect 18346 36902 18962 37198
rect 19006 37172 19302 37198
rect 19006 36928 19032 37172
rect 19032 36928 19276 37172
rect 19276 36928 19302 37172
rect 19006 36902 19302 36928
rect 19346 36902 19962 37198
rect 20006 37172 20302 37198
rect 20006 36928 20032 37172
rect 20032 36928 20276 37172
rect 20276 36928 20302 37172
rect 20006 36902 20302 36928
rect 20346 36902 20962 37198
rect 21006 37172 21302 37198
rect 21006 36928 21032 37172
rect 21032 36928 21276 37172
rect 21276 36928 21302 37172
rect 21006 36902 21302 36928
rect 21346 36902 21962 37198
rect 22006 37172 22302 37198
rect 22006 36928 22032 37172
rect 22032 36928 22276 37172
rect 22276 36928 22302 37172
rect 22006 36902 22302 36928
rect 22346 36902 22962 37198
rect 23006 37172 23302 37198
rect 23006 36928 23032 37172
rect 23032 36928 23276 37172
rect 23276 36928 23302 37172
rect 23006 36902 23302 36928
rect 23346 36902 23962 37198
rect 24006 37172 24302 37198
rect 24006 36928 24032 37172
rect 24032 36928 24276 37172
rect 24276 36928 24302 37172
rect 24006 36902 24302 36928
rect 24346 36902 24962 37198
rect 25006 37172 25302 37198
rect 25006 36928 25032 37172
rect 25032 36928 25276 37172
rect 25276 36928 25302 37172
rect 25006 36902 25302 36928
rect 25346 36902 25962 37198
rect 26006 37172 26302 37198
rect 26006 36928 26032 37172
rect 26032 36928 26276 37172
rect 26276 36928 26302 37172
rect 26006 36902 26302 36928
rect 26346 36902 26962 37198
rect 27006 37172 27302 37198
rect 27006 36928 27032 37172
rect 27032 36928 27276 37172
rect 27276 36928 27302 37172
rect 27006 36902 27302 36928
rect 27346 36902 27962 37198
rect 28006 37172 28302 37198
rect 28006 36928 28032 37172
rect 28032 36928 28276 37172
rect 28276 36928 28302 37172
rect 28006 36902 28302 36928
rect 28346 36902 28962 37198
rect 29006 37172 29302 37198
rect 29006 36928 29032 37172
rect 29032 36928 29276 37172
rect 29276 36928 29302 37172
rect 29006 36902 29302 36928
rect 29346 36902 29962 37198
rect 30006 37172 30302 37198
rect 30006 36928 30032 37172
rect 30032 36928 30276 37172
rect 30276 36928 30302 37172
rect 30006 36902 30302 36928
rect 30346 36902 30962 37198
rect 31006 37172 31302 37198
rect 31006 36928 31032 37172
rect 31032 36928 31276 37172
rect 31276 36928 31302 37172
rect 31006 36902 31302 36928
rect 31346 36902 31962 37198
rect 32006 37172 32302 37198
rect 32006 36928 32032 37172
rect 32032 36928 32276 37172
rect 32276 36928 32302 37172
rect 32006 36902 32302 36928
rect 32346 36902 32962 37198
rect 33006 37172 33302 37198
rect 33006 36928 33032 37172
rect 33032 36928 33276 37172
rect 33276 36928 33302 37172
rect 33006 36902 33302 36928
rect 33346 36902 33962 37198
rect 34006 37172 34302 37198
rect 34006 36928 34032 37172
rect 34032 36928 34276 37172
rect 34276 36928 34302 37172
rect 34006 36902 34302 36928
rect 34346 36902 34642 37198
rect -74473 36242 -74177 36858
rect -73473 36242 -73177 36858
rect -72473 36242 -72177 36858
rect -71473 36242 -71177 36858
rect -70473 36242 -70177 36858
rect -69473 36242 -69177 36858
rect -68473 36242 -68177 36858
rect -67473 36242 -67177 36858
rect -66473 36242 -66177 36858
rect -65473 36242 -65177 36858
rect -64473 36242 -64177 36858
rect -63473 36242 -63177 36858
rect -62473 36242 -62177 36858
rect -61473 36242 -61177 36858
rect -60473 36242 -60177 36858
rect -59473 36242 -59177 36858
rect 10006 36242 10302 36858
rect 11006 36242 11302 36858
rect 12006 36242 12302 36858
rect 13006 36242 13302 36858
rect 14006 36242 14302 36858
rect 15006 36242 15302 36858
rect 16006 36242 16302 36858
rect 17006 36242 17302 36858
rect 18006 36242 18302 36858
rect 19006 36242 19302 36858
rect 20006 36242 20302 36858
rect 21006 36242 21302 36858
rect 22006 36242 22302 36858
rect 23006 36242 23302 36858
rect 24006 36242 24302 36858
rect 25006 36242 25302 36858
rect 26006 36242 26302 36858
rect 27006 36242 27302 36858
rect 28006 36242 28302 36858
rect 29006 36242 29302 36858
rect 30006 36242 30302 36858
rect 31006 36242 31302 36858
rect 32006 36242 32302 36858
rect 33006 36242 33302 36858
rect 34006 36242 34302 36858
rect -74813 35902 -74517 36198
rect -74473 36172 -74177 36198
rect -74473 35928 -74447 36172
rect -74447 35928 -74203 36172
rect -74203 35928 -74177 36172
rect -74473 35902 -74177 35928
rect -74133 35902 -73517 36198
rect -73473 36172 -73177 36198
rect -73473 35928 -73447 36172
rect -73447 35928 -73203 36172
rect -73203 35928 -73177 36172
rect -73473 35902 -73177 35928
rect -73133 35902 -72517 36198
rect -72473 36172 -72177 36198
rect -72473 35928 -72447 36172
rect -72447 35928 -72203 36172
rect -72203 35928 -72177 36172
rect -72473 35902 -72177 35928
rect -72133 35902 -71517 36198
rect -71473 36172 -71177 36198
rect -71473 35928 -71447 36172
rect -71447 35928 -71203 36172
rect -71203 35928 -71177 36172
rect -71473 35902 -71177 35928
rect -71133 35902 -70517 36198
rect -70473 36172 -70177 36198
rect -70473 35928 -70447 36172
rect -70447 35928 -70203 36172
rect -70203 35928 -70177 36172
rect -70473 35902 -70177 35928
rect -70133 35902 -69517 36198
rect -69473 36172 -69177 36198
rect -69473 35928 -69447 36172
rect -69447 35928 -69203 36172
rect -69203 35928 -69177 36172
rect -69473 35902 -69177 35928
rect -69133 35902 -68517 36198
rect -68473 36172 -68177 36198
rect -68473 35928 -68447 36172
rect -68447 35928 -68203 36172
rect -68203 35928 -68177 36172
rect -68473 35902 -68177 35928
rect -68133 35902 -67517 36198
rect -67473 36172 -67177 36198
rect -67473 35928 -67447 36172
rect -67447 35928 -67203 36172
rect -67203 35928 -67177 36172
rect -67473 35902 -67177 35928
rect -67133 35902 -66517 36198
rect -66473 36172 -66177 36198
rect -66473 35928 -66447 36172
rect -66447 35928 -66203 36172
rect -66203 35928 -66177 36172
rect -66473 35902 -66177 35928
rect -66133 35902 -65517 36198
rect -65473 36172 -65177 36198
rect -65473 35928 -65447 36172
rect -65447 35928 -65203 36172
rect -65203 35928 -65177 36172
rect -65473 35902 -65177 35928
rect -65133 35902 -64517 36198
rect -64473 36172 -64177 36198
rect -64473 35928 -64447 36172
rect -64447 35928 -64203 36172
rect -64203 35928 -64177 36172
rect -64473 35902 -64177 35928
rect -64133 35902 -63517 36198
rect -63473 36172 -63177 36198
rect -63473 35928 -63447 36172
rect -63447 35928 -63203 36172
rect -63203 35928 -63177 36172
rect -63473 35902 -63177 35928
rect -63133 35902 -62517 36198
rect -62473 36172 -62177 36198
rect -62473 35928 -62447 36172
rect -62447 35928 -62203 36172
rect -62203 35928 -62177 36172
rect -62473 35902 -62177 35928
rect -62133 35902 -61517 36198
rect -61473 36172 -61177 36198
rect -61473 35928 -61447 36172
rect -61447 35928 -61203 36172
rect -61203 35928 -61177 36172
rect -61473 35902 -61177 35928
rect -61133 35902 -60517 36198
rect -60473 36172 -60177 36198
rect -60473 35928 -60447 36172
rect -60447 35928 -60203 36172
rect -60203 35928 -60177 36172
rect -60473 35902 -60177 35928
rect -60133 35902 -59517 36198
rect -59473 36172 -59177 36198
rect -59473 35928 -59447 36172
rect -59447 35928 -59203 36172
rect -59203 35928 -59177 36172
rect -59473 35902 -59177 35928
rect -59133 35902 -58837 36198
rect 9666 35902 9962 36198
rect 10006 36172 10302 36198
rect 10006 35928 10032 36172
rect 10032 35928 10276 36172
rect 10276 35928 10302 36172
rect 10006 35902 10302 35928
rect 10346 35902 10962 36198
rect 11006 36172 11302 36198
rect 11006 35928 11032 36172
rect 11032 35928 11276 36172
rect 11276 35928 11302 36172
rect 11006 35902 11302 35928
rect 11346 35902 11962 36198
rect 12006 36172 12302 36198
rect 12006 35928 12032 36172
rect 12032 35928 12276 36172
rect 12276 35928 12302 36172
rect 12006 35902 12302 35928
rect 12346 35902 12962 36198
rect 13006 36172 13302 36198
rect 13006 35928 13032 36172
rect 13032 35928 13276 36172
rect 13276 35928 13302 36172
rect 13006 35902 13302 35928
rect 13346 35902 13962 36198
rect 14006 36172 14302 36198
rect 14006 35928 14032 36172
rect 14032 35928 14276 36172
rect 14276 35928 14302 36172
rect 14006 35902 14302 35928
rect 14346 35902 14962 36198
rect 15006 36172 15302 36198
rect 15006 35928 15032 36172
rect 15032 35928 15276 36172
rect 15276 35928 15302 36172
rect 15006 35902 15302 35928
rect 15346 35902 15962 36198
rect 16006 36172 16302 36198
rect 16006 35928 16032 36172
rect 16032 35928 16276 36172
rect 16276 35928 16302 36172
rect 16006 35902 16302 35928
rect 16346 35902 16962 36198
rect 17006 36172 17302 36198
rect 17006 35928 17032 36172
rect 17032 35928 17276 36172
rect 17276 35928 17302 36172
rect 17006 35902 17302 35928
rect 17346 35902 17962 36198
rect 18006 36172 18302 36198
rect 18006 35928 18032 36172
rect 18032 35928 18276 36172
rect 18276 35928 18302 36172
rect 18006 35902 18302 35928
rect 18346 35902 18962 36198
rect 19006 36172 19302 36198
rect 19006 35928 19032 36172
rect 19032 35928 19276 36172
rect 19276 35928 19302 36172
rect 19006 35902 19302 35928
rect 19346 35902 19962 36198
rect 20006 36172 20302 36198
rect 20006 35928 20032 36172
rect 20032 35928 20276 36172
rect 20276 35928 20302 36172
rect 20006 35902 20302 35928
rect 20346 35902 20962 36198
rect 21006 36172 21302 36198
rect 21006 35928 21032 36172
rect 21032 35928 21276 36172
rect 21276 35928 21302 36172
rect 21006 35902 21302 35928
rect 21346 35902 21962 36198
rect 22006 36172 22302 36198
rect 22006 35928 22032 36172
rect 22032 35928 22276 36172
rect 22276 35928 22302 36172
rect 22006 35902 22302 35928
rect 22346 35902 22962 36198
rect 23006 36172 23302 36198
rect 23006 35928 23032 36172
rect 23032 35928 23276 36172
rect 23276 35928 23302 36172
rect 23006 35902 23302 35928
rect 23346 35902 23962 36198
rect 24006 36172 24302 36198
rect 24006 35928 24032 36172
rect 24032 35928 24276 36172
rect 24276 35928 24302 36172
rect 24006 35902 24302 35928
rect 24346 35902 24962 36198
rect 25006 36172 25302 36198
rect 25006 35928 25032 36172
rect 25032 35928 25276 36172
rect 25276 35928 25302 36172
rect 25006 35902 25302 35928
rect 25346 35902 25962 36198
rect 26006 36172 26302 36198
rect 26006 35928 26032 36172
rect 26032 35928 26276 36172
rect 26276 35928 26302 36172
rect 26006 35902 26302 35928
rect 26346 35902 26962 36198
rect 27006 36172 27302 36198
rect 27006 35928 27032 36172
rect 27032 35928 27276 36172
rect 27276 35928 27302 36172
rect 27006 35902 27302 35928
rect 27346 35902 27962 36198
rect 28006 36172 28302 36198
rect 28006 35928 28032 36172
rect 28032 35928 28276 36172
rect 28276 35928 28302 36172
rect 28006 35902 28302 35928
rect 28346 35902 28962 36198
rect 29006 36172 29302 36198
rect 29006 35928 29032 36172
rect 29032 35928 29276 36172
rect 29276 35928 29302 36172
rect 29006 35902 29302 35928
rect 29346 35902 29962 36198
rect 30006 36172 30302 36198
rect 30006 35928 30032 36172
rect 30032 35928 30276 36172
rect 30276 35928 30302 36172
rect 30006 35902 30302 35928
rect 30346 35902 30962 36198
rect 31006 36172 31302 36198
rect 31006 35928 31032 36172
rect 31032 35928 31276 36172
rect 31276 35928 31302 36172
rect 31006 35902 31302 35928
rect 31346 35902 31962 36198
rect 32006 36172 32302 36198
rect 32006 35928 32032 36172
rect 32032 35928 32276 36172
rect 32276 35928 32302 36172
rect 32006 35902 32302 35928
rect 32346 35902 32962 36198
rect 33006 36172 33302 36198
rect 33006 35928 33032 36172
rect 33032 35928 33276 36172
rect 33276 35928 33302 36172
rect 33006 35902 33302 35928
rect 33346 35902 33962 36198
rect 34006 36172 34302 36198
rect 34006 35928 34032 36172
rect 34032 35928 34276 36172
rect 34276 35928 34302 36172
rect 34006 35902 34302 35928
rect 34346 35902 34642 36198
rect -74473 35242 -74177 35858
rect -73473 35242 -73177 35858
rect -72473 35242 -72177 35858
rect -71473 35242 -71177 35858
rect -70473 35242 -70177 35858
rect -69473 35242 -69177 35858
rect -68473 35242 -68177 35858
rect -67473 35242 -67177 35858
rect -66473 35242 -66177 35858
rect -65473 35242 -65177 35858
rect -64473 35242 -64177 35858
rect -63473 35242 -63177 35858
rect -62473 35242 -62177 35858
rect -61473 35242 -61177 35858
rect -60473 35242 -60177 35858
rect -59473 35242 -59177 35858
rect 10006 35242 10302 35858
rect 11006 35242 11302 35858
rect 12006 35242 12302 35858
rect 13006 35242 13302 35858
rect 14006 35242 14302 35858
rect 15006 35242 15302 35858
rect 16006 35242 16302 35858
rect 17006 35242 17302 35858
rect 18006 35242 18302 35858
rect 19006 35242 19302 35858
rect 20006 35242 20302 35858
rect 21006 35242 21302 35858
rect 22006 35242 22302 35858
rect 23006 35242 23302 35858
rect 24006 35242 24302 35858
rect 25006 35242 25302 35858
rect 26006 35242 26302 35858
rect 27006 35242 27302 35858
rect 28006 35242 28302 35858
rect 29006 35242 29302 35858
rect 30006 35242 30302 35858
rect 31006 35242 31302 35858
rect 32006 35242 32302 35858
rect 33006 35242 33302 35858
rect 34006 35242 34302 35858
rect -74813 34902 -74517 35198
rect -74473 35172 -74177 35198
rect -74473 34928 -74447 35172
rect -74447 34928 -74203 35172
rect -74203 34928 -74177 35172
rect -74473 34902 -74177 34928
rect -74133 34902 -73517 35198
rect -73473 35172 -73177 35198
rect -73473 34928 -73447 35172
rect -73447 34928 -73203 35172
rect -73203 34928 -73177 35172
rect -73473 34902 -73177 34928
rect -73133 34902 -72517 35198
rect -72473 35172 -72177 35198
rect -72473 34928 -72447 35172
rect -72447 34928 -72203 35172
rect -72203 34928 -72177 35172
rect -72473 34902 -72177 34928
rect -72133 34902 -71517 35198
rect -71473 35172 -71177 35198
rect -71473 34928 -71447 35172
rect -71447 34928 -71203 35172
rect -71203 34928 -71177 35172
rect -71473 34902 -71177 34928
rect -71133 34902 -70517 35198
rect -70473 35172 -70177 35198
rect -70473 34928 -70447 35172
rect -70447 34928 -70203 35172
rect -70203 34928 -70177 35172
rect -70473 34902 -70177 34928
rect -70133 34902 -69517 35198
rect -69473 35172 -69177 35198
rect -69473 34928 -69447 35172
rect -69447 34928 -69203 35172
rect -69203 34928 -69177 35172
rect -69473 34902 -69177 34928
rect -69133 34902 -68517 35198
rect -68473 35172 -68177 35198
rect -68473 34928 -68447 35172
rect -68447 34928 -68203 35172
rect -68203 34928 -68177 35172
rect -68473 34902 -68177 34928
rect -68133 34902 -67517 35198
rect -67473 35172 -67177 35198
rect -67473 34928 -67447 35172
rect -67447 34928 -67203 35172
rect -67203 34928 -67177 35172
rect -67473 34902 -67177 34928
rect -67133 34902 -66517 35198
rect -66473 35172 -66177 35198
rect -66473 34928 -66447 35172
rect -66447 34928 -66203 35172
rect -66203 34928 -66177 35172
rect -66473 34902 -66177 34928
rect -66133 34902 -65517 35198
rect -65473 35172 -65177 35198
rect -65473 34928 -65447 35172
rect -65447 34928 -65203 35172
rect -65203 34928 -65177 35172
rect -65473 34902 -65177 34928
rect -65133 34902 -64517 35198
rect -64473 35172 -64177 35198
rect -64473 34928 -64447 35172
rect -64447 34928 -64203 35172
rect -64203 34928 -64177 35172
rect -64473 34902 -64177 34928
rect -64133 34902 -63517 35198
rect -63473 35172 -63177 35198
rect -63473 34928 -63447 35172
rect -63447 34928 -63203 35172
rect -63203 34928 -63177 35172
rect -63473 34902 -63177 34928
rect -63133 34902 -62517 35198
rect -62473 35172 -62177 35198
rect -62473 34928 -62447 35172
rect -62447 34928 -62203 35172
rect -62203 34928 -62177 35172
rect -62473 34902 -62177 34928
rect -62133 34902 -61517 35198
rect -61473 35172 -61177 35198
rect -61473 34928 -61447 35172
rect -61447 34928 -61203 35172
rect -61203 34928 -61177 35172
rect -61473 34902 -61177 34928
rect -61133 34902 -60517 35198
rect -60473 35172 -60177 35198
rect -60473 34928 -60447 35172
rect -60447 34928 -60203 35172
rect -60203 34928 -60177 35172
rect -60473 34902 -60177 34928
rect -60133 34902 -59517 35198
rect -59473 35172 -59177 35198
rect -59473 34928 -59447 35172
rect -59447 34928 -59203 35172
rect -59203 34928 -59177 35172
rect -59473 34902 -59177 34928
rect -59133 34902 -58837 35198
rect 9666 34902 9962 35198
rect 10006 35172 10302 35198
rect 10006 34928 10032 35172
rect 10032 34928 10276 35172
rect 10276 34928 10302 35172
rect 10006 34902 10302 34928
rect 10346 34902 10962 35198
rect 11006 35172 11302 35198
rect 11006 34928 11032 35172
rect 11032 34928 11276 35172
rect 11276 34928 11302 35172
rect 11006 34902 11302 34928
rect 11346 34902 11962 35198
rect 12006 35172 12302 35198
rect 12006 34928 12032 35172
rect 12032 34928 12276 35172
rect 12276 34928 12302 35172
rect 12006 34902 12302 34928
rect 12346 34902 12962 35198
rect 13006 35172 13302 35198
rect 13006 34928 13032 35172
rect 13032 34928 13276 35172
rect 13276 34928 13302 35172
rect 13006 34902 13302 34928
rect 13346 34902 13962 35198
rect 14006 35172 14302 35198
rect 14006 34928 14032 35172
rect 14032 34928 14276 35172
rect 14276 34928 14302 35172
rect 14006 34902 14302 34928
rect 14346 34902 14962 35198
rect 15006 35172 15302 35198
rect 15006 34928 15032 35172
rect 15032 34928 15276 35172
rect 15276 34928 15302 35172
rect 15006 34902 15302 34928
rect 15346 34902 15962 35198
rect 16006 35172 16302 35198
rect 16006 34928 16032 35172
rect 16032 34928 16276 35172
rect 16276 34928 16302 35172
rect 16006 34902 16302 34928
rect 16346 34902 16962 35198
rect 17006 35172 17302 35198
rect 17006 34928 17032 35172
rect 17032 34928 17276 35172
rect 17276 34928 17302 35172
rect 17006 34902 17302 34928
rect 17346 34902 17962 35198
rect 18006 35172 18302 35198
rect 18006 34928 18032 35172
rect 18032 34928 18276 35172
rect 18276 34928 18302 35172
rect 18006 34902 18302 34928
rect 18346 34902 18962 35198
rect 19006 35172 19302 35198
rect 19006 34928 19032 35172
rect 19032 34928 19276 35172
rect 19276 34928 19302 35172
rect 19006 34902 19302 34928
rect 19346 34902 19962 35198
rect 20006 35172 20302 35198
rect 20006 34928 20032 35172
rect 20032 34928 20276 35172
rect 20276 34928 20302 35172
rect 20006 34902 20302 34928
rect 20346 34902 20962 35198
rect 21006 35172 21302 35198
rect 21006 34928 21032 35172
rect 21032 34928 21276 35172
rect 21276 34928 21302 35172
rect 21006 34902 21302 34928
rect 21346 34902 21962 35198
rect 22006 35172 22302 35198
rect 22006 34928 22032 35172
rect 22032 34928 22276 35172
rect 22276 34928 22302 35172
rect 22006 34902 22302 34928
rect 22346 34902 22962 35198
rect 23006 35172 23302 35198
rect 23006 34928 23032 35172
rect 23032 34928 23276 35172
rect 23276 34928 23302 35172
rect 23006 34902 23302 34928
rect 23346 34902 23962 35198
rect 24006 35172 24302 35198
rect 24006 34928 24032 35172
rect 24032 34928 24276 35172
rect 24276 34928 24302 35172
rect 24006 34902 24302 34928
rect 24346 34902 24962 35198
rect 25006 35172 25302 35198
rect 25006 34928 25032 35172
rect 25032 34928 25276 35172
rect 25276 34928 25302 35172
rect 25006 34902 25302 34928
rect 25346 34902 25962 35198
rect 26006 35172 26302 35198
rect 26006 34928 26032 35172
rect 26032 34928 26276 35172
rect 26276 34928 26302 35172
rect 26006 34902 26302 34928
rect 26346 34902 26962 35198
rect 27006 35172 27302 35198
rect 27006 34928 27032 35172
rect 27032 34928 27276 35172
rect 27276 34928 27302 35172
rect 27006 34902 27302 34928
rect 27346 34902 27962 35198
rect 28006 35172 28302 35198
rect 28006 34928 28032 35172
rect 28032 34928 28276 35172
rect 28276 34928 28302 35172
rect 28006 34902 28302 34928
rect 28346 34902 28962 35198
rect 29006 35172 29302 35198
rect 29006 34928 29032 35172
rect 29032 34928 29276 35172
rect 29276 34928 29302 35172
rect 29006 34902 29302 34928
rect 29346 34902 29962 35198
rect 30006 35172 30302 35198
rect 30006 34928 30032 35172
rect 30032 34928 30276 35172
rect 30276 34928 30302 35172
rect 30006 34902 30302 34928
rect 30346 34902 30962 35198
rect 31006 35172 31302 35198
rect 31006 34928 31032 35172
rect 31032 34928 31276 35172
rect 31276 34928 31302 35172
rect 31006 34902 31302 34928
rect 31346 34902 31962 35198
rect 32006 35172 32302 35198
rect 32006 34928 32032 35172
rect 32032 34928 32276 35172
rect 32276 34928 32302 35172
rect 32006 34902 32302 34928
rect 32346 34902 32962 35198
rect 33006 35172 33302 35198
rect 33006 34928 33032 35172
rect 33032 34928 33276 35172
rect 33276 34928 33302 35172
rect 33006 34902 33302 34928
rect 33346 34902 33962 35198
rect 34006 35172 34302 35198
rect 34006 34928 34032 35172
rect 34032 34928 34276 35172
rect 34276 34928 34302 35172
rect 34006 34902 34302 34928
rect 34346 34902 34642 35198
rect -74473 34242 -74177 34858
rect -73473 34242 -73177 34858
rect -72473 34242 -72177 34858
rect -71473 34242 -71177 34858
rect -70473 34242 -70177 34858
rect -69473 34242 -69177 34858
rect -68473 34242 -68177 34858
rect -67473 34242 -67177 34858
rect -66473 34242 -66177 34858
rect -65473 34242 -65177 34858
rect -64473 34242 -64177 34858
rect -63473 34242 -63177 34858
rect -62473 34242 -62177 34858
rect -61473 34242 -61177 34858
rect -60473 34242 -60177 34858
rect -59473 34242 -59177 34858
rect 10006 34242 10302 34858
rect 11006 34242 11302 34858
rect 12006 34242 12302 34858
rect 13006 34242 13302 34858
rect 14006 34242 14302 34858
rect 15006 34242 15302 34858
rect 16006 34242 16302 34858
rect 17006 34242 17302 34858
rect 18006 34242 18302 34858
rect 19006 34242 19302 34858
rect 20006 34242 20302 34858
rect 21006 34242 21302 34858
rect 22006 34242 22302 34858
rect 23006 34242 23302 34858
rect 24006 34242 24302 34858
rect 25006 34242 25302 34858
rect 26006 34242 26302 34858
rect 27006 34242 27302 34858
rect 28006 34242 28302 34858
rect 29006 34242 29302 34858
rect 30006 34242 30302 34858
rect 31006 34242 31302 34858
rect 32006 34242 32302 34858
rect 33006 34242 33302 34858
rect 34006 34242 34302 34858
rect -74813 33902 -74517 34198
rect -74473 34172 -74177 34198
rect -74473 33928 -74447 34172
rect -74447 33928 -74203 34172
rect -74203 33928 -74177 34172
rect -74473 33902 -74177 33928
rect -74133 33902 -73517 34198
rect -73473 34172 -73177 34198
rect -73473 33928 -73447 34172
rect -73447 33928 -73203 34172
rect -73203 33928 -73177 34172
rect -73473 33902 -73177 33928
rect -73133 33902 -72517 34198
rect -72473 34172 -72177 34198
rect -72473 33928 -72447 34172
rect -72447 33928 -72203 34172
rect -72203 33928 -72177 34172
rect -72473 33902 -72177 33928
rect -72133 33902 -71517 34198
rect -71473 34172 -71177 34198
rect -71473 33928 -71447 34172
rect -71447 33928 -71203 34172
rect -71203 33928 -71177 34172
rect -71473 33902 -71177 33928
rect -71133 33902 -70517 34198
rect -70473 34172 -70177 34198
rect -70473 33928 -70447 34172
rect -70447 33928 -70203 34172
rect -70203 33928 -70177 34172
rect -70473 33902 -70177 33928
rect -70133 33902 -69517 34198
rect -69473 34172 -69177 34198
rect -69473 33928 -69447 34172
rect -69447 33928 -69203 34172
rect -69203 33928 -69177 34172
rect -69473 33902 -69177 33928
rect -69133 33902 -68517 34198
rect -68473 34172 -68177 34198
rect -68473 33928 -68447 34172
rect -68447 33928 -68203 34172
rect -68203 33928 -68177 34172
rect -68473 33902 -68177 33928
rect -68133 33902 -67517 34198
rect -67473 34172 -67177 34198
rect -67473 33928 -67447 34172
rect -67447 33928 -67203 34172
rect -67203 33928 -67177 34172
rect -67473 33902 -67177 33928
rect -67133 33902 -66517 34198
rect -66473 34172 -66177 34198
rect -66473 33928 -66447 34172
rect -66447 33928 -66203 34172
rect -66203 33928 -66177 34172
rect -66473 33902 -66177 33928
rect -66133 33902 -65517 34198
rect -65473 34172 -65177 34198
rect -65473 33928 -65447 34172
rect -65447 33928 -65203 34172
rect -65203 33928 -65177 34172
rect -65473 33902 -65177 33928
rect -65133 33902 -64517 34198
rect -64473 34172 -64177 34198
rect -64473 33928 -64447 34172
rect -64447 33928 -64203 34172
rect -64203 33928 -64177 34172
rect -64473 33902 -64177 33928
rect -64133 33902 -63517 34198
rect -63473 34172 -63177 34198
rect -63473 33928 -63447 34172
rect -63447 33928 -63203 34172
rect -63203 33928 -63177 34172
rect -63473 33902 -63177 33928
rect -63133 33902 -62517 34198
rect -62473 34172 -62177 34198
rect -62473 33928 -62447 34172
rect -62447 33928 -62203 34172
rect -62203 33928 -62177 34172
rect -62473 33902 -62177 33928
rect -62133 33902 -61517 34198
rect -61473 34172 -61177 34198
rect -61473 33928 -61447 34172
rect -61447 33928 -61203 34172
rect -61203 33928 -61177 34172
rect -61473 33902 -61177 33928
rect -61133 33902 -60517 34198
rect -60473 34172 -60177 34198
rect -60473 33928 -60447 34172
rect -60447 33928 -60203 34172
rect -60203 33928 -60177 34172
rect -60473 33902 -60177 33928
rect -60133 33902 -59517 34198
rect -59473 34172 -59177 34198
rect -59473 33928 -59447 34172
rect -59447 33928 -59203 34172
rect -59203 33928 -59177 34172
rect -59473 33902 -59177 33928
rect -59133 33902 -58837 34198
rect -74473 33242 -74177 33858
rect -73473 33242 -73177 33858
rect -72473 33242 -72177 33858
rect -71473 33242 -71177 33858
rect -70473 33242 -70177 33858
rect -69473 33242 -69177 33858
rect -68473 33242 -68177 33858
rect -67473 33242 -67177 33858
rect -66473 33242 -66177 33858
rect -65473 33242 -65177 33858
rect -64473 33242 -64177 33858
rect -63473 33242 -63177 33858
rect -62473 33242 -62177 33858
rect -61473 33242 -61177 33858
rect -60473 33242 -60177 33858
rect -59473 33242 -59177 33858
rect -50428 33548 -48852 34164
rect 2919 33548 4495 34164
rect 9666 33902 9962 34198
rect 10006 34172 10302 34198
rect 10006 33928 10032 34172
rect 10032 33928 10276 34172
rect 10276 33928 10302 34172
rect 10006 33902 10302 33928
rect 10346 33902 10962 34198
rect 11006 34172 11302 34198
rect 11006 33928 11032 34172
rect 11032 33928 11276 34172
rect 11276 33928 11302 34172
rect 11006 33902 11302 33928
rect 11346 33902 11962 34198
rect 12006 34172 12302 34198
rect 12006 33928 12032 34172
rect 12032 33928 12276 34172
rect 12276 33928 12302 34172
rect 12006 33902 12302 33928
rect 12346 33902 12962 34198
rect 13006 34172 13302 34198
rect 13006 33928 13032 34172
rect 13032 33928 13276 34172
rect 13276 33928 13302 34172
rect 13006 33902 13302 33928
rect 13346 33902 13962 34198
rect 14006 34172 14302 34198
rect 14006 33928 14032 34172
rect 14032 33928 14276 34172
rect 14276 33928 14302 34172
rect 14006 33902 14302 33928
rect 14346 33902 14962 34198
rect 15006 34172 15302 34198
rect 15006 33928 15032 34172
rect 15032 33928 15276 34172
rect 15276 33928 15302 34172
rect 15006 33902 15302 33928
rect 15346 33902 15962 34198
rect 16006 34172 16302 34198
rect 16006 33928 16032 34172
rect 16032 33928 16276 34172
rect 16276 33928 16302 34172
rect 16006 33902 16302 33928
rect 16346 33902 16962 34198
rect 17006 34172 17302 34198
rect 17006 33928 17032 34172
rect 17032 33928 17276 34172
rect 17276 33928 17302 34172
rect 17006 33902 17302 33928
rect 17346 33902 17962 34198
rect 18006 34172 18302 34198
rect 18006 33928 18032 34172
rect 18032 33928 18276 34172
rect 18276 33928 18302 34172
rect 18006 33902 18302 33928
rect 18346 33902 18962 34198
rect 19006 34172 19302 34198
rect 19006 33928 19032 34172
rect 19032 33928 19276 34172
rect 19276 33928 19302 34172
rect 19006 33902 19302 33928
rect 19346 33902 19962 34198
rect 20006 34172 20302 34198
rect 20006 33928 20032 34172
rect 20032 33928 20276 34172
rect 20276 33928 20302 34172
rect 20006 33902 20302 33928
rect 20346 33902 20962 34198
rect 21006 34172 21302 34198
rect 21006 33928 21032 34172
rect 21032 33928 21276 34172
rect 21276 33928 21302 34172
rect 21006 33902 21302 33928
rect 21346 33902 21962 34198
rect 22006 34172 22302 34198
rect 22006 33928 22032 34172
rect 22032 33928 22276 34172
rect 22276 33928 22302 34172
rect 22006 33902 22302 33928
rect 22346 33902 22962 34198
rect 23006 34172 23302 34198
rect 23006 33928 23032 34172
rect 23032 33928 23276 34172
rect 23276 33928 23302 34172
rect 23006 33902 23302 33928
rect 23346 33902 23962 34198
rect 24006 34172 24302 34198
rect 24006 33928 24032 34172
rect 24032 33928 24276 34172
rect 24276 33928 24302 34172
rect 24006 33902 24302 33928
rect 24346 33902 24962 34198
rect 25006 34172 25302 34198
rect 25006 33928 25032 34172
rect 25032 33928 25276 34172
rect 25276 33928 25302 34172
rect 25006 33902 25302 33928
rect 25346 33902 25962 34198
rect 26006 34172 26302 34198
rect 26006 33928 26032 34172
rect 26032 33928 26276 34172
rect 26276 33928 26302 34172
rect 26006 33902 26302 33928
rect 26346 33902 26962 34198
rect 27006 34172 27302 34198
rect 27006 33928 27032 34172
rect 27032 33928 27276 34172
rect 27276 33928 27302 34172
rect 27006 33902 27302 33928
rect 27346 33902 27962 34198
rect 28006 34172 28302 34198
rect 28006 33928 28032 34172
rect 28032 33928 28276 34172
rect 28276 33928 28302 34172
rect 28006 33902 28302 33928
rect 28346 33902 28962 34198
rect 29006 34172 29302 34198
rect 29006 33928 29032 34172
rect 29032 33928 29276 34172
rect 29276 33928 29302 34172
rect 29006 33902 29302 33928
rect 29346 33902 29962 34198
rect 30006 34172 30302 34198
rect 30006 33928 30032 34172
rect 30032 33928 30276 34172
rect 30276 33928 30302 34172
rect 30006 33902 30302 33928
rect 30346 33902 30962 34198
rect 31006 34172 31302 34198
rect 31006 33928 31032 34172
rect 31032 33928 31276 34172
rect 31276 33928 31302 34172
rect 31006 33902 31302 33928
rect 31346 33902 31962 34198
rect 32006 34172 32302 34198
rect 32006 33928 32032 34172
rect 32032 33928 32276 34172
rect 32276 33928 32302 34172
rect 32006 33902 32302 33928
rect 32346 33902 32962 34198
rect 33006 34172 33302 34198
rect 33006 33928 33032 34172
rect 33032 33928 33276 34172
rect 33276 33928 33302 34172
rect 33006 33902 33302 33928
rect 33346 33902 33962 34198
rect 34006 34172 34302 34198
rect 34006 33928 34032 34172
rect 34032 33928 34276 34172
rect 34276 33928 34302 34172
rect 34006 33902 34302 33928
rect 34346 33902 34642 34198
rect -74813 32902 -74517 33198
rect -74473 33172 -74177 33198
rect -74473 32928 -74447 33172
rect -74447 32928 -74203 33172
rect -74203 32928 -74177 33172
rect -74473 32902 -74177 32928
rect -74133 32902 -73517 33198
rect -73473 33172 -73177 33198
rect -73473 32928 -73447 33172
rect -73447 32928 -73203 33172
rect -73203 32928 -73177 33172
rect -73473 32902 -73177 32928
rect -73133 32902 -72517 33198
rect -72473 33172 -72177 33198
rect -72473 32928 -72447 33172
rect -72447 32928 -72203 33172
rect -72203 32928 -72177 33172
rect -72473 32902 -72177 32928
rect -72133 32902 -71517 33198
rect -71473 33172 -71177 33198
rect -71473 32928 -71447 33172
rect -71447 32928 -71203 33172
rect -71203 32928 -71177 33172
rect -71473 32902 -71177 32928
rect -71133 32902 -70517 33198
rect -70473 33172 -70177 33198
rect -70473 32928 -70447 33172
rect -70447 32928 -70203 33172
rect -70203 32928 -70177 33172
rect -70473 32902 -70177 32928
rect -70133 32902 -69517 33198
rect -69473 33172 -69177 33198
rect -69473 32928 -69447 33172
rect -69447 32928 -69203 33172
rect -69203 32928 -69177 33172
rect -69473 32902 -69177 32928
rect -69133 32902 -68517 33198
rect -68473 33172 -68177 33198
rect -68473 32928 -68447 33172
rect -68447 32928 -68203 33172
rect -68203 32928 -68177 33172
rect -68473 32902 -68177 32928
rect -68133 32902 -67517 33198
rect -67473 33172 -67177 33198
rect -67473 32928 -67447 33172
rect -67447 32928 -67203 33172
rect -67203 32928 -67177 33172
rect -67473 32902 -67177 32928
rect -67133 32902 -66517 33198
rect -66473 33172 -66177 33198
rect -66473 32928 -66447 33172
rect -66447 32928 -66203 33172
rect -66203 32928 -66177 33172
rect -66473 32902 -66177 32928
rect -66133 32902 -65517 33198
rect -65473 33172 -65177 33198
rect -65473 32928 -65447 33172
rect -65447 32928 -65203 33172
rect -65203 32928 -65177 33172
rect -65473 32902 -65177 32928
rect -65133 32902 -64517 33198
rect -64473 33172 -64177 33198
rect -64473 32928 -64447 33172
rect -64447 32928 -64203 33172
rect -64203 32928 -64177 33172
rect -64473 32902 -64177 32928
rect -64133 32902 -63517 33198
rect -63473 33172 -63177 33198
rect -63473 32928 -63447 33172
rect -63447 32928 -63203 33172
rect -63203 32928 -63177 33172
rect -63473 32902 -63177 32928
rect -63133 32902 -62517 33198
rect -62473 33172 -62177 33198
rect -62473 32928 -62447 33172
rect -62447 32928 -62203 33172
rect -62203 32928 -62177 33172
rect -62473 32902 -62177 32928
rect -62133 32902 -61517 33198
rect -61473 33172 -61177 33198
rect -61473 32928 -61447 33172
rect -61447 32928 -61203 33172
rect -61203 32928 -61177 33172
rect -61473 32902 -61177 32928
rect -61133 32902 -60517 33198
rect -60473 33172 -60177 33198
rect -60473 32928 -60447 33172
rect -60447 32928 -60203 33172
rect -60203 32928 -60177 33172
rect -60473 32902 -60177 32928
rect -60133 32902 -59517 33198
rect -59473 33172 -59177 33198
rect -59473 32928 -59447 33172
rect -59447 32928 -59203 33172
rect -59203 32928 -59177 33172
rect -59473 32902 -59177 32928
rect -59133 32902 -58837 33198
rect -74473 32242 -74177 32858
rect -73473 32242 -73177 32858
rect -72473 32242 -72177 32858
rect -71473 32242 -71177 32858
rect -70473 32242 -70177 32858
rect -69473 32242 -69177 32858
rect -68473 32242 -68177 32858
rect -67473 32242 -67177 32858
rect -66473 32242 -66177 32858
rect -65473 32242 -65177 32858
rect -64473 32242 -64177 32858
rect -63473 32242 -63177 32858
rect -62473 32242 -62177 32858
rect -61473 32242 -61177 32858
rect -60473 32242 -60177 32858
rect -59473 32242 -59177 32858
rect -50955 32965 -50579 32967
rect -50955 32593 -50951 32965
rect -50951 32593 -50579 32965
rect -50955 32591 -50579 32593
rect 10006 33242 10302 33858
rect 11006 33242 11302 33858
rect 12006 33242 12302 33858
rect 13006 33242 13302 33858
rect 14006 33242 14302 33858
rect 15006 33242 15302 33858
rect 16006 33242 16302 33858
rect 17006 33242 17302 33858
rect 18006 33242 18302 33858
rect 19006 33242 19302 33858
rect 20006 33242 20302 33858
rect 21006 33242 21302 33858
rect 22006 33242 22302 33858
rect 23006 33242 23302 33858
rect 24006 33242 24302 33858
rect 25006 33242 25302 33858
rect 26006 33242 26302 33858
rect 27006 33242 27302 33858
rect 28006 33242 28302 33858
rect 29006 33242 29302 33858
rect 30006 33242 30302 33858
rect 31006 33242 31302 33858
rect 32006 33242 32302 33858
rect 33006 33242 33302 33858
rect 34006 33242 34302 33858
rect 9666 32902 9962 33198
rect 10006 33172 10302 33198
rect 10006 32928 10032 33172
rect 10032 32928 10276 33172
rect 10276 32928 10302 33172
rect 10006 32902 10302 32928
rect 10346 32902 10962 33198
rect 11006 33172 11302 33198
rect 11006 32928 11032 33172
rect 11032 32928 11276 33172
rect 11276 32928 11302 33172
rect 11006 32902 11302 32928
rect 11346 32902 11962 33198
rect 12006 33172 12302 33198
rect 12006 32928 12032 33172
rect 12032 32928 12276 33172
rect 12276 32928 12302 33172
rect 12006 32902 12302 32928
rect 12346 32902 12962 33198
rect 13006 33172 13302 33198
rect 13006 32928 13032 33172
rect 13032 32928 13276 33172
rect 13276 32928 13302 33172
rect 13006 32902 13302 32928
rect 13346 32902 13962 33198
rect 14006 33172 14302 33198
rect 14006 32928 14032 33172
rect 14032 32928 14276 33172
rect 14276 32928 14302 33172
rect 14006 32902 14302 32928
rect 14346 32902 14962 33198
rect 15006 33172 15302 33198
rect 15006 32928 15032 33172
rect 15032 32928 15276 33172
rect 15276 32928 15302 33172
rect 15006 32902 15302 32928
rect 15346 32902 15962 33198
rect 16006 33172 16302 33198
rect 16006 32928 16032 33172
rect 16032 32928 16276 33172
rect 16276 32928 16302 33172
rect 16006 32902 16302 32928
rect 16346 32902 16962 33198
rect 17006 33172 17302 33198
rect 17006 32928 17032 33172
rect 17032 32928 17276 33172
rect 17276 32928 17302 33172
rect 17006 32902 17302 32928
rect 17346 32902 17962 33198
rect 18006 33172 18302 33198
rect 18006 32928 18032 33172
rect 18032 32928 18276 33172
rect 18276 32928 18302 33172
rect 18006 32902 18302 32928
rect 18346 32902 18962 33198
rect 19006 33172 19302 33198
rect 19006 32928 19032 33172
rect 19032 32928 19276 33172
rect 19276 32928 19302 33172
rect 19006 32902 19302 32928
rect 19346 32902 19962 33198
rect 20006 33172 20302 33198
rect 20006 32928 20032 33172
rect 20032 32928 20276 33172
rect 20276 32928 20302 33172
rect 20006 32902 20302 32928
rect 20346 32902 20962 33198
rect 21006 33172 21302 33198
rect 21006 32928 21032 33172
rect 21032 32928 21276 33172
rect 21276 32928 21302 33172
rect 21006 32902 21302 32928
rect 21346 32902 21962 33198
rect 22006 33172 22302 33198
rect 22006 32928 22032 33172
rect 22032 32928 22276 33172
rect 22276 32928 22302 33172
rect 22006 32902 22302 32928
rect 22346 32902 22962 33198
rect 23006 33172 23302 33198
rect 23006 32928 23032 33172
rect 23032 32928 23276 33172
rect 23276 32928 23302 33172
rect 23006 32902 23302 32928
rect 23346 32902 23962 33198
rect 24006 33172 24302 33198
rect 24006 32928 24032 33172
rect 24032 32928 24276 33172
rect 24276 32928 24302 33172
rect 24006 32902 24302 32928
rect 24346 32902 24962 33198
rect 25006 33172 25302 33198
rect 25006 32928 25032 33172
rect 25032 32928 25276 33172
rect 25276 32928 25302 33172
rect 25006 32902 25302 32928
rect 25346 32902 25962 33198
rect 26006 33172 26302 33198
rect 26006 32928 26032 33172
rect 26032 32928 26276 33172
rect 26276 32928 26302 33172
rect 26006 32902 26302 32928
rect 26346 32902 26962 33198
rect 27006 33172 27302 33198
rect 27006 32928 27032 33172
rect 27032 32928 27276 33172
rect 27276 32928 27302 33172
rect 27006 32902 27302 32928
rect 27346 32902 27962 33198
rect 28006 33172 28302 33198
rect 28006 32928 28032 33172
rect 28032 32928 28276 33172
rect 28276 32928 28302 33172
rect 28006 32902 28302 32928
rect 28346 32902 28962 33198
rect 29006 33172 29302 33198
rect 29006 32928 29032 33172
rect 29032 32928 29276 33172
rect 29276 32928 29302 33172
rect 29006 32902 29302 32928
rect 29346 32902 29962 33198
rect 30006 33172 30302 33198
rect 30006 32928 30032 33172
rect 30032 32928 30276 33172
rect 30276 32928 30302 33172
rect 30006 32902 30302 32928
rect 30346 32902 30962 33198
rect 31006 33172 31302 33198
rect 31006 32928 31032 33172
rect 31032 32928 31276 33172
rect 31276 32928 31302 33172
rect 31006 32902 31302 32928
rect 31346 32902 31962 33198
rect 32006 33172 32302 33198
rect 32006 32928 32032 33172
rect 32032 32928 32276 33172
rect 32276 32928 32302 33172
rect 32006 32902 32302 32928
rect 32346 32902 32962 33198
rect 33006 33172 33302 33198
rect 33006 32928 33032 33172
rect 33032 32928 33276 33172
rect 33276 32928 33302 33172
rect 33006 32902 33302 32928
rect 33346 32902 33962 33198
rect 34006 33172 34302 33198
rect 34006 32928 34032 33172
rect 34032 32928 34276 33172
rect 34276 32928 34302 33172
rect 34006 32902 34302 32928
rect 34346 32902 34642 33198
rect -74813 31902 -74517 32198
rect -74473 32172 -74177 32198
rect -74473 31928 -74447 32172
rect -74447 31928 -74203 32172
rect -74203 31928 -74177 32172
rect -74473 31902 -74177 31928
rect -74133 31902 -73517 32198
rect -73473 32172 -73177 32198
rect -73473 31928 -73447 32172
rect -73447 31928 -73203 32172
rect -73203 31928 -73177 32172
rect -73473 31902 -73177 31928
rect -73133 31902 -72517 32198
rect -72473 32172 -72177 32198
rect -72473 31928 -72447 32172
rect -72447 31928 -72203 32172
rect -72203 31928 -72177 32172
rect -72473 31902 -72177 31928
rect -72133 31902 -71517 32198
rect -71473 32172 -71177 32198
rect -71473 31928 -71447 32172
rect -71447 31928 -71203 32172
rect -71203 31928 -71177 32172
rect -71473 31902 -71177 31928
rect -71133 31902 -70517 32198
rect -70473 32172 -70177 32198
rect -70473 31928 -70447 32172
rect -70447 31928 -70203 32172
rect -70203 31928 -70177 32172
rect -70473 31902 -70177 31928
rect -70133 31902 -69517 32198
rect -69473 32172 -69177 32198
rect -69473 31928 -69447 32172
rect -69447 31928 -69203 32172
rect -69203 31928 -69177 32172
rect -69473 31902 -69177 31928
rect -69133 31902 -68517 32198
rect -68473 32172 -68177 32198
rect -68473 31928 -68447 32172
rect -68447 31928 -68203 32172
rect -68203 31928 -68177 32172
rect -68473 31902 -68177 31928
rect -68133 31902 -67517 32198
rect -67473 32172 -67177 32198
rect -67473 31928 -67447 32172
rect -67447 31928 -67203 32172
rect -67203 31928 -67177 32172
rect -67473 31902 -67177 31928
rect -67133 31902 -66517 32198
rect -66473 32172 -66177 32198
rect -66473 31928 -66447 32172
rect -66447 31928 -66203 32172
rect -66203 31928 -66177 32172
rect -66473 31902 -66177 31928
rect -66133 31902 -65517 32198
rect -65473 32172 -65177 32198
rect -65473 31928 -65447 32172
rect -65447 31928 -65203 32172
rect -65203 31928 -65177 32172
rect -65473 31902 -65177 31928
rect -65133 31902 -64517 32198
rect -64473 32172 -64177 32198
rect -64473 31928 -64447 32172
rect -64447 31928 -64203 32172
rect -64203 31928 -64177 32172
rect -64473 31902 -64177 31928
rect -64133 31902 -63517 32198
rect -63473 32172 -63177 32198
rect -63473 31928 -63447 32172
rect -63447 31928 -63203 32172
rect -63203 31928 -63177 32172
rect -63473 31902 -63177 31928
rect -63133 31902 -62517 32198
rect -62473 32172 -62177 32198
rect -62473 31928 -62447 32172
rect -62447 31928 -62203 32172
rect -62203 31928 -62177 32172
rect -62473 31902 -62177 31928
rect -62133 31902 -61517 32198
rect -61473 32172 -61177 32198
rect -61473 31928 -61447 32172
rect -61447 31928 -61203 32172
rect -61203 31928 -61177 32172
rect -61473 31902 -61177 31928
rect -61133 31902 -60517 32198
rect -60473 32172 -60177 32198
rect -60473 31928 -60447 32172
rect -60447 31928 -60203 32172
rect -60203 31928 -60177 32172
rect -60473 31902 -60177 31928
rect -60133 31902 -59517 32198
rect -59473 32172 -59177 32198
rect -59473 31928 -59447 32172
rect -59447 31928 -59203 32172
rect -59203 31928 -59177 32172
rect -59473 31902 -59177 31928
rect -59133 31902 -58837 32198
rect -74473 31242 -74177 31858
rect -73473 31242 -73177 31858
rect -72473 31242 -72177 31858
rect -71473 31242 -71177 31858
rect -70473 31242 -70177 31858
rect -69473 31242 -69177 31858
rect -68473 31242 -68177 31858
rect -67473 31242 -67177 31858
rect -66473 31242 -66177 31858
rect -65473 31242 -65177 31858
rect -64473 31242 -64177 31858
rect -63473 31242 -63177 31858
rect -62473 31242 -62177 31858
rect -61473 31242 -61177 31858
rect -60473 31242 -60177 31858
rect -59473 31242 -59177 31858
rect -74813 30902 -74517 31198
rect -74473 31172 -74177 31198
rect -74473 30928 -74447 31172
rect -74447 30928 -74203 31172
rect -74203 30928 -74177 31172
rect -74473 30902 -74177 30928
rect -74133 30902 -73517 31198
rect -73473 31172 -73177 31198
rect -73473 30928 -73447 31172
rect -73447 30928 -73203 31172
rect -73203 30928 -73177 31172
rect -73473 30902 -73177 30928
rect -73133 30902 -72517 31198
rect -72473 31172 -72177 31198
rect -72473 30928 -72447 31172
rect -72447 30928 -72203 31172
rect -72203 30928 -72177 31172
rect -72473 30902 -72177 30928
rect -72133 30902 -71517 31198
rect -71473 31172 -71177 31198
rect -71473 30928 -71447 31172
rect -71447 30928 -71203 31172
rect -71203 30928 -71177 31172
rect -71473 30902 -71177 30928
rect -71133 30902 -70517 31198
rect -70473 31172 -70177 31198
rect -70473 30928 -70447 31172
rect -70447 30928 -70203 31172
rect -70203 30928 -70177 31172
rect -70473 30902 -70177 30928
rect -70133 30902 -69517 31198
rect -69473 31172 -69177 31198
rect -69473 30928 -69447 31172
rect -69447 30928 -69203 31172
rect -69203 30928 -69177 31172
rect -69473 30902 -69177 30928
rect -69133 30902 -68517 31198
rect -68473 31172 -68177 31198
rect -68473 30928 -68447 31172
rect -68447 30928 -68203 31172
rect -68203 30928 -68177 31172
rect -68473 30902 -68177 30928
rect -68133 30902 -67517 31198
rect -67473 31172 -67177 31198
rect -67473 30928 -67447 31172
rect -67447 30928 -67203 31172
rect -67203 30928 -67177 31172
rect -67473 30902 -67177 30928
rect -67133 30902 -66517 31198
rect -66473 31172 -66177 31198
rect -66473 30928 -66447 31172
rect -66447 30928 -66203 31172
rect -66203 30928 -66177 31172
rect -66473 30902 -66177 30928
rect -66133 30902 -65517 31198
rect -65473 31172 -65177 31198
rect -65473 30928 -65447 31172
rect -65447 30928 -65203 31172
rect -65203 30928 -65177 31172
rect -65473 30902 -65177 30928
rect -65133 30902 -64517 31198
rect -64473 31172 -64177 31198
rect -64473 30928 -64447 31172
rect -64447 30928 -64203 31172
rect -64203 30928 -64177 31172
rect -64473 30902 -64177 30928
rect -64133 30902 -63517 31198
rect -63473 31172 -63177 31198
rect -63473 30928 -63447 31172
rect -63447 30928 -63203 31172
rect -63203 30928 -63177 31172
rect -63473 30902 -63177 30928
rect -63133 30902 -62517 31198
rect -62473 31172 -62177 31198
rect -62473 30928 -62447 31172
rect -62447 30928 -62203 31172
rect -62203 30928 -62177 31172
rect -62473 30902 -62177 30928
rect -62133 30902 -61517 31198
rect -61473 31172 -61177 31198
rect -61473 30928 -61447 31172
rect -61447 30928 -61203 31172
rect -61203 30928 -61177 31172
rect -61473 30902 -61177 30928
rect -61133 30902 -60517 31198
rect -60473 31172 -60177 31198
rect -60473 30928 -60447 31172
rect -60447 30928 -60203 31172
rect -60203 30928 -60177 31172
rect -60473 30902 -60177 30928
rect -60133 30902 -59517 31198
rect -59473 31172 -59177 31198
rect -59473 30928 -59447 31172
rect -59447 30928 -59203 31172
rect -59203 30928 -59177 31172
rect -59473 30902 -59177 30928
rect -59133 30902 -58837 31198
rect -74473 30242 -74177 30858
rect -73473 30242 -73177 30858
rect -72473 30242 -72177 30858
rect -71473 30242 -71177 30858
rect -70473 30242 -70177 30858
rect -69473 30242 -69177 30858
rect -68473 30242 -68177 30858
rect -67473 30242 -67177 30858
rect -66473 30242 -66177 30858
rect -65473 30242 -65177 30858
rect -64473 30242 -64177 30858
rect -63473 30242 -63177 30858
rect -62473 30242 -62177 30858
rect -61473 30242 -61177 30858
rect -60473 30242 -60177 30858
rect -59473 30242 -59177 30858
rect -74813 29902 -74517 30198
rect -74473 30172 -74177 30198
rect -74473 29928 -74447 30172
rect -74447 29928 -74203 30172
rect -74203 29928 -74177 30172
rect -74473 29902 -74177 29928
rect -74133 29902 -73517 30198
rect -73473 30172 -73177 30198
rect -73473 29928 -73447 30172
rect -73447 29928 -73203 30172
rect -73203 29928 -73177 30172
rect -73473 29902 -73177 29928
rect -73133 29902 -72517 30198
rect -72473 30172 -72177 30198
rect -72473 29928 -72447 30172
rect -72447 29928 -72203 30172
rect -72203 29928 -72177 30172
rect -72473 29902 -72177 29928
rect -72133 29902 -71517 30198
rect -71473 30172 -71177 30198
rect -71473 29928 -71447 30172
rect -71447 29928 -71203 30172
rect -71203 29928 -71177 30172
rect -71473 29902 -71177 29928
rect -71133 29902 -70517 30198
rect -70473 30172 -70177 30198
rect -70473 29928 -70447 30172
rect -70447 29928 -70203 30172
rect -70203 29928 -70177 30172
rect -70473 29902 -70177 29928
rect -70133 29902 -69517 30198
rect -69473 30172 -69177 30198
rect -69473 29928 -69447 30172
rect -69447 29928 -69203 30172
rect -69203 29928 -69177 30172
rect -69473 29902 -69177 29928
rect -69133 29902 -68517 30198
rect -68473 30172 -68177 30198
rect -68473 29928 -68447 30172
rect -68447 29928 -68203 30172
rect -68203 29928 -68177 30172
rect -68473 29902 -68177 29928
rect -68133 29902 -67517 30198
rect -67473 30172 -67177 30198
rect -67473 29928 -67447 30172
rect -67447 29928 -67203 30172
rect -67203 29928 -67177 30172
rect -67473 29902 -67177 29928
rect -67133 29902 -66517 30198
rect -66473 30172 -66177 30198
rect -66473 29928 -66447 30172
rect -66447 29928 -66203 30172
rect -66203 29928 -66177 30172
rect -66473 29902 -66177 29928
rect -66133 29902 -65517 30198
rect -65473 30172 -65177 30198
rect -65473 29928 -65447 30172
rect -65447 29928 -65203 30172
rect -65203 29928 -65177 30172
rect -65473 29902 -65177 29928
rect -65133 29902 -64517 30198
rect -64473 30172 -64177 30198
rect -64473 29928 -64447 30172
rect -64447 29928 -64203 30172
rect -64203 29928 -64177 30172
rect -64473 29902 -64177 29928
rect -64133 29902 -63517 30198
rect -63473 30172 -63177 30198
rect -63473 29928 -63447 30172
rect -63447 29928 -63203 30172
rect -63203 29928 -63177 30172
rect -63473 29902 -63177 29928
rect -63133 29902 -62517 30198
rect -62473 30172 -62177 30198
rect -62473 29928 -62447 30172
rect -62447 29928 -62203 30172
rect -62203 29928 -62177 30172
rect -62473 29902 -62177 29928
rect -62133 29902 -61517 30198
rect -61473 30172 -61177 30198
rect -61473 29928 -61447 30172
rect -61447 29928 -61203 30172
rect -61203 29928 -61177 30172
rect -61473 29902 -61177 29928
rect -61133 29902 -60517 30198
rect -60473 30172 -60177 30198
rect -60473 29928 -60447 30172
rect -60447 29928 -60203 30172
rect -60203 29928 -60177 30172
rect -60473 29902 -60177 29928
rect -60133 29902 -59517 30198
rect -59473 30172 -59177 30198
rect -59473 29928 -59447 30172
rect -59447 29928 -59203 30172
rect -59203 29928 -59177 30172
rect -59473 29902 -59177 29928
rect -59133 29902 -58837 30198
rect -74473 29242 -74177 29858
rect -73473 29242 -73177 29858
rect -72473 29242 -72177 29858
rect -71473 29242 -71177 29858
rect -70473 29242 -70177 29858
rect -69473 29242 -69177 29858
rect -68473 29242 -68177 29858
rect -67473 29242 -67177 29858
rect -66473 29242 -66177 29858
rect -65473 29242 -65177 29858
rect -64473 29242 -64177 29858
rect -63473 29242 -63177 29858
rect -62473 29242 -62177 29858
rect -61473 29242 -61177 29858
rect -60473 29242 -60177 29858
rect -59473 29242 -59177 29858
rect -74813 28902 -74517 29198
rect -74473 29172 -74177 29198
rect -74473 28928 -74447 29172
rect -74447 28928 -74203 29172
rect -74203 28928 -74177 29172
rect -74473 28902 -74177 28928
rect -74133 28902 -73517 29198
rect -73473 29172 -73177 29198
rect -73473 28928 -73447 29172
rect -73447 28928 -73203 29172
rect -73203 28928 -73177 29172
rect -73473 28902 -73177 28928
rect -73133 28902 -72517 29198
rect -72473 29172 -72177 29198
rect -72473 28928 -72447 29172
rect -72447 28928 -72203 29172
rect -72203 28928 -72177 29172
rect -72473 28902 -72177 28928
rect -72133 28902 -71517 29198
rect -71473 29172 -71177 29198
rect -71473 28928 -71447 29172
rect -71447 28928 -71203 29172
rect -71203 28928 -71177 29172
rect -71473 28902 -71177 28928
rect -71133 28902 -70517 29198
rect -70473 29172 -70177 29198
rect -70473 28928 -70447 29172
rect -70447 28928 -70203 29172
rect -70203 28928 -70177 29172
rect -70473 28902 -70177 28928
rect -70133 28902 -69517 29198
rect -69473 29172 -69177 29198
rect -69473 28928 -69447 29172
rect -69447 28928 -69203 29172
rect -69203 28928 -69177 29172
rect -69473 28902 -69177 28928
rect -69133 28902 -68517 29198
rect -68473 29172 -68177 29198
rect -68473 28928 -68447 29172
rect -68447 28928 -68203 29172
rect -68203 28928 -68177 29172
rect -68473 28902 -68177 28928
rect -68133 28902 -67517 29198
rect -67473 29172 -67177 29198
rect -67473 28928 -67447 29172
rect -67447 28928 -67203 29172
rect -67203 28928 -67177 29172
rect -67473 28902 -67177 28928
rect -67133 28902 -66517 29198
rect -66473 29172 -66177 29198
rect -66473 28928 -66447 29172
rect -66447 28928 -66203 29172
rect -66203 28928 -66177 29172
rect -66473 28902 -66177 28928
rect -66133 28902 -65517 29198
rect -65473 29172 -65177 29198
rect -65473 28928 -65447 29172
rect -65447 28928 -65203 29172
rect -65203 28928 -65177 29172
rect -65473 28902 -65177 28928
rect -65133 28902 -64517 29198
rect -64473 29172 -64177 29198
rect -64473 28928 -64447 29172
rect -64447 28928 -64203 29172
rect -64203 28928 -64177 29172
rect -64473 28902 -64177 28928
rect -64133 28902 -63517 29198
rect -63473 29172 -63177 29198
rect -63473 28928 -63447 29172
rect -63447 28928 -63203 29172
rect -63203 28928 -63177 29172
rect -63473 28902 -63177 28928
rect -63133 28902 -62517 29198
rect -62473 29172 -62177 29198
rect -62473 28928 -62447 29172
rect -62447 28928 -62203 29172
rect -62203 28928 -62177 29172
rect -62473 28902 -62177 28928
rect -62133 28902 -61517 29198
rect -61473 29172 -61177 29198
rect -61473 28928 -61447 29172
rect -61447 28928 -61203 29172
rect -61203 28928 -61177 29172
rect -61473 28902 -61177 28928
rect -61133 28902 -60517 29198
rect -60473 29172 -60177 29198
rect -60473 28928 -60447 29172
rect -60447 28928 -60203 29172
rect -60203 28928 -60177 29172
rect -60473 28902 -60177 28928
rect -60133 28902 -59517 29198
rect -59473 29172 -59177 29198
rect -59473 28928 -59447 29172
rect -59447 28928 -59203 29172
rect -59203 28928 -59177 29172
rect -59473 28902 -59177 28928
rect -59133 28902 -58837 29198
rect -74473 28562 -74177 28858
rect -73473 28562 -73177 28858
rect -72473 28562 -72177 28858
rect -71473 28562 -71177 28858
rect -70473 28562 -70177 28858
rect -69473 28562 -69177 28858
rect -68473 28562 -68177 28858
rect -67473 28562 -67177 28858
rect -66473 28562 -66177 28858
rect -65473 28562 -65177 28858
rect -64473 28562 -64177 28858
rect -63473 28562 -63177 28858
rect -62473 28562 -62177 28858
rect -61473 28562 -61177 28858
rect -60473 28562 -60177 28858
rect -59473 28562 -59177 28858
rect -72778 16047 -72776 25943
rect -72776 16047 -60884 25943
rect -60884 16047 -60882 25943
rect 10006 32242 10302 32858
rect 11006 32242 11302 32858
rect 12006 32242 12302 32858
rect 13006 32242 13302 32858
rect 14006 32242 14302 32858
rect 15006 32242 15302 32858
rect 16006 32242 16302 32858
rect 17006 32242 17302 32858
rect 18006 32242 18302 32858
rect 19006 32242 19302 32858
rect 20006 32242 20302 32858
rect 21006 32242 21302 32858
rect 22006 32242 22302 32858
rect 23006 32242 23302 32858
rect 24006 32242 24302 32858
rect 25006 32242 25302 32858
rect 26006 32242 26302 32858
rect 27006 32242 27302 32858
rect 28006 32242 28302 32858
rect 29006 32242 29302 32858
rect 30006 32242 30302 32858
rect 31006 32242 31302 32858
rect 32006 32242 32302 32858
rect 33006 32242 33302 32858
rect 34006 32242 34302 32858
rect 9666 31902 9962 32198
rect 10006 32172 10302 32198
rect 10006 31928 10032 32172
rect 10032 31928 10276 32172
rect 10276 31928 10302 32172
rect 10006 31902 10302 31928
rect 10346 31902 10962 32198
rect 11006 32172 11302 32198
rect 11006 31928 11032 32172
rect 11032 31928 11276 32172
rect 11276 31928 11302 32172
rect 11006 31902 11302 31928
rect 11346 31902 11962 32198
rect 12006 32172 12302 32198
rect 12006 31928 12032 32172
rect 12032 31928 12276 32172
rect 12276 31928 12302 32172
rect 12006 31902 12302 31928
rect 12346 31902 12962 32198
rect 13006 32172 13302 32198
rect 13006 31928 13032 32172
rect 13032 31928 13276 32172
rect 13276 31928 13302 32172
rect 13006 31902 13302 31928
rect 13346 31902 13962 32198
rect 14006 32172 14302 32198
rect 14006 31928 14032 32172
rect 14032 31928 14276 32172
rect 14276 31928 14302 32172
rect 14006 31902 14302 31928
rect 14346 31902 14962 32198
rect 15006 32172 15302 32198
rect 15006 31928 15032 32172
rect 15032 31928 15276 32172
rect 15276 31928 15302 32172
rect 15006 31902 15302 31928
rect 15346 31902 15962 32198
rect 16006 32172 16302 32198
rect 16006 31928 16032 32172
rect 16032 31928 16276 32172
rect 16276 31928 16302 32172
rect 16006 31902 16302 31928
rect 16346 31902 16962 32198
rect 17006 32172 17302 32198
rect 17006 31928 17032 32172
rect 17032 31928 17276 32172
rect 17276 31928 17302 32172
rect 17006 31902 17302 31928
rect 17346 31902 17962 32198
rect 18006 32172 18302 32198
rect 18006 31928 18032 32172
rect 18032 31928 18276 32172
rect 18276 31928 18302 32172
rect 18006 31902 18302 31928
rect 18346 31902 18962 32198
rect 19006 32172 19302 32198
rect 19006 31928 19032 32172
rect 19032 31928 19276 32172
rect 19276 31928 19302 32172
rect 19006 31902 19302 31928
rect 19346 31902 19962 32198
rect 20006 32172 20302 32198
rect 20006 31928 20032 32172
rect 20032 31928 20276 32172
rect 20276 31928 20302 32172
rect 20006 31902 20302 31928
rect 20346 31902 20962 32198
rect 21006 32172 21302 32198
rect 21006 31928 21032 32172
rect 21032 31928 21276 32172
rect 21276 31928 21302 32172
rect 21006 31902 21302 31928
rect 21346 31902 21962 32198
rect 22006 32172 22302 32198
rect 22006 31928 22032 32172
rect 22032 31928 22276 32172
rect 22276 31928 22302 32172
rect 22006 31902 22302 31928
rect 22346 31902 22962 32198
rect 23006 32172 23302 32198
rect 23006 31928 23032 32172
rect 23032 31928 23276 32172
rect 23276 31928 23302 32172
rect 23006 31902 23302 31928
rect 23346 31902 23962 32198
rect 24006 32172 24302 32198
rect 24006 31928 24032 32172
rect 24032 31928 24276 32172
rect 24276 31928 24302 32172
rect 24006 31902 24302 31928
rect 24346 31902 24962 32198
rect 25006 32172 25302 32198
rect 25006 31928 25032 32172
rect 25032 31928 25276 32172
rect 25276 31928 25302 32172
rect 25006 31902 25302 31928
rect 25346 31902 25962 32198
rect 26006 32172 26302 32198
rect 26006 31928 26032 32172
rect 26032 31928 26276 32172
rect 26276 31928 26302 32172
rect 26006 31902 26302 31928
rect 26346 31902 26962 32198
rect 27006 32172 27302 32198
rect 27006 31928 27032 32172
rect 27032 31928 27276 32172
rect 27276 31928 27302 32172
rect 27006 31902 27302 31928
rect 27346 31902 27962 32198
rect 28006 32172 28302 32198
rect 28006 31928 28032 32172
rect 28032 31928 28276 32172
rect 28276 31928 28302 32172
rect 28006 31902 28302 31928
rect 28346 31902 28962 32198
rect 29006 32172 29302 32198
rect 29006 31928 29032 32172
rect 29032 31928 29276 32172
rect 29276 31928 29302 32172
rect 29006 31902 29302 31928
rect 29346 31902 29962 32198
rect 30006 32172 30302 32198
rect 30006 31928 30032 32172
rect 30032 31928 30276 32172
rect 30276 31928 30302 32172
rect 30006 31902 30302 31928
rect 30346 31902 30962 32198
rect 31006 32172 31302 32198
rect 31006 31928 31032 32172
rect 31032 31928 31276 32172
rect 31276 31928 31302 32172
rect 31006 31902 31302 31928
rect 31346 31902 31962 32198
rect 32006 32172 32302 32198
rect 32006 31928 32032 32172
rect 32032 31928 32276 32172
rect 32276 31928 32302 32172
rect 32006 31902 32302 31928
rect 32346 31902 32962 32198
rect 33006 32172 33302 32198
rect 33006 31928 33032 32172
rect 33032 31928 33276 32172
rect 33276 31928 33302 32172
rect 33006 31902 33302 31928
rect 33346 31902 33962 32198
rect 34006 32172 34302 32198
rect 34006 31928 34032 32172
rect 34032 31928 34276 32172
rect 34276 31928 34302 32172
rect 34006 31902 34302 31928
rect 34346 31902 34642 32198
rect 10006 31242 10302 31858
rect 11006 31242 11302 31858
rect 12006 31242 12302 31858
rect 13006 31242 13302 31858
rect 14006 31242 14302 31858
rect 15006 31242 15302 31858
rect 16006 31242 16302 31858
rect 17006 31242 17302 31858
rect 18006 31242 18302 31858
rect 19006 31242 19302 31858
rect 20006 31242 20302 31858
rect 21006 31242 21302 31858
rect 22006 31242 22302 31858
rect 23006 31242 23302 31858
rect 24006 31242 24302 31858
rect 25006 31242 25302 31858
rect 26006 31242 26302 31858
rect 27006 31242 27302 31858
rect 28006 31242 28302 31858
rect 29006 31242 29302 31858
rect 30006 31242 30302 31858
rect 31006 31242 31302 31858
rect 32006 31242 32302 31858
rect 33006 31242 33302 31858
rect 34006 31242 34302 31858
rect 9666 30902 9962 31198
rect 10006 31172 10302 31198
rect 10006 30928 10032 31172
rect 10032 30928 10276 31172
rect 10276 30928 10302 31172
rect 10006 30902 10302 30928
rect 10346 30902 10962 31198
rect 11006 31172 11302 31198
rect 11006 30928 11032 31172
rect 11032 30928 11276 31172
rect 11276 30928 11302 31172
rect 11006 30902 11302 30928
rect 11346 30902 11962 31198
rect 12006 31172 12302 31198
rect 12006 30928 12032 31172
rect 12032 30928 12276 31172
rect 12276 30928 12302 31172
rect 12006 30902 12302 30928
rect 12346 30902 12962 31198
rect 13006 31172 13302 31198
rect 13006 30928 13032 31172
rect 13032 30928 13276 31172
rect 13276 30928 13302 31172
rect 13006 30902 13302 30928
rect 13346 30902 13962 31198
rect 14006 31172 14302 31198
rect 14006 30928 14032 31172
rect 14032 30928 14276 31172
rect 14276 30928 14302 31172
rect 14006 30902 14302 30928
rect 14346 30902 14962 31198
rect 15006 31172 15302 31198
rect 15006 30928 15032 31172
rect 15032 30928 15276 31172
rect 15276 30928 15302 31172
rect 15006 30902 15302 30928
rect 15346 30902 15962 31198
rect 16006 31172 16302 31198
rect 16006 30928 16032 31172
rect 16032 30928 16276 31172
rect 16276 30928 16302 31172
rect 16006 30902 16302 30928
rect 16346 30902 16962 31198
rect 17006 31172 17302 31198
rect 17006 30928 17032 31172
rect 17032 30928 17276 31172
rect 17276 30928 17302 31172
rect 17006 30902 17302 30928
rect 17346 30902 17962 31198
rect 18006 31172 18302 31198
rect 18006 30928 18032 31172
rect 18032 30928 18276 31172
rect 18276 30928 18302 31172
rect 18006 30902 18302 30928
rect 18346 30902 18962 31198
rect 19006 31172 19302 31198
rect 19006 30928 19032 31172
rect 19032 30928 19276 31172
rect 19276 30928 19302 31172
rect 19006 30902 19302 30928
rect 19346 30902 19962 31198
rect 20006 31172 20302 31198
rect 20006 30928 20032 31172
rect 20032 30928 20276 31172
rect 20276 30928 20302 31172
rect 20006 30902 20302 30928
rect 20346 30902 20962 31198
rect 21006 31172 21302 31198
rect 21006 30928 21032 31172
rect 21032 30928 21276 31172
rect 21276 30928 21302 31172
rect 21006 30902 21302 30928
rect 21346 30902 21962 31198
rect 22006 31172 22302 31198
rect 22006 30928 22032 31172
rect 22032 30928 22276 31172
rect 22276 30928 22302 31172
rect 22006 30902 22302 30928
rect 22346 30902 22962 31198
rect 23006 31172 23302 31198
rect 23006 30928 23032 31172
rect 23032 30928 23276 31172
rect 23276 30928 23302 31172
rect 23006 30902 23302 30928
rect 23346 30902 23962 31198
rect 24006 31172 24302 31198
rect 24006 30928 24032 31172
rect 24032 30928 24276 31172
rect 24276 30928 24302 31172
rect 24006 30902 24302 30928
rect 24346 30902 24962 31198
rect 25006 31172 25302 31198
rect 25006 30928 25032 31172
rect 25032 30928 25276 31172
rect 25276 30928 25302 31172
rect 25006 30902 25302 30928
rect 25346 30902 25962 31198
rect 26006 31172 26302 31198
rect 26006 30928 26032 31172
rect 26032 30928 26276 31172
rect 26276 30928 26302 31172
rect 26006 30902 26302 30928
rect 26346 30902 26962 31198
rect 27006 31172 27302 31198
rect 27006 30928 27032 31172
rect 27032 30928 27276 31172
rect 27276 30928 27302 31172
rect 27006 30902 27302 30928
rect 27346 30902 27962 31198
rect 28006 31172 28302 31198
rect 28006 30928 28032 31172
rect 28032 30928 28276 31172
rect 28276 30928 28302 31172
rect 28006 30902 28302 30928
rect 28346 30902 28962 31198
rect 29006 31172 29302 31198
rect 29006 30928 29032 31172
rect 29032 30928 29276 31172
rect 29276 30928 29302 31172
rect 29006 30902 29302 30928
rect 29346 30902 29962 31198
rect 30006 31172 30302 31198
rect 30006 30928 30032 31172
rect 30032 30928 30276 31172
rect 30276 30928 30302 31172
rect 30006 30902 30302 30928
rect 30346 30902 30962 31198
rect 31006 31172 31302 31198
rect 31006 30928 31032 31172
rect 31032 30928 31276 31172
rect 31276 30928 31302 31172
rect 31006 30902 31302 30928
rect 31346 30902 31962 31198
rect 32006 31172 32302 31198
rect 32006 30928 32032 31172
rect 32032 30928 32276 31172
rect 32276 30928 32302 31172
rect 32006 30902 32302 30928
rect 32346 30902 32962 31198
rect 33006 31172 33302 31198
rect 33006 30928 33032 31172
rect 33032 30928 33276 31172
rect 33276 30928 33302 31172
rect 33006 30902 33302 30928
rect 33346 30902 33962 31198
rect 34006 31172 34302 31198
rect 34006 30928 34032 31172
rect 34032 30928 34276 31172
rect 34276 30928 34302 31172
rect 34006 30902 34302 30928
rect 34346 30902 34642 31198
rect 10006 30242 10302 30858
rect 11006 30242 11302 30858
rect 12006 30242 12302 30858
rect 13006 30242 13302 30858
rect 14006 30242 14302 30858
rect 15006 30242 15302 30858
rect 16006 30242 16302 30858
rect 17006 30242 17302 30858
rect 18006 30242 18302 30858
rect 19006 30242 19302 30858
rect 20006 30242 20302 30858
rect 21006 30242 21302 30858
rect 22006 30242 22302 30858
rect 23006 30242 23302 30858
rect 24006 30242 24302 30858
rect 25006 30242 25302 30858
rect 26006 30242 26302 30858
rect 27006 30242 27302 30858
rect 28006 30242 28302 30858
rect 29006 30242 29302 30858
rect 30006 30242 30302 30858
rect 31006 30242 31302 30858
rect 32006 30242 32302 30858
rect 33006 30242 33302 30858
rect 34006 30242 34302 30858
rect 9666 29902 9962 30198
rect 10006 30172 10302 30198
rect 10006 29928 10032 30172
rect 10032 29928 10276 30172
rect 10276 29928 10302 30172
rect 10006 29902 10302 29928
rect 10346 29902 10962 30198
rect 11006 30172 11302 30198
rect 11006 29928 11032 30172
rect 11032 29928 11276 30172
rect 11276 29928 11302 30172
rect 11006 29902 11302 29928
rect 11346 29902 11962 30198
rect 12006 30172 12302 30198
rect 12006 29928 12032 30172
rect 12032 29928 12276 30172
rect 12276 29928 12302 30172
rect 12006 29902 12302 29928
rect 12346 29902 12962 30198
rect 13006 30172 13302 30198
rect 13006 29928 13032 30172
rect 13032 29928 13276 30172
rect 13276 29928 13302 30172
rect 13006 29902 13302 29928
rect 13346 29902 13962 30198
rect 14006 30172 14302 30198
rect 14006 29928 14032 30172
rect 14032 29928 14276 30172
rect 14276 29928 14302 30172
rect 14006 29902 14302 29928
rect 14346 29902 14962 30198
rect 15006 30172 15302 30198
rect 15006 29928 15032 30172
rect 15032 29928 15276 30172
rect 15276 29928 15302 30172
rect 15006 29902 15302 29928
rect 15346 29902 15962 30198
rect 16006 30172 16302 30198
rect 16006 29928 16032 30172
rect 16032 29928 16276 30172
rect 16276 29928 16302 30172
rect 16006 29902 16302 29928
rect 16346 29902 16962 30198
rect 17006 30172 17302 30198
rect 17006 29928 17032 30172
rect 17032 29928 17276 30172
rect 17276 29928 17302 30172
rect 17006 29902 17302 29928
rect 17346 29902 17962 30198
rect 18006 30172 18302 30198
rect 18006 29928 18032 30172
rect 18032 29928 18276 30172
rect 18276 29928 18302 30172
rect 18006 29902 18302 29928
rect 18346 29902 18962 30198
rect 19006 30172 19302 30198
rect 19006 29928 19032 30172
rect 19032 29928 19276 30172
rect 19276 29928 19302 30172
rect 19006 29902 19302 29928
rect 19346 29902 19962 30198
rect 20006 30172 20302 30198
rect 20006 29928 20032 30172
rect 20032 29928 20276 30172
rect 20276 29928 20302 30172
rect 20006 29902 20302 29928
rect 20346 29902 20962 30198
rect 21006 30172 21302 30198
rect 21006 29928 21032 30172
rect 21032 29928 21276 30172
rect 21276 29928 21302 30172
rect 21006 29902 21302 29928
rect 21346 29902 21962 30198
rect 22006 30172 22302 30198
rect 22006 29928 22032 30172
rect 22032 29928 22276 30172
rect 22276 29928 22302 30172
rect 22006 29902 22302 29928
rect 22346 29902 22962 30198
rect 23006 30172 23302 30198
rect 23006 29928 23032 30172
rect 23032 29928 23276 30172
rect 23276 29928 23302 30172
rect 23006 29902 23302 29928
rect 23346 29902 23962 30198
rect 24006 30172 24302 30198
rect 24006 29928 24032 30172
rect 24032 29928 24276 30172
rect 24276 29928 24302 30172
rect 24006 29902 24302 29928
rect 24346 29902 24962 30198
rect 25006 30172 25302 30198
rect 25006 29928 25032 30172
rect 25032 29928 25276 30172
rect 25276 29928 25302 30172
rect 25006 29902 25302 29928
rect 25346 29902 25962 30198
rect 26006 30172 26302 30198
rect 26006 29928 26032 30172
rect 26032 29928 26276 30172
rect 26276 29928 26302 30172
rect 26006 29902 26302 29928
rect 26346 29902 26962 30198
rect 27006 30172 27302 30198
rect 27006 29928 27032 30172
rect 27032 29928 27276 30172
rect 27276 29928 27302 30172
rect 27006 29902 27302 29928
rect 27346 29902 27962 30198
rect 28006 30172 28302 30198
rect 28006 29928 28032 30172
rect 28032 29928 28276 30172
rect 28276 29928 28302 30172
rect 28006 29902 28302 29928
rect 28346 29902 28962 30198
rect 29006 30172 29302 30198
rect 29006 29928 29032 30172
rect 29032 29928 29276 30172
rect 29276 29928 29302 30172
rect 29006 29902 29302 29928
rect 29346 29902 29962 30198
rect 30006 30172 30302 30198
rect 30006 29928 30032 30172
rect 30032 29928 30276 30172
rect 30276 29928 30302 30172
rect 30006 29902 30302 29928
rect 30346 29902 30962 30198
rect 31006 30172 31302 30198
rect 31006 29928 31032 30172
rect 31032 29928 31276 30172
rect 31276 29928 31302 30172
rect 31006 29902 31302 29928
rect 31346 29902 31962 30198
rect 32006 30172 32302 30198
rect 32006 29928 32032 30172
rect 32032 29928 32276 30172
rect 32276 29928 32302 30172
rect 32006 29902 32302 29928
rect 32346 29902 32962 30198
rect 33006 30172 33302 30198
rect 33006 29928 33032 30172
rect 33032 29928 33276 30172
rect 33276 29928 33302 30172
rect 33006 29902 33302 29928
rect 33346 29902 33962 30198
rect 34006 30172 34302 30198
rect 34006 29928 34032 30172
rect 34032 29928 34276 30172
rect 34276 29928 34302 30172
rect 34006 29902 34302 29928
rect 34346 29902 34642 30198
rect 10006 29242 10302 29858
rect 11006 29242 11302 29858
rect 12006 29242 12302 29858
rect 13006 29242 13302 29858
rect 14006 29242 14302 29858
rect 15006 29242 15302 29858
rect 16006 29242 16302 29858
rect 17006 29242 17302 29858
rect 18006 29242 18302 29858
rect 19006 29242 19302 29858
rect 20006 29242 20302 29858
rect 21006 29242 21302 29858
rect 22006 29242 22302 29858
rect 23006 29242 23302 29858
rect 24006 29242 24302 29858
rect 25006 29242 25302 29858
rect 26006 29242 26302 29858
rect 27006 29242 27302 29858
rect 28006 29242 28302 29858
rect 29006 29242 29302 29858
rect 30006 29242 30302 29858
rect 31006 29242 31302 29858
rect 32006 29242 32302 29858
rect 33006 29242 33302 29858
rect 34006 29242 34302 29858
rect 9666 28902 9962 29198
rect 10006 29172 10302 29198
rect 10006 28928 10032 29172
rect 10032 28928 10276 29172
rect 10276 28928 10302 29172
rect 10006 28902 10302 28928
rect 10346 28902 10962 29198
rect 11006 29172 11302 29198
rect 11006 28928 11032 29172
rect 11032 28928 11276 29172
rect 11276 28928 11302 29172
rect 11006 28902 11302 28928
rect 11346 28902 11962 29198
rect 12006 29172 12302 29198
rect 12006 28928 12032 29172
rect 12032 28928 12276 29172
rect 12276 28928 12302 29172
rect 12006 28902 12302 28928
rect 12346 28902 12962 29198
rect 13006 29172 13302 29198
rect 13006 28928 13032 29172
rect 13032 28928 13276 29172
rect 13276 28928 13302 29172
rect 13006 28902 13302 28928
rect 13346 28902 13962 29198
rect 14006 29172 14302 29198
rect 14006 28928 14032 29172
rect 14032 28928 14276 29172
rect 14276 28928 14302 29172
rect 14006 28902 14302 28928
rect 14346 28902 14962 29198
rect 15006 29172 15302 29198
rect 15006 28928 15032 29172
rect 15032 28928 15276 29172
rect 15276 28928 15302 29172
rect 15006 28902 15302 28928
rect 15346 28902 15962 29198
rect 16006 29172 16302 29198
rect 16006 28928 16032 29172
rect 16032 28928 16276 29172
rect 16276 28928 16302 29172
rect 16006 28902 16302 28928
rect 16346 28902 16962 29198
rect 17006 29172 17302 29198
rect 17006 28928 17032 29172
rect 17032 28928 17276 29172
rect 17276 28928 17302 29172
rect 17006 28902 17302 28928
rect 17346 28902 17962 29198
rect 18006 29172 18302 29198
rect 18006 28928 18032 29172
rect 18032 28928 18276 29172
rect 18276 28928 18302 29172
rect 18006 28902 18302 28928
rect 18346 28902 18962 29198
rect 19006 29172 19302 29198
rect 19006 28928 19032 29172
rect 19032 28928 19276 29172
rect 19276 28928 19302 29172
rect 19006 28902 19302 28928
rect 19346 28902 19962 29198
rect 20006 29172 20302 29198
rect 20006 28928 20032 29172
rect 20032 28928 20276 29172
rect 20276 28928 20302 29172
rect 20006 28902 20302 28928
rect 20346 28902 20962 29198
rect 21006 29172 21302 29198
rect 21006 28928 21032 29172
rect 21032 28928 21276 29172
rect 21276 28928 21302 29172
rect 21006 28902 21302 28928
rect 21346 28902 21962 29198
rect 22006 29172 22302 29198
rect 22006 28928 22032 29172
rect 22032 28928 22276 29172
rect 22276 28928 22302 29172
rect 22006 28902 22302 28928
rect 22346 28902 22962 29198
rect 23006 29172 23302 29198
rect 23006 28928 23032 29172
rect 23032 28928 23276 29172
rect 23276 28928 23302 29172
rect 23006 28902 23302 28928
rect 23346 28902 23962 29198
rect 24006 29172 24302 29198
rect 24006 28928 24032 29172
rect 24032 28928 24276 29172
rect 24276 28928 24302 29172
rect 24006 28902 24302 28928
rect 24346 28902 24962 29198
rect 25006 29172 25302 29198
rect 25006 28928 25032 29172
rect 25032 28928 25276 29172
rect 25276 28928 25302 29172
rect 25006 28902 25302 28928
rect 25346 28902 25962 29198
rect 26006 29172 26302 29198
rect 26006 28928 26032 29172
rect 26032 28928 26276 29172
rect 26276 28928 26302 29172
rect 26006 28902 26302 28928
rect 26346 28902 26962 29198
rect 27006 29172 27302 29198
rect 27006 28928 27032 29172
rect 27032 28928 27276 29172
rect 27276 28928 27302 29172
rect 27006 28902 27302 28928
rect 27346 28902 27962 29198
rect 28006 29172 28302 29198
rect 28006 28928 28032 29172
rect 28032 28928 28276 29172
rect 28276 28928 28302 29172
rect 28006 28902 28302 28928
rect 28346 28902 28962 29198
rect 29006 29172 29302 29198
rect 29006 28928 29032 29172
rect 29032 28928 29276 29172
rect 29276 28928 29302 29172
rect 29006 28902 29302 28928
rect 29346 28902 29962 29198
rect 30006 29172 30302 29198
rect 30006 28928 30032 29172
rect 30032 28928 30276 29172
rect 30276 28928 30302 29172
rect 30006 28902 30302 28928
rect 30346 28902 30962 29198
rect 31006 29172 31302 29198
rect 31006 28928 31032 29172
rect 31032 28928 31276 29172
rect 31276 28928 31302 29172
rect 31006 28902 31302 28928
rect 31346 28902 31962 29198
rect 32006 29172 32302 29198
rect 32006 28928 32032 29172
rect 32032 28928 32276 29172
rect 32276 28928 32302 29172
rect 32006 28902 32302 28928
rect 32346 28902 32962 29198
rect 33006 29172 33302 29198
rect 33006 28928 33032 29172
rect 33032 28928 33276 29172
rect 33276 28928 33302 29172
rect 33006 28902 33302 28928
rect 33346 28902 33962 29198
rect 34006 29172 34302 29198
rect 34006 28928 34032 29172
rect 34032 28928 34276 29172
rect 34276 28928 34302 29172
rect 34006 28902 34302 28928
rect 34346 28902 34642 29198
rect 10006 28562 10302 28858
rect 11006 28562 11302 28858
rect 12006 28562 12302 28858
rect 13006 28562 13302 28858
rect 14006 28562 14302 28858
rect 15006 28562 15302 28858
rect 16006 28562 16302 28858
rect 17006 28562 17302 28858
rect 18006 28562 18302 28858
rect 19006 28562 19302 28858
rect 20006 28562 20302 28858
rect 21006 28562 21302 28858
rect 22006 28562 22302 28858
rect 23006 28562 23302 28858
rect 24006 28562 24302 28858
rect 25006 28562 25302 28858
rect 26006 28562 26302 28858
rect 27006 28562 27302 28858
rect 28006 28562 28302 28858
rect 29006 28562 29302 28858
rect 30006 28562 30302 28858
rect 31006 28562 31302 28858
rect 32006 28562 32302 28858
rect 33006 28562 33302 28858
rect 34006 28562 34302 28858
rect 20322 16052 20324 25948
rect 20324 16052 32216 25948
rect 32216 16052 32218 25948
rect -21206 13862 -19310 15118
rect -42378 7902 -40722 13798
rect 172 7902 1828 13798
rect -42378 2298 -40722 2308
rect -42378 -2298 -40722 2298
rect -42378 -2308 -40722 -2298
rect 172 2298 1828 2308
rect 172 -2298 1828 2298
rect 172 -2308 1828 -2298
rect -42378 -13798 -40722 -7902
rect 172 -13798 1828 -7902
rect -72778 -25948 -72776 -16052
rect -72776 -25948 -60884 -16052
rect -60884 -25948 -60882 -16052
rect 20322 -25948 20324 -16052
rect 20324 -25948 32216 -16052
rect 32216 -25948 32218 -16052
rect -74473 -28858 -74177 -28562
rect -73473 -28858 -73177 -28562
rect -72473 -28858 -72177 -28562
rect -71473 -28858 -71177 -28562
rect -70473 -28858 -70177 -28562
rect -69473 -28858 -69177 -28562
rect -68473 -28858 -68177 -28562
rect -67473 -28858 -67177 -28562
rect -66473 -28858 -66177 -28562
rect -65473 -28858 -65177 -28562
rect -64473 -28858 -64177 -28562
rect -63473 -28858 -63177 -28562
rect -62473 -28858 -62177 -28562
rect -61473 -28858 -61177 -28562
rect -60473 -28858 -60177 -28562
rect -59473 -28858 -59177 -28562
rect -58473 -28858 -58177 -28562
rect -57473 -28858 -57177 -28562
rect -56473 -28858 -56177 -28562
rect -55473 -28858 -55177 -28562
rect -54473 -28858 -54177 -28562
rect -53473 -28858 -53177 -28562
rect -52473 -28858 -52177 -28562
rect -51473 -28858 -51177 -28562
rect -50473 -28858 -50177 -28562
rect -49473 -28858 -49177 -28562
rect 8627 -28858 8923 -28562
rect 9627 -28858 9923 -28562
rect 10627 -28858 10923 -28562
rect 11627 -28858 11923 -28562
rect 12627 -28858 12923 -28562
rect 13627 -28858 13923 -28562
rect 14627 -28858 14923 -28562
rect 15627 -28858 15923 -28562
rect 16627 -28858 16923 -28562
rect 17627 -28858 17923 -28562
rect 18627 -28858 18923 -28562
rect 19627 -28858 19923 -28562
rect 20627 -28858 20923 -28562
rect 21627 -28858 21923 -28562
rect 22627 -28858 22923 -28562
rect 23627 -28858 23923 -28562
rect 24627 -28858 24923 -28562
rect 25627 -28858 25923 -28562
rect 26627 -28858 26923 -28562
rect 27627 -28858 27923 -28562
rect 28627 -28858 28923 -28562
rect 29627 -28858 29923 -28562
rect 30627 -28858 30923 -28562
rect 31627 -28858 31923 -28562
rect 32627 -28858 32923 -28562
rect 33627 -28858 33923 -28562
rect -74813 -29198 -74517 -28902
rect -74473 -28928 -74177 -28902
rect -74473 -29172 -74447 -28928
rect -74447 -29172 -74203 -28928
rect -74203 -29172 -74177 -28928
rect -74473 -29198 -74177 -29172
rect -74133 -29198 -73517 -28902
rect -73473 -28928 -73177 -28902
rect -73473 -29172 -73447 -28928
rect -73447 -29172 -73203 -28928
rect -73203 -29172 -73177 -28928
rect -73473 -29198 -73177 -29172
rect -73133 -29198 -72517 -28902
rect -72473 -28928 -72177 -28902
rect -72473 -29172 -72447 -28928
rect -72447 -29172 -72203 -28928
rect -72203 -29172 -72177 -28928
rect -72473 -29198 -72177 -29172
rect -72133 -29198 -71517 -28902
rect -71473 -28928 -71177 -28902
rect -71473 -29172 -71447 -28928
rect -71447 -29172 -71203 -28928
rect -71203 -29172 -71177 -28928
rect -71473 -29198 -71177 -29172
rect -71133 -29198 -70517 -28902
rect -70473 -28928 -70177 -28902
rect -70473 -29172 -70447 -28928
rect -70447 -29172 -70203 -28928
rect -70203 -29172 -70177 -28928
rect -70473 -29198 -70177 -29172
rect -70133 -29198 -69517 -28902
rect -69473 -28928 -69177 -28902
rect -69473 -29172 -69447 -28928
rect -69447 -29172 -69203 -28928
rect -69203 -29172 -69177 -28928
rect -69473 -29198 -69177 -29172
rect -69133 -29198 -68517 -28902
rect -68473 -28928 -68177 -28902
rect -68473 -29172 -68447 -28928
rect -68447 -29172 -68203 -28928
rect -68203 -29172 -68177 -28928
rect -68473 -29198 -68177 -29172
rect -68133 -29198 -67517 -28902
rect -67473 -28928 -67177 -28902
rect -67473 -29172 -67447 -28928
rect -67447 -29172 -67203 -28928
rect -67203 -29172 -67177 -28928
rect -67473 -29198 -67177 -29172
rect -67133 -29198 -66517 -28902
rect -66473 -28928 -66177 -28902
rect -66473 -29172 -66447 -28928
rect -66447 -29172 -66203 -28928
rect -66203 -29172 -66177 -28928
rect -66473 -29198 -66177 -29172
rect -66133 -29198 -65517 -28902
rect -65473 -28928 -65177 -28902
rect -65473 -29172 -65447 -28928
rect -65447 -29172 -65203 -28928
rect -65203 -29172 -65177 -28928
rect -65473 -29198 -65177 -29172
rect -65133 -29198 -64517 -28902
rect -64473 -28928 -64177 -28902
rect -64473 -29172 -64447 -28928
rect -64447 -29172 -64203 -28928
rect -64203 -29172 -64177 -28928
rect -64473 -29198 -64177 -29172
rect -64133 -29198 -63517 -28902
rect -63473 -28928 -63177 -28902
rect -63473 -29172 -63447 -28928
rect -63447 -29172 -63203 -28928
rect -63203 -29172 -63177 -28928
rect -63473 -29198 -63177 -29172
rect -63133 -29198 -62517 -28902
rect -62473 -28928 -62177 -28902
rect -62473 -29172 -62447 -28928
rect -62447 -29172 -62203 -28928
rect -62203 -29172 -62177 -28928
rect -62473 -29198 -62177 -29172
rect -62133 -29198 -61517 -28902
rect -61473 -28928 -61177 -28902
rect -61473 -29172 -61447 -28928
rect -61447 -29172 -61203 -28928
rect -61203 -29172 -61177 -28928
rect -61473 -29198 -61177 -29172
rect -61133 -29198 -60517 -28902
rect -60473 -28928 -60177 -28902
rect -60473 -29172 -60447 -28928
rect -60447 -29172 -60203 -28928
rect -60203 -29172 -60177 -28928
rect -60473 -29198 -60177 -29172
rect -60133 -29198 -59517 -28902
rect -59473 -28928 -59177 -28902
rect -59473 -29172 -59447 -28928
rect -59447 -29172 -59203 -28928
rect -59203 -29172 -59177 -28928
rect -59473 -29198 -59177 -29172
rect -59133 -29198 -58517 -28902
rect -58473 -28928 -58177 -28902
rect -58473 -29172 -58447 -28928
rect -58447 -29172 -58203 -28928
rect -58203 -29172 -58177 -28928
rect -58473 -29198 -58177 -29172
rect -58133 -29198 -57517 -28902
rect -57473 -28928 -57177 -28902
rect -57473 -29172 -57447 -28928
rect -57447 -29172 -57203 -28928
rect -57203 -29172 -57177 -28928
rect -57473 -29198 -57177 -29172
rect -57133 -29198 -56517 -28902
rect -56473 -28928 -56177 -28902
rect -56473 -29172 -56447 -28928
rect -56447 -29172 -56203 -28928
rect -56203 -29172 -56177 -28928
rect -56473 -29198 -56177 -29172
rect -56133 -29198 -55517 -28902
rect -55473 -28928 -55177 -28902
rect -55473 -29172 -55447 -28928
rect -55447 -29172 -55203 -28928
rect -55203 -29172 -55177 -28928
rect -55473 -29198 -55177 -29172
rect -55133 -29198 -54517 -28902
rect -54473 -28928 -54177 -28902
rect -54473 -29172 -54447 -28928
rect -54447 -29172 -54203 -28928
rect -54203 -29172 -54177 -28928
rect -54473 -29198 -54177 -29172
rect -54133 -29198 -53517 -28902
rect -53473 -28928 -53177 -28902
rect -53473 -29172 -53447 -28928
rect -53447 -29172 -53203 -28928
rect -53203 -29172 -53177 -28928
rect -53473 -29198 -53177 -29172
rect -53133 -29198 -52517 -28902
rect -52473 -28928 -52177 -28902
rect -52473 -29172 -52447 -28928
rect -52447 -29172 -52203 -28928
rect -52203 -29172 -52177 -28928
rect -52473 -29198 -52177 -29172
rect -52133 -29198 -51517 -28902
rect -51473 -28928 -51177 -28902
rect -51473 -29172 -51447 -28928
rect -51447 -29172 -51203 -28928
rect -51203 -29172 -51177 -28928
rect -51473 -29198 -51177 -29172
rect -51133 -29198 -50517 -28902
rect -50473 -28928 -50177 -28902
rect -50473 -29172 -50447 -28928
rect -50447 -29172 -50203 -28928
rect -50203 -29172 -50177 -28928
rect -50473 -29198 -50177 -29172
rect -50133 -29198 -49517 -28902
rect -49473 -28928 -49177 -28902
rect -49473 -29172 -49447 -28928
rect -49447 -29172 -49203 -28928
rect -49203 -29172 -49177 -28928
rect -49473 -29198 -49177 -29172
rect -49133 -29198 -48837 -28902
rect 8287 -29198 8583 -28902
rect 8627 -28928 8923 -28902
rect 8627 -29172 8653 -28928
rect 8653 -29172 8897 -28928
rect 8897 -29172 8923 -28928
rect 8627 -29198 8923 -29172
rect 8967 -29198 9583 -28902
rect 9627 -28928 9923 -28902
rect 9627 -29172 9653 -28928
rect 9653 -29172 9897 -28928
rect 9897 -29172 9923 -28928
rect 9627 -29198 9923 -29172
rect 9967 -29198 10583 -28902
rect 10627 -28928 10923 -28902
rect 10627 -29172 10653 -28928
rect 10653 -29172 10897 -28928
rect 10897 -29172 10923 -28928
rect 10627 -29198 10923 -29172
rect 10967 -29198 11583 -28902
rect 11627 -28928 11923 -28902
rect 11627 -29172 11653 -28928
rect 11653 -29172 11897 -28928
rect 11897 -29172 11923 -28928
rect 11627 -29198 11923 -29172
rect 11967 -29198 12583 -28902
rect 12627 -28928 12923 -28902
rect 12627 -29172 12653 -28928
rect 12653 -29172 12897 -28928
rect 12897 -29172 12923 -28928
rect 12627 -29198 12923 -29172
rect 12967 -29198 13583 -28902
rect 13627 -28928 13923 -28902
rect 13627 -29172 13653 -28928
rect 13653 -29172 13897 -28928
rect 13897 -29172 13923 -28928
rect 13627 -29198 13923 -29172
rect 13967 -29198 14583 -28902
rect 14627 -28928 14923 -28902
rect 14627 -29172 14653 -28928
rect 14653 -29172 14897 -28928
rect 14897 -29172 14923 -28928
rect 14627 -29198 14923 -29172
rect 14967 -29198 15583 -28902
rect 15627 -28928 15923 -28902
rect 15627 -29172 15653 -28928
rect 15653 -29172 15897 -28928
rect 15897 -29172 15923 -28928
rect 15627 -29198 15923 -29172
rect 15967 -29198 16583 -28902
rect 16627 -28928 16923 -28902
rect 16627 -29172 16653 -28928
rect 16653 -29172 16897 -28928
rect 16897 -29172 16923 -28928
rect 16627 -29198 16923 -29172
rect 16967 -29198 17583 -28902
rect 17627 -28928 17923 -28902
rect 17627 -29172 17653 -28928
rect 17653 -29172 17897 -28928
rect 17897 -29172 17923 -28928
rect 17627 -29198 17923 -29172
rect 17967 -29198 18583 -28902
rect 18627 -28928 18923 -28902
rect 18627 -29172 18653 -28928
rect 18653 -29172 18897 -28928
rect 18897 -29172 18923 -28928
rect 18627 -29198 18923 -29172
rect 18967 -29198 19583 -28902
rect 19627 -28928 19923 -28902
rect 19627 -29172 19653 -28928
rect 19653 -29172 19897 -28928
rect 19897 -29172 19923 -28928
rect 19627 -29198 19923 -29172
rect 19967 -29198 20583 -28902
rect 20627 -28928 20923 -28902
rect 20627 -29172 20653 -28928
rect 20653 -29172 20897 -28928
rect 20897 -29172 20923 -28928
rect 20627 -29198 20923 -29172
rect 20967 -29198 21583 -28902
rect 21627 -28928 21923 -28902
rect 21627 -29172 21653 -28928
rect 21653 -29172 21897 -28928
rect 21897 -29172 21923 -28928
rect 21627 -29198 21923 -29172
rect 21967 -29198 22583 -28902
rect 22627 -28928 22923 -28902
rect 22627 -29172 22653 -28928
rect 22653 -29172 22897 -28928
rect 22897 -29172 22923 -28928
rect 22627 -29198 22923 -29172
rect 22967 -29198 23583 -28902
rect 23627 -28928 23923 -28902
rect 23627 -29172 23653 -28928
rect 23653 -29172 23897 -28928
rect 23897 -29172 23923 -28928
rect 23627 -29198 23923 -29172
rect 23967 -29198 24583 -28902
rect 24627 -28928 24923 -28902
rect 24627 -29172 24653 -28928
rect 24653 -29172 24897 -28928
rect 24897 -29172 24923 -28928
rect 24627 -29198 24923 -29172
rect 24967 -29198 25583 -28902
rect 25627 -28928 25923 -28902
rect 25627 -29172 25653 -28928
rect 25653 -29172 25897 -28928
rect 25897 -29172 25923 -28928
rect 25627 -29198 25923 -29172
rect 25967 -29198 26583 -28902
rect 26627 -28928 26923 -28902
rect 26627 -29172 26653 -28928
rect 26653 -29172 26897 -28928
rect 26897 -29172 26923 -28928
rect 26627 -29198 26923 -29172
rect 26967 -29198 27583 -28902
rect 27627 -28928 27923 -28902
rect 27627 -29172 27653 -28928
rect 27653 -29172 27897 -28928
rect 27897 -29172 27923 -28928
rect 27627 -29198 27923 -29172
rect 27967 -29198 28583 -28902
rect 28627 -28928 28923 -28902
rect 28627 -29172 28653 -28928
rect 28653 -29172 28897 -28928
rect 28897 -29172 28923 -28928
rect 28627 -29198 28923 -29172
rect 28967 -29198 29583 -28902
rect 29627 -28928 29923 -28902
rect 29627 -29172 29653 -28928
rect 29653 -29172 29897 -28928
rect 29897 -29172 29923 -28928
rect 29627 -29198 29923 -29172
rect 29967 -29198 30583 -28902
rect 30627 -28928 30923 -28902
rect 30627 -29172 30653 -28928
rect 30653 -29172 30897 -28928
rect 30897 -29172 30923 -28928
rect 30627 -29198 30923 -29172
rect 30967 -29198 31583 -28902
rect 31627 -28928 31923 -28902
rect 31627 -29172 31653 -28928
rect 31653 -29172 31897 -28928
rect 31897 -29172 31923 -28928
rect 31627 -29198 31923 -29172
rect 31967 -29198 32583 -28902
rect 32627 -28928 32923 -28902
rect 32627 -29172 32653 -28928
rect 32653 -29172 32897 -28928
rect 32897 -29172 32923 -28928
rect 32627 -29198 32923 -29172
rect 32967 -29198 33583 -28902
rect 33627 -28928 33923 -28902
rect 33627 -29172 33653 -28928
rect 33653 -29172 33897 -28928
rect 33897 -29172 33923 -28928
rect 33627 -29198 33923 -29172
rect 33967 -29198 34263 -28902
rect -74473 -29858 -74177 -29242
rect -73473 -29858 -73177 -29242
rect -72473 -29858 -72177 -29242
rect -71473 -29858 -71177 -29242
rect -70473 -29858 -70177 -29242
rect -69473 -29858 -69177 -29242
rect -68473 -29858 -68177 -29242
rect -67473 -29858 -67177 -29242
rect -66473 -29858 -66177 -29242
rect -65473 -29858 -65177 -29242
rect -64473 -29858 -64177 -29242
rect -63473 -29858 -63177 -29242
rect -62473 -29858 -62177 -29242
rect -61473 -29858 -61177 -29242
rect -60473 -29858 -60177 -29242
rect -59473 -29858 -59177 -29242
rect -58473 -29858 -58177 -29242
rect -57473 -29858 -57177 -29242
rect -56473 -29858 -56177 -29242
rect -55473 -29858 -55177 -29242
rect -54473 -29858 -54177 -29242
rect -53473 -29858 -53177 -29242
rect -52473 -29858 -52177 -29242
rect -51473 -29858 -51177 -29242
rect -50473 -29858 -50177 -29242
rect -49473 -29858 -49177 -29242
rect 8627 -29858 8923 -29242
rect 9627 -29858 9923 -29242
rect 10627 -29858 10923 -29242
rect 11627 -29858 11923 -29242
rect 12627 -29858 12923 -29242
rect 13627 -29858 13923 -29242
rect 14627 -29858 14923 -29242
rect 15627 -29858 15923 -29242
rect 16627 -29858 16923 -29242
rect 17627 -29858 17923 -29242
rect 18627 -29858 18923 -29242
rect 19627 -29858 19923 -29242
rect 20627 -29858 20923 -29242
rect 21627 -29858 21923 -29242
rect 22627 -29858 22923 -29242
rect 23627 -29858 23923 -29242
rect 24627 -29858 24923 -29242
rect 25627 -29858 25923 -29242
rect 26627 -29858 26923 -29242
rect 27627 -29858 27923 -29242
rect 28627 -29858 28923 -29242
rect 29627 -29858 29923 -29242
rect 30627 -29858 30923 -29242
rect 31627 -29858 31923 -29242
rect 32627 -29858 32923 -29242
rect 33627 -29858 33923 -29242
rect -74813 -30198 -74517 -29902
rect -74473 -29928 -74177 -29902
rect -74473 -30172 -74447 -29928
rect -74447 -30172 -74203 -29928
rect -74203 -30172 -74177 -29928
rect -74473 -30198 -74177 -30172
rect -74133 -30198 -73517 -29902
rect -73473 -29928 -73177 -29902
rect -73473 -30172 -73447 -29928
rect -73447 -30172 -73203 -29928
rect -73203 -30172 -73177 -29928
rect -73473 -30198 -73177 -30172
rect -73133 -30198 -72517 -29902
rect -72473 -29928 -72177 -29902
rect -72473 -30172 -72447 -29928
rect -72447 -30172 -72203 -29928
rect -72203 -30172 -72177 -29928
rect -72473 -30198 -72177 -30172
rect -72133 -30198 -71517 -29902
rect -71473 -29928 -71177 -29902
rect -71473 -30172 -71447 -29928
rect -71447 -30172 -71203 -29928
rect -71203 -30172 -71177 -29928
rect -71473 -30198 -71177 -30172
rect -71133 -30198 -70517 -29902
rect -70473 -29928 -70177 -29902
rect -70473 -30172 -70447 -29928
rect -70447 -30172 -70203 -29928
rect -70203 -30172 -70177 -29928
rect -70473 -30198 -70177 -30172
rect -70133 -30198 -69517 -29902
rect -69473 -29928 -69177 -29902
rect -69473 -30172 -69447 -29928
rect -69447 -30172 -69203 -29928
rect -69203 -30172 -69177 -29928
rect -69473 -30198 -69177 -30172
rect -69133 -30198 -68517 -29902
rect -68473 -29928 -68177 -29902
rect -68473 -30172 -68447 -29928
rect -68447 -30172 -68203 -29928
rect -68203 -30172 -68177 -29928
rect -68473 -30198 -68177 -30172
rect -68133 -30198 -67517 -29902
rect -67473 -29928 -67177 -29902
rect -67473 -30172 -67447 -29928
rect -67447 -30172 -67203 -29928
rect -67203 -30172 -67177 -29928
rect -67473 -30198 -67177 -30172
rect -67133 -30198 -66517 -29902
rect -66473 -29928 -66177 -29902
rect -66473 -30172 -66447 -29928
rect -66447 -30172 -66203 -29928
rect -66203 -30172 -66177 -29928
rect -66473 -30198 -66177 -30172
rect -66133 -30198 -65517 -29902
rect -65473 -29928 -65177 -29902
rect -65473 -30172 -65447 -29928
rect -65447 -30172 -65203 -29928
rect -65203 -30172 -65177 -29928
rect -65473 -30198 -65177 -30172
rect -65133 -30198 -64517 -29902
rect -64473 -29928 -64177 -29902
rect -64473 -30172 -64447 -29928
rect -64447 -30172 -64203 -29928
rect -64203 -30172 -64177 -29928
rect -64473 -30198 -64177 -30172
rect -64133 -30198 -63517 -29902
rect -63473 -29928 -63177 -29902
rect -63473 -30172 -63447 -29928
rect -63447 -30172 -63203 -29928
rect -63203 -30172 -63177 -29928
rect -63473 -30198 -63177 -30172
rect -63133 -30198 -62517 -29902
rect -62473 -29928 -62177 -29902
rect -62473 -30172 -62447 -29928
rect -62447 -30172 -62203 -29928
rect -62203 -30172 -62177 -29928
rect -62473 -30198 -62177 -30172
rect -62133 -30198 -61517 -29902
rect -61473 -29928 -61177 -29902
rect -61473 -30172 -61447 -29928
rect -61447 -30172 -61203 -29928
rect -61203 -30172 -61177 -29928
rect -61473 -30198 -61177 -30172
rect -61133 -30198 -60517 -29902
rect -60473 -29928 -60177 -29902
rect -60473 -30172 -60447 -29928
rect -60447 -30172 -60203 -29928
rect -60203 -30172 -60177 -29928
rect -60473 -30198 -60177 -30172
rect -60133 -30198 -59517 -29902
rect -59473 -29928 -59177 -29902
rect -59473 -30172 -59447 -29928
rect -59447 -30172 -59203 -29928
rect -59203 -30172 -59177 -29928
rect -59473 -30198 -59177 -30172
rect -59133 -30198 -58517 -29902
rect -58473 -29928 -58177 -29902
rect -58473 -30172 -58447 -29928
rect -58447 -30172 -58203 -29928
rect -58203 -30172 -58177 -29928
rect -58473 -30198 -58177 -30172
rect -58133 -30198 -57517 -29902
rect -57473 -29928 -57177 -29902
rect -57473 -30172 -57447 -29928
rect -57447 -30172 -57203 -29928
rect -57203 -30172 -57177 -29928
rect -57473 -30198 -57177 -30172
rect -57133 -30198 -56517 -29902
rect -56473 -29928 -56177 -29902
rect -56473 -30172 -56447 -29928
rect -56447 -30172 -56203 -29928
rect -56203 -30172 -56177 -29928
rect -56473 -30198 -56177 -30172
rect -56133 -30198 -55517 -29902
rect -55473 -29928 -55177 -29902
rect -55473 -30172 -55447 -29928
rect -55447 -30172 -55203 -29928
rect -55203 -30172 -55177 -29928
rect -55473 -30198 -55177 -30172
rect -55133 -30198 -54517 -29902
rect -54473 -29928 -54177 -29902
rect -54473 -30172 -54447 -29928
rect -54447 -30172 -54203 -29928
rect -54203 -30172 -54177 -29928
rect -54473 -30198 -54177 -30172
rect -54133 -30198 -53517 -29902
rect -53473 -29928 -53177 -29902
rect -53473 -30172 -53447 -29928
rect -53447 -30172 -53203 -29928
rect -53203 -30172 -53177 -29928
rect -53473 -30198 -53177 -30172
rect -53133 -30198 -52517 -29902
rect -52473 -29928 -52177 -29902
rect -52473 -30172 -52447 -29928
rect -52447 -30172 -52203 -29928
rect -52203 -30172 -52177 -29928
rect -52473 -30198 -52177 -30172
rect -52133 -30198 -51517 -29902
rect -51473 -29928 -51177 -29902
rect -51473 -30172 -51447 -29928
rect -51447 -30172 -51203 -29928
rect -51203 -30172 -51177 -29928
rect -51473 -30198 -51177 -30172
rect -51133 -30198 -50517 -29902
rect -50473 -29928 -50177 -29902
rect -50473 -30172 -50447 -29928
rect -50447 -30172 -50203 -29928
rect -50203 -30172 -50177 -29928
rect -50473 -30198 -50177 -30172
rect -50133 -30198 -49517 -29902
rect -49473 -29928 -49177 -29902
rect -49473 -30172 -49447 -29928
rect -49447 -30172 -49203 -29928
rect -49203 -30172 -49177 -29928
rect -49473 -30198 -49177 -30172
rect -49133 -30198 -48837 -29902
rect 8287 -30198 8583 -29902
rect 8627 -29928 8923 -29902
rect 8627 -30172 8653 -29928
rect 8653 -30172 8897 -29928
rect 8897 -30172 8923 -29928
rect 8627 -30198 8923 -30172
rect 8967 -30198 9583 -29902
rect 9627 -29928 9923 -29902
rect 9627 -30172 9653 -29928
rect 9653 -30172 9897 -29928
rect 9897 -30172 9923 -29928
rect 9627 -30198 9923 -30172
rect 9967 -30198 10583 -29902
rect 10627 -29928 10923 -29902
rect 10627 -30172 10653 -29928
rect 10653 -30172 10897 -29928
rect 10897 -30172 10923 -29928
rect 10627 -30198 10923 -30172
rect 10967 -30198 11583 -29902
rect 11627 -29928 11923 -29902
rect 11627 -30172 11653 -29928
rect 11653 -30172 11897 -29928
rect 11897 -30172 11923 -29928
rect 11627 -30198 11923 -30172
rect 11967 -30198 12583 -29902
rect 12627 -29928 12923 -29902
rect 12627 -30172 12653 -29928
rect 12653 -30172 12897 -29928
rect 12897 -30172 12923 -29928
rect 12627 -30198 12923 -30172
rect 12967 -30198 13583 -29902
rect 13627 -29928 13923 -29902
rect 13627 -30172 13653 -29928
rect 13653 -30172 13897 -29928
rect 13897 -30172 13923 -29928
rect 13627 -30198 13923 -30172
rect 13967 -30198 14583 -29902
rect 14627 -29928 14923 -29902
rect 14627 -30172 14653 -29928
rect 14653 -30172 14897 -29928
rect 14897 -30172 14923 -29928
rect 14627 -30198 14923 -30172
rect 14967 -30198 15583 -29902
rect 15627 -29928 15923 -29902
rect 15627 -30172 15653 -29928
rect 15653 -30172 15897 -29928
rect 15897 -30172 15923 -29928
rect 15627 -30198 15923 -30172
rect 15967 -30198 16583 -29902
rect 16627 -29928 16923 -29902
rect 16627 -30172 16653 -29928
rect 16653 -30172 16897 -29928
rect 16897 -30172 16923 -29928
rect 16627 -30198 16923 -30172
rect 16967 -30198 17583 -29902
rect 17627 -29928 17923 -29902
rect 17627 -30172 17653 -29928
rect 17653 -30172 17897 -29928
rect 17897 -30172 17923 -29928
rect 17627 -30198 17923 -30172
rect 17967 -30198 18583 -29902
rect 18627 -29928 18923 -29902
rect 18627 -30172 18653 -29928
rect 18653 -30172 18897 -29928
rect 18897 -30172 18923 -29928
rect 18627 -30198 18923 -30172
rect 18967 -30198 19583 -29902
rect 19627 -29928 19923 -29902
rect 19627 -30172 19653 -29928
rect 19653 -30172 19897 -29928
rect 19897 -30172 19923 -29928
rect 19627 -30198 19923 -30172
rect 19967 -30198 20583 -29902
rect 20627 -29928 20923 -29902
rect 20627 -30172 20653 -29928
rect 20653 -30172 20897 -29928
rect 20897 -30172 20923 -29928
rect 20627 -30198 20923 -30172
rect 20967 -30198 21583 -29902
rect 21627 -29928 21923 -29902
rect 21627 -30172 21653 -29928
rect 21653 -30172 21897 -29928
rect 21897 -30172 21923 -29928
rect 21627 -30198 21923 -30172
rect 21967 -30198 22583 -29902
rect 22627 -29928 22923 -29902
rect 22627 -30172 22653 -29928
rect 22653 -30172 22897 -29928
rect 22897 -30172 22923 -29928
rect 22627 -30198 22923 -30172
rect 22967 -30198 23583 -29902
rect 23627 -29928 23923 -29902
rect 23627 -30172 23653 -29928
rect 23653 -30172 23897 -29928
rect 23897 -30172 23923 -29928
rect 23627 -30198 23923 -30172
rect 23967 -30198 24583 -29902
rect 24627 -29928 24923 -29902
rect 24627 -30172 24653 -29928
rect 24653 -30172 24897 -29928
rect 24897 -30172 24923 -29928
rect 24627 -30198 24923 -30172
rect 24967 -30198 25583 -29902
rect 25627 -29928 25923 -29902
rect 25627 -30172 25653 -29928
rect 25653 -30172 25897 -29928
rect 25897 -30172 25923 -29928
rect 25627 -30198 25923 -30172
rect 25967 -30198 26583 -29902
rect 26627 -29928 26923 -29902
rect 26627 -30172 26653 -29928
rect 26653 -30172 26897 -29928
rect 26897 -30172 26923 -29928
rect 26627 -30198 26923 -30172
rect 26967 -30198 27583 -29902
rect 27627 -29928 27923 -29902
rect 27627 -30172 27653 -29928
rect 27653 -30172 27897 -29928
rect 27897 -30172 27923 -29928
rect 27627 -30198 27923 -30172
rect 27967 -30198 28583 -29902
rect 28627 -29928 28923 -29902
rect 28627 -30172 28653 -29928
rect 28653 -30172 28897 -29928
rect 28897 -30172 28923 -29928
rect 28627 -30198 28923 -30172
rect 28967 -30198 29583 -29902
rect 29627 -29928 29923 -29902
rect 29627 -30172 29653 -29928
rect 29653 -30172 29897 -29928
rect 29897 -30172 29923 -29928
rect 29627 -30198 29923 -30172
rect 29967 -30198 30583 -29902
rect 30627 -29928 30923 -29902
rect 30627 -30172 30653 -29928
rect 30653 -30172 30897 -29928
rect 30897 -30172 30923 -29928
rect 30627 -30198 30923 -30172
rect 30967 -30198 31583 -29902
rect 31627 -29928 31923 -29902
rect 31627 -30172 31653 -29928
rect 31653 -30172 31897 -29928
rect 31897 -30172 31923 -29928
rect 31627 -30198 31923 -30172
rect 31967 -30198 32583 -29902
rect 32627 -29928 32923 -29902
rect 32627 -30172 32653 -29928
rect 32653 -30172 32897 -29928
rect 32897 -30172 32923 -29928
rect 32627 -30198 32923 -30172
rect 32967 -30198 33583 -29902
rect 33627 -29928 33923 -29902
rect 33627 -30172 33653 -29928
rect 33653 -30172 33897 -29928
rect 33897 -30172 33923 -29928
rect 33627 -30198 33923 -30172
rect 33967 -30198 34263 -29902
rect -74473 -30858 -74177 -30242
rect -73473 -30858 -73177 -30242
rect -72473 -30858 -72177 -30242
rect -71473 -30858 -71177 -30242
rect -70473 -30858 -70177 -30242
rect -69473 -30858 -69177 -30242
rect -68473 -30858 -68177 -30242
rect -67473 -30858 -67177 -30242
rect -66473 -30858 -66177 -30242
rect -65473 -30858 -65177 -30242
rect -64473 -30858 -64177 -30242
rect -63473 -30858 -63177 -30242
rect -62473 -30858 -62177 -30242
rect -61473 -30858 -61177 -30242
rect -60473 -30858 -60177 -30242
rect -59473 -30858 -59177 -30242
rect -58473 -30858 -58177 -30242
rect -57473 -30858 -57177 -30242
rect -56473 -30858 -56177 -30242
rect -55473 -30858 -55177 -30242
rect -54473 -30858 -54177 -30242
rect -53473 -30858 -53177 -30242
rect -52473 -30858 -52177 -30242
rect -51473 -30858 -51177 -30242
rect -50473 -30858 -50177 -30242
rect -49473 -30858 -49177 -30242
rect 8627 -30858 8923 -30242
rect 9627 -30858 9923 -30242
rect 10627 -30858 10923 -30242
rect 11627 -30858 11923 -30242
rect 12627 -30858 12923 -30242
rect 13627 -30858 13923 -30242
rect 14627 -30858 14923 -30242
rect 15627 -30858 15923 -30242
rect 16627 -30858 16923 -30242
rect 17627 -30858 17923 -30242
rect 18627 -30858 18923 -30242
rect 19627 -30858 19923 -30242
rect 20627 -30858 20923 -30242
rect 21627 -30858 21923 -30242
rect 22627 -30858 22923 -30242
rect 23627 -30858 23923 -30242
rect 24627 -30858 24923 -30242
rect 25627 -30858 25923 -30242
rect 26627 -30858 26923 -30242
rect 27627 -30858 27923 -30242
rect 28627 -30858 28923 -30242
rect 29627 -30858 29923 -30242
rect 30627 -30858 30923 -30242
rect 31627 -30858 31923 -30242
rect 32627 -30858 32923 -30242
rect 33627 -30858 33923 -30242
rect -74813 -31198 -74517 -30902
rect -74473 -30928 -74177 -30902
rect -74473 -31172 -74447 -30928
rect -74447 -31172 -74203 -30928
rect -74203 -31172 -74177 -30928
rect -74473 -31198 -74177 -31172
rect -74133 -31198 -73517 -30902
rect -73473 -30928 -73177 -30902
rect -73473 -31172 -73447 -30928
rect -73447 -31172 -73203 -30928
rect -73203 -31172 -73177 -30928
rect -73473 -31198 -73177 -31172
rect -73133 -31198 -72517 -30902
rect -72473 -30928 -72177 -30902
rect -72473 -31172 -72447 -30928
rect -72447 -31172 -72203 -30928
rect -72203 -31172 -72177 -30928
rect -72473 -31198 -72177 -31172
rect -72133 -31198 -71517 -30902
rect -71473 -30928 -71177 -30902
rect -71473 -31172 -71447 -30928
rect -71447 -31172 -71203 -30928
rect -71203 -31172 -71177 -30928
rect -71473 -31198 -71177 -31172
rect -71133 -31198 -70517 -30902
rect -70473 -30928 -70177 -30902
rect -70473 -31172 -70447 -30928
rect -70447 -31172 -70203 -30928
rect -70203 -31172 -70177 -30928
rect -70473 -31198 -70177 -31172
rect -70133 -31198 -69517 -30902
rect -69473 -30928 -69177 -30902
rect -69473 -31172 -69447 -30928
rect -69447 -31172 -69203 -30928
rect -69203 -31172 -69177 -30928
rect -69473 -31198 -69177 -31172
rect -69133 -31198 -68517 -30902
rect -68473 -30928 -68177 -30902
rect -68473 -31172 -68447 -30928
rect -68447 -31172 -68203 -30928
rect -68203 -31172 -68177 -30928
rect -68473 -31198 -68177 -31172
rect -68133 -31198 -67517 -30902
rect -67473 -30928 -67177 -30902
rect -67473 -31172 -67447 -30928
rect -67447 -31172 -67203 -30928
rect -67203 -31172 -67177 -30928
rect -67473 -31198 -67177 -31172
rect -67133 -31198 -66517 -30902
rect -66473 -30928 -66177 -30902
rect -66473 -31172 -66447 -30928
rect -66447 -31172 -66203 -30928
rect -66203 -31172 -66177 -30928
rect -66473 -31198 -66177 -31172
rect -66133 -31198 -65517 -30902
rect -65473 -30928 -65177 -30902
rect -65473 -31172 -65447 -30928
rect -65447 -31172 -65203 -30928
rect -65203 -31172 -65177 -30928
rect -65473 -31198 -65177 -31172
rect -65133 -31198 -64517 -30902
rect -64473 -30928 -64177 -30902
rect -64473 -31172 -64447 -30928
rect -64447 -31172 -64203 -30928
rect -64203 -31172 -64177 -30928
rect -64473 -31198 -64177 -31172
rect -64133 -31198 -63517 -30902
rect -63473 -30928 -63177 -30902
rect -63473 -31172 -63447 -30928
rect -63447 -31172 -63203 -30928
rect -63203 -31172 -63177 -30928
rect -63473 -31198 -63177 -31172
rect -63133 -31198 -62517 -30902
rect -62473 -30928 -62177 -30902
rect -62473 -31172 -62447 -30928
rect -62447 -31172 -62203 -30928
rect -62203 -31172 -62177 -30928
rect -62473 -31198 -62177 -31172
rect -62133 -31198 -61517 -30902
rect -61473 -30928 -61177 -30902
rect -61473 -31172 -61447 -30928
rect -61447 -31172 -61203 -30928
rect -61203 -31172 -61177 -30928
rect -61473 -31198 -61177 -31172
rect -61133 -31198 -60517 -30902
rect -60473 -30928 -60177 -30902
rect -60473 -31172 -60447 -30928
rect -60447 -31172 -60203 -30928
rect -60203 -31172 -60177 -30928
rect -60473 -31198 -60177 -31172
rect -60133 -31198 -59517 -30902
rect -59473 -30928 -59177 -30902
rect -59473 -31172 -59447 -30928
rect -59447 -31172 -59203 -30928
rect -59203 -31172 -59177 -30928
rect -59473 -31198 -59177 -31172
rect -59133 -31198 -58517 -30902
rect -58473 -30928 -58177 -30902
rect -58473 -31172 -58447 -30928
rect -58447 -31172 -58203 -30928
rect -58203 -31172 -58177 -30928
rect -58473 -31198 -58177 -31172
rect -58133 -31198 -57517 -30902
rect -57473 -30928 -57177 -30902
rect -57473 -31172 -57447 -30928
rect -57447 -31172 -57203 -30928
rect -57203 -31172 -57177 -30928
rect -57473 -31198 -57177 -31172
rect -57133 -31198 -56517 -30902
rect -56473 -30928 -56177 -30902
rect -56473 -31172 -56447 -30928
rect -56447 -31172 -56203 -30928
rect -56203 -31172 -56177 -30928
rect -56473 -31198 -56177 -31172
rect -56133 -31198 -55517 -30902
rect -55473 -30928 -55177 -30902
rect -55473 -31172 -55447 -30928
rect -55447 -31172 -55203 -30928
rect -55203 -31172 -55177 -30928
rect -55473 -31198 -55177 -31172
rect -55133 -31198 -54517 -30902
rect -54473 -30928 -54177 -30902
rect -54473 -31172 -54447 -30928
rect -54447 -31172 -54203 -30928
rect -54203 -31172 -54177 -30928
rect -54473 -31198 -54177 -31172
rect -54133 -31198 -53517 -30902
rect -53473 -30928 -53177 -30902
rect -53473 -31172 -53447 -30928
rect -53447 -31172 -53203 -30928
rect -53203 -31172 -53177 -30928
rect -53473 -31198 -53177 -31172
rect -53133 -31198 -52517 -30902
rect -52473 -30928 -52177 -30902
rect -52473 -31172 -52447 -30928
rect -52447 -31172 -52203 -30928
rect -52203 -31172 -52177 -30928
rect -52473 -31198 -52177 -31172
rect -52133 -31198 -51517 -30902
rect -51473 -30928 -51177 -30902
rect -51473 -31172 -51447 -30928
rect -51447 -31172 -51203 -30928
rect -51203 -31172 -51177 -30928
rect -51473 -31198 -51177 -31172
rect -51133 -31198 -50517 -30902
rect -50473 -30928 -50177 -30902
rect -50473 -31172 -50447 -30928
rect -50447 -31172 -50203 -30928
rect -50203 -31172 -50177 -30928
rect -50473 -31198 -50177 -31172
rect -50133 -31198 -49517 -30902
rect -49473 -30928 -49177 -30902
rect -49473 -31172 -49447 -30928
rect -49447 -31172 -49203 -30928
rect -49203 -31172 -49177 -30928
rect -49473 -31198 -49177 -31172
rect -49133 -31198 -48837 -30902
rect 8287 -31198 8583 -30902
rect 8627 -30928 8923 -30902
rect 8627 -31172 8653 -30928
rect 8653 -31172 8897 -30928
rect 8897 -31172 8923 -30928
rect 8627 -31198 8923 -31172
rect 8967 -31198 9583 -30902
rect 9627 -30928 9923 -30902
rect 9627 -31172 9653 -30928
rect 9653 -31172 9897 -30928
rect 9897 -31172 9923 -30928
rect 9627 -31198 9923 -31172
rect 9967 -31198 10583 -30902
rect 10627 -30928 10923 -30902
rect 10627 -31172 10653 -30928
rect 10653 -31172 10897 -30928
rect 10897 -31172 10923 -30928
rect 10627 -31198 10923 -31172
rect 10967 -31198 11583 -30902
rect 11627 -30928 11923 -30902
rect 11627 -31172 11653 -30928
rect 11653 -31172 11897 -30928
rect 11897 -31172 11923 -30928
rect 11627 -31198 11923 -31172
rect 11967 -31198 12583 -30902
rect 12627 -30928 12923 -30902
rect 12627 -31172 12653 -30928
rect 12653 -31172 12897 -30928
rect 12897 -31172 12923 -30928
rect 12627 -31198 12923 -31172
rect 12967 -31198 13583 -30902
rect 13627 -30928 13923 -30902
rect 13627 -31172 13653 -30928
rect 13653 -31172 13897 -30928
rect 13897 -31172 13923 -30928
rect 13627 -31198 13923 -31172
rect 13967 -31198 14583 -30902
rect 14627 -30928 14923 -30902
rect 14627 -31172 14653 -30928
rect 14653 -31172 14897 -30928
rect 14897 -31172 14923 -30928
rect 14627 -31198 14923 -31172
rect 14967 -31198 15583 -30902
rect 15627 -30928 15923 -30902
rect 15627 -31172 15653 -30928
rect 15653 -31172 15897 -30928
rect 15897 -31172 15923 -30928
rect 15627 -31198 15923 -31172
rect 15967 -31198 16583 -30902
rect 16627 -30928 16923 -30902
rect 16627 -31172 16653 -30928
rect 16653 -31172 16897 -30928
rect 16897 -31172 16923 -30928
rect 16627 -31198 16923 -31172
rect 16967 -31198 17583 -30902
rect 17627 -30928 17923 -30902
rect 17627 -31172 17653 -30928
rect 17653 -31172 17897 -30928
rect 17897 -31172 17923 -30928
rect 17627 -31198 17923 -31172
rect 17967 -31198 18583 -30902
rect 18627 -30928 18923 -30902
rect 18627 -31172 18653 -30928
rect 18653 -31172 18897 -30928
rect 18897 -31172 18923 -30928
rect 18627 -31198 18923 -31172
rect 18967 -31198 19583 -30902
rect 19627 -30928 19923 -30902
rect 19627 -31172 19653 -30928
rect 19653 -31172 19897 -30928
rect 19897 -31172 19923 -30928
rect 19627 -31198 19923 -31172
rect 19967 -31198 20583 -30902
rect 20627 -30928 20923 -30902
rect 20627 -31172 20653 -30928
rect 20653 -31172 20897 -30928
rect 20897 -31172 20923 -30928
rect 20627 -31198 20923 -31172
rect 20967 -31198 21583 -30902
rect 21627 -30928 21923 -30902
rect 21627 -31172 21653 -30928
rect 21653 -31172 21897 -30928
rect 21897 -31172 21923 -30928
rect 21627 -31198 21923 -31172
rect 21967 -31198 22583 -30902
rect 22627 -30928 22923 -30902
rect 22627 -31172 22653 -30928
rect 22653 -31172 22897 -30928
rect 22897 -31172 22923 -30928
rect 22627 -31198 22923 -31172
rect 22967 -31198 23583 -30902
rect 23627 -30928 23923 -30902
rect 23627 -31172 23653 -30928
rect 23653 -31172 23897 -30928
rect 23897 -31172 23923 -30928
rect 23627 -31198 23923 -31172
rect 23967 -31198 24583 -30902
rect 24627 -30928 24923 -30902
rect 24627 -31172 24653 -30928
rect 24653 -31172 24897 -30928
rect 24897 -31172 24923 -30928
rect 24627 -31198 24923 -31172
rect 24967 -31198 25583 -30902
rect 25627 -30928 25923 -30902
rect 25627 -31172 25653 -30928
rect 25653 -31172 25897 -30928
rect 25897 -31172 25923 -30928
rect 25627 -31198 25923 -31172
rect 25967 -31198 26583 -30902
rect 26627 -30928 26923 -30902
rect 26627 -31172 26653 -30928
rect 26653 -31172 26897 -30928
rect 26897 -31172 26923 -30928
rect 26627 -31198 26923 -31172
rect 26967 -31198 27583 -30902
rect 27627 -30928 27923 -30902
rect 27627 -31172 27653 -30928
rect 27653 -31172 27897 -30928
rect 27897 -31172 27923 -30928
rect 27627 -31198 27923 -31172
rect 27967 -31198 28583 -30902
rect 28627 -30928 28923 -30902
rect 28627 -31172 28653 -30928
rect 28653 -31172 28897 -30928
rect 28897 -31172 28923 -30928
rect 28627 -31198 28923 -31172
rect 28967 -31198 29583 -30902
rect 29627 -30928 29923 -30902
rect 29627 -31172 29653 -30928
rect 29653 -31172 29897 -30928
rect 29897 -31172 29923 -30928
rect 29627 -31198 29923 -31172
rect 29967 -31198 30583 -30902
rect 30627 -30928 30923 -30902
rect 30627 -31172 30653 -30928
rect 30653 -31172 30897 -30928
rect 30897 -31172 30923 -30928
rect 30627 -31198 30923 -31172
rect 30967 -31198 31583 -30902
rect 31627 -30928 31923 -30902
rect 31627 -31172 31653 -30928
rect 31653 -31172 31897 -30928
rect 31897 -31172 31923 -30928
rect 31627 -31198 31923 -31172
rect 31967 -31198 32583 -30902
rect 32627 -30928 32923 -30902
rect 32627 -31172 32653 -30928
rect 32653 -31172 32897 -30928
rect 32897 -31172 32923 -30928
rect 32627 -31198 32923 -31172
rect 32967 -31198 33583 -30902
rect 33627 -30928 33923 -30902
rect 33627 -31172 33653 -30928
rect 33653 -31172 33897 -30928
rect 33897 -31172 33923 -30928
rect 33627 -31198 33923 -31172
rect 33967 -31198 34263 -30902
rect -74473 -31858 -74177 -31242
rect -73473 -31858 -73177 -31242
rect -72473 -31858 -72177 -31242
rect -71473 -31858 -71177 -31242
rect -70473 -31858 -70177 -31242
rect -69473 -31858 -69177 -31242
rect -68473 -31858 -68177 -31242
rect -67473 -31858 -67177 -31242
rect -66473 -31858 -66177 -31242
rect -65473 -31858 -65177 -31242
rect -64473 -31858 -64177 -31242
rect -63473 -31858 -63177 -31242
rect -62473 -31858 -62177 -31242
rect -61473 -31858 -61177 -31242
rect -60473 -31858 -60177 -31242
rect -59473 -31858 -59177 -31242
rect -58473 -31858 -58177 -31242
rect -57473 -31858 -57177 -31242
rect -56473 -31858 -56177 -31242
rect -55473 -31858 -55177 -31242
rect -54473 -31858 -54177 -31242
rect -53473 -31858 -53177 -31242
rect -52473 -31858 -52177 -31242
rect -51473 -31858 -51177 -31242
rect -50473 -31858 -50177 -31242
rect -49473 -31858 -49177 -31242
rect 8627 -31858 8923 -31242
rect 9627 -31858 9923 -31242
rect 10627 -31858 10923 -31242
rect 11627 -31858 11923 -31242
rect 12627 -31858 12923 -31242
rect 13627 -31858 13923 -31242
rect 14627 -31858 14923 -31242
rect 15627 -31858 15923 -31242
rect 16627 -31858 16923 -31242
rect 17627 -31858 17923 -31242
rect 18627 -31858 18923 -31242
rect 19627 -31858 19923 -31242
rect 20627 -31858 20923 -31242
rect 21627 -31858 21923 -31242
rect 22627 -31858 22923 -31242
rect 23627 -31858 23923 -31242
rect 24627 -31858 24923 -31242
rect 25627 -31858 25923 -31242
rect 26627 -31858 26923 -31242
rect 27627 -31858 27923 -31242
rect 28627 -31858 28923 -31242
rect 29627 -31858 29923 -31242
rect 30627 -31858 30923 -31242
rect 31627 -31858 31923 -31242
rect 32627 -31858 32923 -31242
rect 33627 -31858 33923 -31242
rect -74813 -32198 -74517 -31902
rect -74473 -31928 -74177 -31902
rect -74473 -32172 -74447 -31928
rect -74447 -32172 -74203 -31928
rect -74203 -32172 -74177 -31928
rect -74473 -32198 -74177 -32172
rect -74133 -32198 -73517 -31902
rect -73473 -31928 -73177 -31902
rect -73473 -32172 -73447 -31928
rect -73447 -32172 -73203 -31928
rect -73203 -32172 -73177 -31928
rect -73473 -32198 -73177 -32172
rect -73133 -32198 -72517 -31902
rect -72473 -31928 -72177 -31902
rect -72473 -32172 -72447 -31928
rect -72447 -32172 -72203 -31928
rect -72203 -32172 -72177 -31928
rect -72473 -32198 -72177 -32172
rect -72133 -32198 -71517 -31902
rect -71473 -31928 -71177 -31902
rect -71473 -32172 -71447 -31928
rect -71447 -32172 -71203 -31928
rect -71203 -32172 -71177 -31928
rect -71473 -32198 -71177 -32172
rect -71133 -32198 -70517 -31902
rect -70473 -31928 -70177 -31902
rect -70473 -32172 -70447 -31928
rect -70447 -32172 -70203 -31928
rect -70203 -32172 -70177 -31928
rect -70473 -32198 -70177 -32172
rect -70133 -32198 -69517 -31902
rect -69473 -31928 -69177 -31902
rect -69473 -32172 -69447 -31928
rect -69447 -32172 -69203 -31928
rect -69203 -32172 -69177 -31928
rect -69473 -32198 -69177 -32172
rect -69133 -32198 -68517 -31902
rect -68473 -31928 -68177 -31902
rect -68473 -32172 -68447 -31928
rect -68447 -32172 -68203 -31928
rect -68203 -32172 -68177 -31928
rect -68473 -32198 -68177 -32172
rect -68133 -32198 -67517 -31902
rect -67473 -31928 -67177 -31902
rect -67473 -32172 -67447 -31928
rect -67447 -32172 -67203 -31928
rect -67203 -32172 -67177 -31928
rect -67473 -32198 -67177 -32172
rect -67133 -32198 -66517 -31902
rect -66473 -31928 -66177 -31902
rect -66473 -32172 -66447 -31928
rect -66447 -32172 -66203 -31928
rect -66203 -32172 -66177 -31928
rect -66473 -32198 -66177 -32172
rect -66133 -32198 -65517 -31902
rect -65473 -31928 -65177 -31902
rect -65473 -32172 -65447 -31928
rect -65447 -32172 -65203 -31928
rect -65203 -32172 -65177 -31928
rect -65473 -32198 -65177 -32172
rect -65133 -32198 -64517 -31902
rect -64473 -31928 -64177 -31902
rect -64473 -32172 -64447 -31928
rect -64447 -32172 -64203 -31928
rect -64203 -32172 -64177 -31928
rect -64473 -32198 -64177 -32172
rect -64133 -32198 -63517 -31902
rect -63473 -31928 -63177 -31902
rect -63473 -32172 -63447 -31928
rect -63447 -32172 -63203 -31928
rect -63203 -32172 -63177 -31928
rect -63473 -32198 -63177 -32172
rect -63133 -32198 -62517 -31902
rect -62473 -31928 -62177 -31902
rect -62473 -32172 -62447 -31928
rect -62447 -32172 -62203 -31928
rect -62203 -32172 -62177 -31928
rect -62473 -32198 -62177 -32172
rect -62133 -32198 -61517 -31902
rect -61473 -31928 -61177 -31902
rect -61473 -32172 -61447 -31928
rect -61447 -32172 -61203 -31928
rect -61203 -32172 -61177 -31928
rect -61473 -32198 -61177 -32172
rect -61133 -32198 -60517 -31902
rect -60473 -31928 -60177 -31902
rect -60473 -32172 -60447 -31928
rect -60447 -32172 -60203 -31928
rect -60203 -32172 -60177 -31928
rect -60473 -32198 -60177 -32172
rect -60133 -32198 -59517 -31902
rect -59473 -31928 -59177 -31902
rect -59473 -32172 -59447 -31928
rect -59447 -32172 -59203 -31928
rect -59203 -32172 -59177 -31928
rect -59473 -32198 -59177 -32172
rect -59133 -32198 -58517 -31902
rect -58473 -31928 -58177 -31902
rect -58473 -32172 -58447 -31928
rect -58447 -32172 -58203 -31928
rect -58203 -32172 -58177 -31928
rect -58473 -32198 -58177 -32172
rect -58133 -32198 -57517 -31902
rect -57473 -31928 -57177 -31902
rect -57473 -32172 -57447 -31928
rect -57447 -32172 -57203 -31928
rect -57203 -32172 -57177 -31928
rect -57473 -32198 -57177 -32172
rect -57133 -32198 -56517 -31902
rect -56473 -31928 -56177 -31902
rect -56473 -32172 -56447 -31928
rect -56447 -32172 -56203 -31928
rect -56203 -32172 -56177 -31928
rect -56473 -32198 -56177 -32172
rect -56133 -32198 -55517 -31902
rect -55473 -31928 -55177 -31902
rect -55473 -32172 -55447 -31928
rect -55447 -32172 -55203 -31928
rect -55203 -32172 -55177 -31928
rect -55473 -32198 -55177 -32172
rect -55133 -32198 -54517 -31902
rect -54473 -31928 -54177 -31902
rect -54473 -32172 -54447 -31928
rect -54447 -32172 -54203 -31928
rect -54203 -32172 -54177 -31928
rect -54473 -32198 -54177 -32172
rect -54133 -32198 -53517 -31902
rect -53473 -31928 -53177 -31902
rect -53473 -32172 -53447 -31928
rect -53447 -32172 -53203 -31928
rect -53203 -32172 -53177 -31928
rect -53473 -32198 -53177 -32172
rect -53133 -32198 -52517 -31902
rect -52473 -31928 -52177 -31902
rect -52473 -32172 -52447 -31928
rect -52447 -32172 -52203 -31928
rect -52203 -32172 -52177 -31928
rect -52473 -32198 -52177 -32172
rect -52133 -32198 -51517 -31902
rect -51473 -31928 -51177 -31902
rect -51473 -32172 -51447 -31928
rect -51447 -32172 -51203 -31928
rect -51203 -32172 -51177 -31928
rect -51473 -32198 -51177 -32172
rect -51133 -32198 -50517 -31902
rect -50473 -31928 -50177 -31902
rect -50473 -32172 -50447 -31928
rect -50447 -32172 -50203 -31928
rect -50203 -32172 -50177 -31928
rect -50473 -32198 -50177 -32172
rect -50133 -32198 -49517 -31902
rect -49473 -31928 -49177 -31902
rect -49473 -32172 -49447 -31928
rect -49447 -32172 -49203 -31928
rect -49203 -32172 -49177 -31928
rect -49473 -32198 -49177 -32172
rect -49133 -32198 -48837 -31902
rect 8287 -32198 8583 -31902
rect 8627 -31928 8923 -31902
rect 8627 -32172 8653 -31928
rect 8653 -32172 8897 -31928
rect 8897 -32172 8923 -31928
rect 8627 -32198 8923 -32172
rect 8967 -32198 9583 -31902
rect 9627 -31928 9923 -31902
rect 9627 -32172 9653 -31928
rect 9653 -32172 9897 -31928
rect 9897 -32172 9923 -31928
rect 9627 -32198 9923 -32172
rect 9967 -32198 10583 -31902
rect 10627 -31928 10923 -31902
rect 10627 -32172 10653 -31928
rect 10653 -32172 10897 -31928
rect 10897 -32172 10923 -31928
rect 10627 -32198 10923 -32172
rect 10967 -32198 11583 -31902
rect 11627 -31928 11923 -31902
rect 11627 -32172 11653 -31928
rect 11653 -32172 11897 -31928
rect 11897 -32172 11923 -31928
rect 11627 -32198 11923 -32172
rect 11967 -32198 12583 -31902
rect 12627 -31928 12923 -31902
rect 12627 -32172 12653 -31928
rect 12653 -32172 12897 -31928
rect 12897 -32172 12923 -31928
rect 12627 -32198 12923 -32172
rect 12967 -32198 13583 -31902
rect 13627 -31928 13923 -31902
rect 13627 -32172 13653 -31928
rect 13653 -32172 13897 -31928
rect 13897 -32172 13923 -31928
rect 13627 -32198 13923 -32172
rect 13967 -32198 14583 -31902
rect 14627 -31928 14923 -31902
rect 14627 -32172 14653 -31928
rect 14653 -32172 14897 -31928
rect 14897 -32172 14923 -31928
rect 14627 -32198 14923 -32172
rect 14967 -32198 15583 -31902
rect 15627 -31928 15923 -31902
rect 15627 -32172 15653 -31928
rect 15653 -32172 15897 -31928
rect 15897 -32172 15923 -31928
rect 15627 -32198 15923 -32172
rect 15967 -32198 16583 -31902
rect 16627 -31928 16923 -31902
rect 16627 -32172 16653 -31928
rect 16653 -32172 16897 -31928
rect 16897 -32172 16923 -31928
rect 16627 -32198 16923 -32172
rect 16967 -32198 17583 -31902
rect 17627 -31928 17923 -31902
rect 17627 -32172 17653 -31928
rect 17653 -32172 17897 -31928
rect 17897 -32172 17923 -31928
rect 17627 -32198 17923 -32172
rect 17967 -32198 18583 -31902
rect 18627 -31928 18923 -31902
rect 18627 -32172 18653 -31928
rect 18653 -32172 18897 -31928
rect 18897 -32172 18923 -31928
rect 18627 -32198 18923 -32172
rect 18967 -32198 19583 -31902
rect 19627 -31928 19923 -31902
rect 19627 -32172 19653 -31928
rect 19653 -32172 19897 -31928
rect 19897 -32172 19923 -31928
rect 19627 -32198 19923 -32172
rect 19967 -32198 20583 -31902
rect 20627 -31928 20923 -31902
rect 20627 -32172 20653 -31928
rect 20653 -32172 20897 -31928
rect 20897 -32172 20923 -31928
rect 20627 -32198 20923 -32172
rect 20967 -32198 21583 -31902
rect 21627 -31928 21923 -31902
rect 21627 -32172 21653 -31928
rect 21653 -32172 21897 -31928
rect 21897 -32172 21923 -31928
rect 21627 -32198 21923 -32172
rect 21967 -32198 22583 -31902
rect 22627 -31928 22923 -31902
rect 22627 -32172 22653 -31928
rect 22653 -32172 22897 -31928
rect 22897 -32172 22923 -31928
rect 22627 -32198 22923 -32172
rect 22967 -32198 23583 -31902
rect 23627 -31928 23923 -31902
rect 23627 -32172 23653 -31928
rect 23653 -32172 23897 -31928
rect 23897 -32172 23923 -31928
rect 23627 -32198 23923 -32172
rect 23967 -32198 24583 -31902
rect 24627 -31928 24923 -31902
rect 24627 -32172 24653 -31928
rect 24653 -32172 24897 -31928
rect 24897 -32172 24923 -31928
rect 24627 -32198 24923 -32172
rect 24967 -32198 25583 -31902
rect 25627 -31928 25923 -31902
rect 25627 -32172 25653 -31928
rect 25653 -32172 25897 -31928
rect 25897 -32172 25923 -31928
rect 25627 -32198 25923 -32172
rect 25967 -32198 26583 -31902
rect 26627 -31928 26923 -31902
rect 26627 -32172 26653 -31928
rect 26653 -32172 26897 -31928
rect 26897 -32172 26923 -31928
rect 26627 -32198 26923 -32172
rect 26967 -32198 27583 -31902
rect 27627 -31928 27923 -31902
rect 27627 -32172 27653 -31928
rect 27653 -32172 27897 -31928
rect 27897 -32172 27923 -31928
rect 27627 -32198 27923 -32172
rect 27967 -32198 28583 -31902
rect 28627 -31928 28923 -31902
rect 28627 -32172 28653 -31928
rect 28653 -32172 28897 -31928
rect 28897 -32172 28923 -31928
rect 28627 -32198 28923 -32172
rect 28967 -32198 29583 -31902
rect 29627 -31928 29923 -31902
rect 29627 -32172 29653 -31928
rect 29653 -32172 29897 -31928
rect 29897 -32172 29923 -31928
rect 29627 -32198 29923 -32172
rect 29967 -32198 30583 -31902
rect 30627 -31928 30923 -31902
rect 30627 -32172 30653 -31928
rect 30653 -32172 30897 -31928
rect 30897 -32172 30923 -31928
rect 30627 -32198 30923 -32172
rect 30967 -32198 31583 -31902
rect 31627 -31928 31923 -31902
rect 31627 -32172 31653 -31928
rect 31653 -32172 31897 -31928
rect 31897 -32172 31923 -31928
rect 31627 -32198 31923 -32172
rect 31967 -32198 32583 -31902
rect 32627 -31928 32923 -31902
rect 32627 -32172 32653 -31928
rect 32653 -32172 32897 -31928
rect 32897 -32172 32923 -31928
rect 32627 -32198 32923 -32172
rect 32967 -32198 33583 -31902
rect 33627 -31928 33923 -31902
rect 33627 -32172 33653 -31928
rect 33653 -32172 33897 -31928
rect 33897 -32172 33923 -31928
rect 33627 -32198 33923 -32172
rect 33967 -32198 34263 -31902
rect -74473 -32858 -74177 -32242
rect -73473 -32858 -73177 -32242
rect -72473 -32858 -72177 -32242
rect -71473 -32858 -71177 -32242
rect -70473 -32858 -70177 -32242
rect -69473 -32858 -69177 -32242
rect -68473 -32858 -68177 -32242
rect -67473 -32858 -67177 -32242
rect -66473 -32858 -66177 -32242
rect -65473 -32858 -65177 -32242
rect -64473 -32858 -64177 -32242
rect -63473 -32858 -63177 -32242
rect -62473 -32858 -62177 -32242
rect -61473 -32858 -61177 -32242
rect -60473 -32858 -60177 -32242
rect -59473 -32858 -59177 -32242
rect -58473 -32858 -58177 -32242
rect -57473 -32858 -57177 -32242
rect -56473 -32858 -56177 -32242
rect -55473 -32858 -55177 -32242
rect -54473 -32858 -54177 -32242
rect -53473 -32858 -53177 -32242
rect -52473 -32858 -52177 -32242
rect -51473 -32858 -51177 -32242
rect -50473 -32858 -50177 -32242
rect -49473 -32858 -49177 -32242
rect -46228 -32604 -36332 -32602
rect -74813 -33198 -74517 -32902
rect -74473 -32928 -74177 -32902
rect -74473 -33172 -74447 -32928
rect -74447 -33172 -74203 -32928
rect -74203 -33172 -74177 -32928
rect -74473 -33198 -74177 -33172
rect -74133 -33198 -73517 -32902
rect -73473 -32928 -73177 -32902
rect -73473 -33172 -73447 -32928
rect -73447 -33172 -73203 -32928
rect -73203 -33172 -73177 -32928
rect -73473 -33198 -73177 -33172
rect -73133 -33198 -72517 -32902
rect -72473 -32928 -72177 -32902
rect -72473 -33172 -72447 -32928
rect -72447 -33172 -72203 -32928
rect -72203 -33172 -72177 -32928
rect -72473 -33198 -72177 -33172
rect -72133 -33198 -71517 -32902
rect -71473 -32928 -71177 -32902
rect -71473 -33172 -71447 -32928
rect -71447 -33172 -71203 -32928
rect -71203 -33172 -71177 -32928
rect -71473 -33198 -71177 -33172
rect -71133 -33198 -70517 -32902
rect -70473 -32928 -70177 -32902
rect -70473 -33172 -70447 -32928
rect -70447 -33172 -70203 -32928
rect -70203 -33172 -70177 -32928
rect -70473 -33198 -70177 -33172
rect -70133 -33198 -69517 -32902
rect -69473 -32928 -69177 -32902
rect -69473 -33172 -69447 -32928
rect -69447 -33172 -69203 -32928
rect -69203 -33172 -69177 -32928
rect -69473 -33198 -69177 -33172
rect -69133 -33198 -68517 -32902
rect -68473 -32928 -68177 -32902
rect -68473 -33172 -68447 -32928
rect -68447 -33172 -68203 -32928
rect -68203 -33172 -68177 -32928
rect -68473 -33198 -68177 -33172
rect -68133 -33198 -67517 -32902
rect -67473 -32928 -67177 -32902
rect -67473 -33172 -67447 -32928
rect -67447 -33172 -67203 -32928
rect -67203 -33172 -67177 -32928
rect -67473 -33198 -67177 -33172
rect -67133 -33198 -66517 -32902
rect -66473 -32928 -66177 -32902
rect -66473 -33172 -66447 -32928
rect -66447 -33172 -66203 -32928
rect -66203 -33172 -66177 -32928
rect -66473 -33198 -66177 -33172
rect -66133 -33198 -65517 -32902
rect -65473 -32928 -65177 -32902
rect -65473 -33172 -65447 -32928
rect -65447 -33172 -65203 -32928
rect -65203 -33172 -65177 -32928
rect -65473 -33198 -65177 -33172
rect -65133 -33198 -64517 -32902
rect -64473 -32928 -64177 -32902
rect -64473 -33172 -64447 -32928
rect -64447 -33172 -64203 -32928
rect -64203 -33172 -64177 -32928
rect -64473 -33198 -64177 -33172
rect -64133 -33198 -63517 -32902
rect -63473 -32928 -63177 -32902
rect -63473 -33172 -63447 -32928
rect -63447 -33172 -63203 -32928
rect -63203 -33172 -63177 -32928
rect -63473 -33198 -63177 -33172
rect -63133 -33198 -62517 -32902
rect -62473 -32928 -62177 -32902
rect -62473 -33172 -62447 -32928
rect -62447 -33172 -62203 -32928
rect -62203 -33172 -62177 -32928
rect -62473 -33198 -62177 -33172
rect -62133 -33198 -61517 -32902
rect -61473 -32928 -61177 -32902
rect -61473 -33172 -61447 -32928
rect -61447 -33172 -61203 -32928
rect -61203 -33172 -61177 -32928
rect -61473 -33198 -61177 -33172
rect -61133 -33198 -60517 -32902
rect -60473 -32928 -60177 -32902
rect -60473 -33172 -60447 -32928
rect -60447 -33172 -60203 -32928
rect -60203 -33172 -60177 -32928
rect -60473 -33198 -60177 -33172
rect -60133 -33198 -59517 -32902
rect -59473 -32928 -59177 -32902
rect -59473 -33172 -59447 -32928
rect -59447 -33172 -59203 -32928
rect -59203 -33172 -59177 -32928
rect -59473 -33198 -59177 -33172
rect -59133 -33198 -58517 -32902
rect -58473 -32928 -58177 -32902
rect -58473 -33172 -58447 -32928
rect -58447 -33172 -58203 -32928
rect -58203 -33172 -58177 -32928
rect -58473 -33198 -58177 -33172
rect -58133 -33198 -57517 -32902
rect -57473 -32928 -57177 -32902
rect -57473 -33172 -57447 -32928
rect -57447 -33172 -57203 -32928
rect -57203 -33172 -57177 -32928
rect -57473 -33198 -57177 -33172
rect -57133 -33198 -56517 -32902
rect -56473 -32928 -56177 -32902
rect -56473 -33172 -56447 -32928
rect -56447 -33172 -56203 -32928
rect -56203 -33172 -56177 -32928
rect -56473 -33198 -56177 -33172
rect -56133 -33198 -55517 -32902
rect -55473 -32928 -55177 -32902
rect -55473 -33172 -55447 -32928
rect -55447 -33172 -55203 -32928
rect -55203 -33172 -55177 -32928
rect -55473 -33198 -55177 -33172
rect -55133 -33198 -54517 -32902
rect -54473 -32928 -54177 -32902
rect -54473 -33172 -54447 -32928
rect -54447 -33172 -54203 -32928
rect -54203 -33172 -54177 -32928
rect -54473 -33198 -54177 -33172
rect -54133 -33198 -53517 -32902
rect -53473 -32928 -53177 -32902
rect -53473 -33172 -53447 -32928
rect -53447 -33172 -53203 -32928
rect -53203 -33172 -53177 -32928
rect -53473 -33198 -53177 -33172
rect -53133 -33198 -52517 -32902
rect -52473 -32928 -52177 -32902
rect -52473 -33172 -52447 -32928
rect -52447 -33172 -52203 -32928
rect -52203 -33172 -52177 -32928
rect -52473 -33198 -52177 -33172
rect -52133 -33198 -51517 -32902
rect -51473 -32928 -51177 -32902
rect -51473 -33172 -51447 -32928
rect -51447 -33172 -51203 -32928
rect -51203 -33172 -51177 -32928
rect -51473 -33198 -51177 -33172
rect -51133 -33198 -50517 -32902
rect -50473 -32928 -50177 -32902
rect -50473 -33172 -50447 -32928
rect -50447 -33172 -50203 -32928
rect -50203 -33172 -50177 -32928
rect -50473 -33198 -50177 -33172
rect -50133 -33198 -49517 -32902
rect -49473 -32928 -49177 -32902
rect -49473 -33172 -49447 -32928
rect -49447 -33172 -49203 -32928
rect -49203 -33172 -49177 -32928
rect -49473 -33198 -49177 -33172
rect -49133 -33198 -48837 -32902
rect -74473 -33858 -74177 -33242
rect -73473 -33858 -73177 -33242
rect -72473 -33858 -72177 -33242
rect -71473 -33858 -71177 -33242
rect -70473 -33858 -70177 -33242
rect -69473 -33858 -69177 -33242
rect -68473 -33858 -68177 -33242
rect -67473 -33858 -67177 -33242
rect -66473 -33858 -66177 -33242
rect -65473 -33858 -65177 -33242
rect -64473 -33858 -64177 -33242
rect -63473 -33858 -63177 -33242
rect -62473 -33858 -62177 -33242
rect -61473 -33858 -61177 -33242
rect -60473 -33858 -60177 -33242
rect -59473 -33858 -59177 -33242
rect -58473 -33858 -58177 -33242
rect -57473 -33858 -57177 -33242
rect -56473 -33858 -56177 -33242
rect -55473 -33858 -55177 -33242
rect -54473 -33858 -54177 -33242
rect -53473 -33858 -53177 -33242
rect -52473 -33858 -52177 -33242
rect -51473 -33858 -51177 -33242
rect -50473 -33858 -50177 -33242
rect -49473 -33858 -49177 -33242
rect -74813 -34198 -74517 -33902
rect -74473 -33928 -74177 -33902
rect -74473 -34172 -74447 -33928
rect -74447 -34172 -74203 -33928
rect -74203 -34172 -74177 -33928
rect -74473 -34198 -74177 -34172
rect -74133 -34198 -73517 -33902
rect -73473 -33928 -73177 -33902
rect -73473 -34172 -73447 -33928
rect -73447 -34172 -73203 -33928
rect -73203 -34172 -73177 -33928
rect -73473 -34198 -73177 -34172
rect -73133 -34198 -72517 -33902
rect -72473 -33928 -72177 -33902
rect -72473 -34172 -72447 -33928
rect -72447 -34172 -72203 -33928
rect -72203 -34172 -72177 -33928
rect -72473 -34198 -72177 -34172
rect -72133 -34198 -71517 -33902
rect -71473 -33928 -71177 -33902
rect -71473 -34172 -71447 -33928
rect -71447 -34172 -71203 -33928
rect -71203 -34172 -71177 -33928
rect -71473 -34198 -71177 -34172
rect -71133 -34198 -70517 -33902
rect -70473 -33928 -70177 -33902
rect -70473 -34172 -70447 -33928
rect -70447 -34172 -70203 -33928
rect -70203 -34172 -70177 -33928
rect -70473 -34198 -70177 -34172
rect -70133 -34198 -69517 -33902
rect -69473 -33928 -69177 -33902
rect -69473 -34172 -69447 -33928
rect -69447 -34172 -69203 -33928
rect -69203 -34172 -69177 -33928
rect -69473 -34198 -69177 -34172
rect -69133 -34198 -68517 -33902
rect -68473 -33928 -68177 -33902
rect -68473 -34172 -68447 -33928
rect -68447 -34172 -68203 -33928
rect -68203 -34172 -68177 -33928
rect -68473 -34198 -68177 -34172
rect -68133 -34198 -67517 -33902
rect -67473 -33928 -67177 -33902
rect -67473 -34172 -67447 -33928
rect -67447 -34172 -67203 -33928
rect -67203 -34172 -67177 -33928
rect -67473 -34198 -67177 -34172
rect -67133 -34198 -66517 -33902
rect -66473 -33928 -66177 -33902
rect -66473 -34172 -66447 -33928
rect -66447 -34172 -66203 -33928
rect -66203 -34172 -66177 -33928
rect -66473 -34198 -66177 -34172
rect -66133 -34198 -65517 -33902
rect -65473 -33928 -65177 -33902
rect -65473 -34172 -65447 -33928
rect -65447 -34172 -65203 -33928
rect -65203 -34172 -65177 -33928
rect -65473 -34198 -65177 -34172
rect -65133 -34198 -64517 -33902
rect -64473 -33928 -64177 -33902
rect -64473 -34172 -64447 -33928
rect -64447 -34172 -64203 -33928
rect -64203 -34172 -64177 -33928
rect -64473 -34198 -64177 -34172
rect -64133 -34198 -63517 -33902
rect -63473 -33928 -63177 -33902
rect -63473 -34172 -63447 -33928
rect -63447 -34172 -63203 -33928
rect -63203 -34172 -63177 -33928
rect -63473 -34198 -63177 -34172
rect -63133 -34198 -62517 -33902
rect -62473 -33928 -62177 -33902
rect -62473 -34172 -62447 -33928
rect -62447 -34172 -62203 -33928
rect -62203 -34172 -62177 -33928
rect -62473 -34198 -62177 -34172
rect -62133 -34198 -61517 -33902
rect -61473 -33928 -61177 -33902
rect -61473 -34172 -61447 -33928
rect -61447 -34172 -61203 -33928
rect -61203 -34172 -61177 -33928
rect -61473 -34198 -61177 -34172
rect -61133 -34198 -60517 -33902
rect -60473 -33928 -60177 -33902
rect -60473 -34172 -60447 -33928
rect -60447 -34172 -60203 -33928
rect -60203 -34172 -60177 -33928
rect -60473 -34198 -60177 -34172
rect -60133 -34198 -59517 -33902
rect -59473 -33928 -59177 -33902
rect -59473 -34172 -59447 -33928
rect -59447 -34172 -59203 -33928
rect -59203 -34172 -59177 -33928
rect -59473 -34198 -59177 -34172
rect -59133 -34198 -58517 -33902
rect -58473 -33928 -58177 -33902
rect -58473 -34172 -58447 -33928
rect -58447 -34172 -58203 -33928
rect -58203 -34172 -58177 -33928
rect -58473 -34198 -58177 -34172
rect -58133 -34198 -57517 -33902
rect -57473 -33928 -57177 -33902
rect -57473 -34172 -57447 -33928
rect -57447 -34172 -57203 -33928
rect -57203 -34172 -57177 -33928
rect -57473 -34198 -57177 -34172
rect -57133 -34198 -56517 -33902
rect -56473 -33928 -56177 -33902
rect -56473 -34172 -56447 -33928
rect -56447 -34172 -56203 -33928
rect -56203 -34172 -56177 -33928
rect -56473 -34198 -56177 -34172
rect -56133 -34198 -55517 -33902
rect -55473 -33928 -55177 -33902
rect -55473 -34172 -55447 -33928
rect -55447 -34172 -55203 -33928
rect -55203 -34172 -55177 -33928
rect -55473 -34198 -55177 -34172
rect -55133 -34198 -54517 -33902
rect -54473 -33928 -54177 -33902
rect -54473 -34172 -54447 -33928
rect -54447 -34172 -54203 -33928
rect -54203 -34172 -54177 -33928
rect -54473 -34198 -54177 -34172
rect -54133 -34198 -53517 -33902
rect -53473 -33928 -53177 -33902
rect -53473 -34172 -53447 -33928
rect -53447 -34172 -53203 -33928
rect -53203 -34172 -53177 -33928
rect -53473 -34198 -53177 -34172
rect -53133 -34198 -52517 -33902
rect -52473 -33928 -52177 -33902
rect -52473 -34172 -52447 -33928
rect -52447 -34172 -52203 -33928
rect -52203 -34172 -52177 -33928
rect -52473 -34198 -52177 -34172
rect -52133 -34198 -51517 -33902
rect -51473 -33928 -51177 -33902
rect -51473 -34172 -51447 -33928
rect -51447 -34172 -51203 -33928
rect -51203 -34172 -51177 -33928
rect -51473 -34198 -51177 -34172
rect -51133 -34198 -50517 -33902
rect -50473 -33928 -50177 -33902
rect -50473 -34172 -50447 -33928
rect -50447 -34172 -50203 -33928
rect -50203 -34172 -50177 -33928
rect -50473 -34198 -50177 -34172
rect -50133 -34198 -49517 -33902
rect -49473 -33928 -49177 -33902
rect -49473 -34172 -49447 -33928
rect -49447 -34172 -49203 -33928
rect -49203 -34172 -49177 -33928
rect -49473 -34198 -49177 -34172
rect -49133 -34198 -48837 -33902
rect -74473 -34858 -74177 -34242
rect -73473 -34858 -73177 -34242
rect -72473 -34858 -72177 -34242
rect -71473 -34858 -71177 -34242
rect -70473 -34858 -70177 -34242
rect -69473 -34858 -69177 -34242
rect -68473 -34858 -68177 -34242
rect -67473 -34858 -67177 -34242
rect -66473 -34858 -66177 -34242
rect -65473 -34858 -65177 -34242
rect -64473 -34858 -64177 -34242
rect -63473 -34858 -63177 -34242
rect -62473 -34858 -62177 -34242
rect -61473 -34858 -61177 -34242
rect -60473 -34858 -60177 -34242
rect -59473 -34858 -59177 -34242
rect -58473 -34858 -58177 -34242
rect -57473 -34858 -57177 -34242
rect -56473 -34858 -56177 -34242
rect -55473 -34858 -55177 -34242
rect -54473 -34858 -54177 -34242
rect -53473 -34858 -53177 -34242
rect -52473 -34858 -52177 -34242
rect -51473 -34858 -51177 -34242
rect -50473 -34858 -50177 -34242
rect -49473 -34858 -49177 -34242
rect -74813 -35198 -74517 -34902
rect -74473 -34928 -74177 -34902
rect -74473 -35172 -74447 -34928
rect -74447 -35172 -74203 -34928
rect -74203 -35172 -74177 -34928
rect -74473 -35198 -74177 -35172
rect -74133 -35198 -73517 -34902
rect -73473 -34928 -73177 -34902
rect -73473 -35172 -73447 -34928
rect -73447 -35172 -73203 -34928
rect -73203 -35172 -73177 -34928
rect -73473 -35198 -73177 -35172
rect -73133 -35198 -72517 -34902
rect -72473 -34928 -72177 -34902
rect -72473 -35172 -72447 -34928
rect -72447 -35172 -72203 -34928
rect -72203 -35172 -72177 -34928
rect -72473 -35198 -72177 -35172
rect -72133 -35198 -71517 -34902
rect -71473 -34928 -71177 -34902
rect -71473 -35172 -71447 -34928
rect -71447 -35172 -71203 -34928
rect -71203 -35172 -71177 -34928
rect -71473 -35198 -71177 -35172
rect -71133 -35198 -70517 -34902
rect -70473 -34928 -70177 -34902
rect -70473 -35172 -70447 -34928
rect -70447 -35172 -70203 -34928
rect -70203 -35172 -70177 -34928
rect -70473 -35198 -70177 -35172
rect -70133 -35198 -69517 -34902
rect -69473 -34928 -69177 -34902
rect -69473 -35172 -69447 -34928
rect -69447 -35172 -69203 -34928
rect -69203 -35172 -69177 -34928
rect -69473 -35198 -69177 -35172
rect -69133 -35198 -68517 -34902
rect -68473 -34928 -68177 -34902
rect -68473 -35172 -68447 -34928
rect -68447 -35172 -68203 -34928
rect -68203 -35172 -68177 -34928
rect -68473 -35198 -68177 -35172
rect -68133 -35198 -67517 -34902
rect -67473 -34928 -67177 -34902
rect -67473 -35172 -67447 -34928
rect -67447 -35172 -67203 -34928
rect -67203 -35172 -67177 -34928
rect -67473 -35198 -67177 -35172
rect -67133 -35198 -66517 -34902
rect -66473 -34928 -66177 -34902
rect -66473 -35172 -66447 -34928
rect -66447 -35172 -66203 -34928
rect -66203 -35172 -66177 -34928
rect -66473 -35198 -66177 -35172
rect -66133 -35198 -65517 -34902
rect -65473 -34928 -65177 -34902
rect -65473 -35172 -65447 -34928
rect -65447 -35172 -65203 -34928
rect -65203 -35172 -65177 -34928
rect -65473 -35198 -65177 -35172
rect -65133 -35198 -64517 -34902
rect -64473 -34928 -64177 -34902
rect -64473 -35172 -64447 -34928
rect -64447 -35172 -64203 -34928
rect -64203 -35172 -64177 -34928
rect -64473 -35198 -64177 -35172
rect -64133 -35198 -63517 -34902
rect -63473 -34928 -63177 -34902
rect -63473 -35172 -63447 -34928
rect -63447 -35172 -63203 -34928
rect -63203 -35172 -63177 -34928
rect -63473 -35198 -63177 -35172
rect -63133 -35198 -62517 -34902
rect -62473 -34928 -62177 -34902
rect -62473 -35172 -62447 -34928
rect -62447 -35172 -62203 -34928
rect -62203 -35172 -62177 -34928
rect -62473 -35198 -62177 -35172
rect -62133 -35198 -61517 -34902
rect -61473 -34928 -61177 -34902
rect -61473 -35172 -61447 -34928
rect -61447 -35172 -61203 -34928
rect -61203 -35172 -61177 -34928
rect -61473 -35198 -61177 -35172
rect -61133 -35198 -60517 -34902
rect -60473 -34928 -60177 -34902
rect -60473 -35172 -60447 -34928
rect -60447 -35172 -60203 -34928
rect -60203 -35172 -60177 -34928
rect -60473 -35198 -60177 -35172
rect -60133 -35198 -59517 -34902
rect -59473 -34928 -59177 -34902
rect -59473 -35172 -59447 -34928
rect -59447 -35172 -59203 -34928
rect -59203 -35172 -59177 -34928
rect -59473 -35198 -59177 -35172
rect -59133 -35198 -58517 -34902
rect -58473 -34928 -58177 -34902
rect -58473 -35172 -58447 -34928
rect -58447 -35172 -58203 -34928
rect -58203 -35172 -58177 -34928
rect -58473 -35198 -58177 -35172
rect -58133 -35198 -57517 -34902
rect -57473 -34928 -57177 -34902
rect -57473 -35172 -57447 -34928
rect -57447 -35172 -57203 -34928
rect -57203 -35172 -57177 -34928
rect -57473 -35198 -57177 -35172
rect -57133 -35198 -56517 -34902
rect -56473 -34928 -56177 -34902
rect -56473 -35172 -56447 -34928
rect -56447 -35172 -56203 -34928
rect -56203 -35172 -56177 -34928
rect -56473 -35198 -56177 -35172
rect -56133 -35198 -55517 -34902
rect -55473 -34928 -55177 -34902
rect -55473 -35172 -55447 -34928
rect -55447 -35172 -55203 -34928
rect -55203 -35172 -55177 -34928
rect -55473 -35198 -55177 -35172
rect -55133 -35198 -54517 -34902
rect -54473 -34928 -54177 -34902
rect -54473 -35172 -54447 -34928
rect -54447 -35172 -54203 -34928
rect -54203 -35172 -54177 -34928
rect -54473 -35198 -54177 -35172
rect -54133 -35198 -53517 -34902
rect -53473 -34928 -53177 -34902
rect -53473 -35172 -53447 -34928
rect -53447 -35172 -53203 -34928
rect -53203 -35172 -53177 -34928
rect -53473 -35198 -53177 -35172
rect -53133 -35198 -52517 -34902
rect -52473 -34928 -52177 -34902
rect -52473 -35172 -52447 -34928
rect -52447 -35172 -52203 -34928
rect -52203 -35172 -52177 -34928
rect -52473 -35198 -52177 -35172
rect -52133 -35198 -51517 -34902
rect -51473 -34928 -51177 -34902
rect -51473 -35172 -51447 -34928
rect -51447 -35172 -51203 -34928
rect -51203 -35172 -51177 -34928
rect -51473 -35198 -51177 -35172
rect -51133 -35198 -50517 -34902
rect -50473 -34928 -50177 -34902
rect -50473 -35172 -50447 -34928
rect -50447 -35172 -50203 -34928
rect -50203 -35172 -50177 -34928
rect -50473 -35198 -50177 -35172
rect -50133 -35198 -49517 -34902
rect -49473 -34928 -49177 -34902
rect -49473 -35172 -49447 -34928
rect -49447 -35172 -49203 -34928
rect -49203 -35172 -49177 -34928
rect -49473 -35198 -49177 -35172
rect -49133 -35198 -48837 -34902
rect -74473 -35858 -74177 -35242
rect -73473 -35858 -73177 -35242
rect -72473 -35858 -72177 -35242
rect -71473 -35858 -71177 -35242
rect -70473 -35858 -70177 -35242
rect -69473 -35858 -69177 -35242
rect -68473 -35858 -68177 -35242
rect -67473 -35858 -67177 -35242
rect -66473 -35858 -66177 -35242
rect -65473 -35858 -65177 -35242
rect -64473 -35858 -64177 -35242
rect -63473 -35858 -63177 -35242
rect -62473 -35858 -62177 -35242
rect -61473 -35858 -61177 -35242
rect -60473 -35858 -60177 -35242
rect -59473 -35858 -59177 -35242
rect -58473 -35858 -58177 -35242
rect -57473 -35858 -57177 -35242
rect -56473 -35858 -56177 -35242
rect -55473 -35858 -55177 -35242
rect -54473 -35858 -54177 -35242
rect -53473 -35858 -53177 -35242
rect -52473 -35858 -52177 -35242
rect -51473 -35858 -51177 -35242
rect -50473 -35858 -50177 -35242
rect -49473 -35858 -49177 -35242
rect -74813 -36198 -74517 -35902
rect -74473 -35928 -74177 -35902
rect -74473 -36172 -74447 -35928
rect -74447 -36172 -74203 -35928
rect -74203 -36172 -74177 -35928
rect -74473 -36198 -74177 -36172
rect -74133 -36198 -73517 -35902
rect -73473 -35928 -73177 -35902
rect -73473 -36172 -73447 -35928
rect -73447 -36172 -73203 -35928
rect -73203 -36172 -73177 -35928
rect -73473 -36198 -73177 -36172
rect -73133 -36198 -72517 -35902
rect -72473 -35928 -72177 -35902
rect -72473 -36172 -72447 -35928
rect -72447 -36172 -72203 -35928
rect -72203 -36172 -72177 -35928
rect -72473 -36198 -72177 -36172
rect -72133 -36198 -71517 -35902
rect -71473 -35928 -71177 -35902
rect -71473 -36172 -71447 -35928
rect -71447 -36172 -71203 -35928
rect -71203 -36172 -71177 -35928
rect -71473 -36198 -71177 -36172
rect -71133 -36198 -70517 -35902
rect -70473 -35928 -70177 -35902
rect -70473 -36172 -70447 -35928
rect -70447 -36172 -70203 -35928
rect -70203 -36172 -70177 -35928
rect -70473 -36198 -70177 -36172
rect -70133 -36198 -69517 -35902
rect -69473 -35928 -69177 -35902
rect -69473 -36172 -69447 -35928
rect -69447 -36172 -69203 -35928
rect -69203 -36172 -69177 -35928
rect -69473 -36198 -69177 -36172
rect -69133 -36198 -68517 -35902
rect -68473 -35928 -68177 -35902
rect -68473 -36172 -68447 -35928
rect -68447 -36172 -68203 -35928
rect -68203 -36172 -68177 -35928
rect -68473 -36198 -68177 -36172
rect -68133 -36198 -67517 -35902
rect -67473 -35928 -67177 -35902
rect -67473 -36172 -67447 -35928
rect -67447 -36172 -67203 -35928
rect -67203 -36172 -67177 -35928
rect -67473 -36198 -67177 -36172
rect -67133 -36198 -66517 -35902
rect -66473 -35928 -66177 -35902
rect -66473 -36172 -66447 -35928
rect -66447 -36172 -66203 -35928
rect -66203 -36172 -66177 -35928
rect -66473 -36198 -66177 -36172
rect -66133 -36198 -65517 -35902
rect -65473 -35928 -65177 -35902
rect -65473 -36172 -65447 -35928
rect -65447 -36172 -65203 -35928
rect -65203 -36172 -65177 -35928
rect -65473 -36198 -65177 -36172
rect -65133 -36198 -64517 -35902
rect -64473 -35928 -64177 -35902
rect -64473 -36172 -64447 -35928
rect -64447 -36172 -64203 -35928
rect -64203 -36172 -64177 -35928
rect -64473 -36198 -64177 -36172
rect -64133 -36198 -63517 -35902
rect -63473 -35928 -63177 -35902
rect -63473 -36172 -63447 -35928
rect -63447 -36172 -63203 -35928
rect -63203 -36172 -63177 -35928
rect -63473 -36198 -63177 -36172
rect -63133 -36198 -62517 -35902
rect -62473 -35928 -62177 -35902
rect -62473 -36172 -62447 -35928
rect -62447 -36172 -62203 -35928
rect -62203 -36172 -62177 -35928
rect -62473 -36198 -62177 -36172
rect -62133 -36198 -61517 -35902
rect -61473 -35928 -61177 -35902
rect -61473 -36172 -61447 -35928
rect -61447 -36172 -61203 -35928
rect -61203 -36172 -61177 -35928
rect -61473 -36198 -61177 -36172
rect -61133 -36198 -60517 -35902
rect -60473 -35928 -60177 -35902
rect -60473 -36172 -60447 -35928
rect -60447 -36172 -60203 -35928
rect -60203 -36172 -60177 -35928
rect -60473 -36198 -60177 -36172
rect -60133 -36198 -59517 -35902
rect -59473 -35928 -59177 -35902
rect -59473 -36172 -59447 -35928
rect -59447 -36172 -59203 -35928
rect -59203 -36172 -59177 -35928
rect -59473 -36198 -59177 -36172
rect -59133 -36198 -58517 -35902
rect -58473 -35928 -58177 -35902
rect -58473 -36172 -58447 -35928
rect -58447 -36172 -58203 -35928
rect -58203 -36172 -58177 -35928
rect -58473 -36198 -58177 -36172
rect -58133 -36198 -57517 -35902
rect -57473 -35928 -57177 -35902
rect -57473 -36172 -57447 -35928
rect -57447 -36172 -57203 -35928
rect -57203 -36172 -57177 -35928
rect -57473 -36198 -57177 -36172
rect -57133 -36198 -56517 -35902
rect -56473 -35928 -56177 -35902
rect -56473 -36172 -56447 -35928
rect -56447 -36172 -56203 -35928
rect -56203 -36172 -56177 -35928
rect -56473 -36198 -56177 -36172
rect -56133 -36198 -55517 -35902
rect -55473 -35928 -55177 -35902
rect -55473 -36172 -55447 -35928
rect -55447 -36172 -55203 -35928
rect -55203 -36172 -55177 -35928
rect -55473 -36198 -55177 -36172
rect -55133 -36198 -54517 -35902
rect -54473 -35928 -54177 -35902
rect -54473 -36172 -54447 -35928
rect -54447 -36172 -54203 -35928
rect -54203 -36172 -54177 -35928
rect -54473 -36198 -54177 -36172
rect -54133 -36198 -53517 -35902
rect -53473 -35928 -53177 -35902
rect -53473 -36172 -53447 -35928
rect -53447 -36172 -53203 -35928
rect -53203 -36172 -53177 -35928
rect -53473 -36198 -53177 -36172
rect -53133 -36198 -52517 -35902
rect -52473 -35928 -52177 -35902
rect -52473 -36172 -52447 -35928
rect -52447 -36172 -52203 -35928
rect -52203 -36172 -52177 -35928
rect -52473 -36198 -52177 -36172
rect -52133 -36198 -51517 -35902
rect -51473 -35928 -51177 -35902
rect -51473 -36172 -51447 -35928
rect -51447 -36172 -51203 -35928
rect -51203 -36172 -51177 -35928
rect -51473 -36198 -51177 -36172
rect -51133 -36198 -50517 -35902
rect -50473 -35928 -50177 -35902
rect -50473 -36172 -50447 -35928
rect -50447 -36172 -50203 -35928
rect -50203 -36172 -50177 -35928
rect -50473 -36198 -50177 -36172
rect -50133 -36198 -49517 -35902
rect -49473 -35928 -49177 -35902
rect -49473 -36172 -49447 -35928
rect -49447 -36172 -49203 -35928
rect -49203 -36172 -49177 -35928
rect -49473 -36198 -49177 -36172
rect -49133 -36198 -48837 -35902
rect -74473 -36858 -74177 -36242
rect -73473 -36858 -73177 -36242
rect -72473 -36858 -72177 -36242
rect -71473 -36858 -71177 -36242
rect -70473 -36858 -70177 -36242
rect -69473 -36858 -69177 -36242
rect -68473 -36858 -68177 -36242
rect -67473 -36858 -67177 -36242
rect -66473 -36858 -66177 -36242
rect -65473 -36858 -65177 -36242
rect -64473 -36858 -64177 -36242
rect -63473 -36858 -63177 -36242
rect -62473 -36858 -62177 -36242
rect -61473 -36858 -61177 -36242
rect -60473 -36858 -60177 -36242
rect -59473 -36858 -59177 -36242
rect -58473 -36858 -58177 -36242
rect -57473 -36858 -57177 -36242
rect -56473 -36858 -56177 -36242
rect -55473 -36858 -55177 -36242
rect -54473 -36858 -54177 -36242
rect -53473 -36858 -53177 -36242
rect -52473 -36858 -52177 -36242
rect -51473 -36858 -51177 -36242
rect -50473 -36858 -50177 -36242
rect -49473 -36858 -49177 -36242
rect -74813 -37198 -74517 -36902
rect -74473 -36928 -74177 -36902
rect -74473 -37172 -74447 -36928
rect -74447 -37172 -74203 -36928
rect -74203 -37172 -74177 -36928
rect -74473 -37198 -74177 -37172
rect -74133 -37198 -73517 -36902
rect -73473 -36928 -73177 -36902
rect -73473 -37172 -73447 -36928
rect -73447 -37172 -73203 -36928
rect -73203 -37172 -73177 -36928
rect -73473 -37198 -73177 -37172
rect -73133 -37198 -72517 -36902
rect -72473 -36928 -72177 -36902
rect -72473 -37172 -72447 -36928
rect -72447 -37172 -72203 -36928
rect -72203 -37172 -72177 -36928
rect -72473 -37198 -72177 -37172
rect -72133 -37198 -71517 -36902
rect -71473 -36928 -71177 -36902
rect -71473 -37172 -71447 -36928
rect -71447 -37172 -71203 -36928
rect -71203 -37172 -71177 -36928
rect -71473 -37198 -71177 -37172
rect -71133 -37198 -70517 -36902
rect -70473 -36928 -70177 -36902
rect -70473 -37172 -70447 -36928
rect -70447 -37172 -70203 -36928
rect -70203 -37172 -70177 -36928
rect -70473 -37198 -70177 -37172
rect -70133 -37198 -69517 -36902
rect -69473 -36928 -69177 -36902
rect -69473 -37172 -69447 -36928
rect -69447 -37172 -69203 -36928
rect -69203 -37172 -69177 -36928
rect -69473 -37198 -69177 -37172
rect -69133 -37198 -68517 -36902
rect -68473 -36928 -68177 -36902
rect -68473 -37172 -68447 -36928
rect -68447 -37172 -68203 -36928
rect -68203 -37172 -68177 -36928
rect -68473 -37198 -68177 -37172
rect -68133 -37198 -67517 -36902
rect -67473 -36928 -67177 -36902
rect -67473 -37172 -67447 -36928
rect -67447 -37172 -67203 -36928
rect -67203 -37172 -67177 -36928
rect -67473 -37198 -67177 -37172
rect -67133 -37198 -66517 -36902
rect -66473 -36928 -66177 -36902
rect -66473 -37172 -66447 -36928
rect -66447 -37172 -66203 -36928
rect -66203 -37172 -66177 -36928
rect -66473 -37198 -66177 -37172
rect -66133 -37198 -65517 -36902
rect -65473 -36928 -65177 -36902
rect -65473 -37172 -65447 -36928
rect -65447 -37172 -65203 -36928
rect -65203 -37172 -65177 -36928
rect -65473 -37198 -65177 -37172
rect -65133 -37198 -64517 -36902
rect -64473 -36928 -64177 -36902
rect -64473 -37172 -64447 -36928
rect -64447 -37172 -64203 -36928
rect -64203 -37172 -64177 -36928
rect -64473 -37198 -64177 -37172
rect -64133 -37198 -63517 -36902
rect -63473 -36928 -63177 -36902
rect -63473 -37172 -63447 -36928
rect -63447 -37172 -63203 -36928
rect -63203 -37172 -63177 -36928
rect -63473 -37198 -63177 -37172
rect -63133 -37198 -62517 -36902
rect -62473 -36928 -62177 -36902
rect -62473 -37172 -62447 -36928
rect -62447 -37172 -62203 -36928
rect -62203 -37172 -62177 -36928
rect -62473 -37198 -62177 -37172
rect -62133 -37198 -61517 -36902
rect -61473 -36928 -61177 -36902
rect -61473 -37172 -61447 -36928
rect -61447 -37172 -61203 -36928
rect -61203 -37172 -61177 -36928
rect -61473 -37198 -61177 -37172
rect -61133 -37198 -60517 -36902
rect -60473 -36928 -60177 -36902
rect -60473 -37172 -60447 -36928
rect -60447 -37172 -60203 -36928
rect -60203 -37172 -60177 -36928
rect -60473 -37198 -60177 -37172
rect -60133 -37198 -59517 -36902
rect -59473 -36928 -59177 -36902
rect -59473 -37172 -59447 -36928
rect -59447 -37172 -59203 -36928
rect -59203 -37172 -59177 -36928
rect -59473 -37198 -59177 -37172
rect -59133 -37198 -58517 -36902
rect -58473 -36928 -58177 -36902
rect -58473 -37172 -58447 -36928
rect -58447 -37172 -58203 -36928
rect -58203 -37172 -58177 -36928
rect -58473 -37198 -58177 -37172
rect -58133 -37198 -57517 -36902
rect -57473 -36928 -57177 -36902
rect -57473 -37172 -57447 -36928
rect -57447 -37172 -57203 -36928
rect -57203 -37172 -57177 -36928
rect -57473 -37198 -57177 -37172
rect -57133 -37198 -56517 -36902
rect -56473 -36928 -56177 -36902
rect -56473 -37172 -56447 -36928
rect -56447 -37172 -56203 -36928
rect -56203 -37172 -56177 -36928
rect -56473 -37198 -56177 -37172
rect -56133 -37198 -55517 -36902
rect -55473 -36928 -55177 -36902
rect -55473 -37172 -55447 -36928
rect -55447 -37172 -55203 -36928
rect -55203 -37172 -55177 -36928
rect -55473 -37198 -55177 -37172
rect -55133 -37198 -54517 -36902
rect -54473 -36928 -54177 -36902
rect -54473 -37172 -54447 -36928
rect -54447 -37172 -54203 -36928
rect -54203 -37172 -54177 -36928
rect -54473 -37198 -54177 -37172
rect -54133 -37198 -53517 -36902
rect -53473 -36928 -53177 -36902
rect -53473 -37172 -53447 -36928
rect -53447 -37172 -53203 -36928
rect -53203 -37172 -53177 -36928
rect -53473 -37198 -53177 -37172
rect -53133 -37198 -52517 -36902
rect -52473 -36928 -52177 -36902
rect -52473 -37172 -52447 -36928
rect -52447 -37172 -52203 -36928
rect -52203 -37172 -52177 -36928
rect -52473 -37198 -52177 -37172
rect -52133 -37198 -51517 -36902
rect -51473 -36928 -51177 -36902
rect -51473 -37172 -51447 -36928
rect -51447 -37172 -51203 -36928
rect -51203 -37172 -51177 -36928
rect -51473 -37198 -51177 -37172
rect -51133 -37198 -50517 -36902
rect -50473 -36928 -50177 -36902
rect -50473 -37172 -50447 -36928
rect -50447 -37172 -50203 -36928
rect -50203 -37172 -50177 -36928
rect -50473 -37198 -50177 -37172
rect -50133 -37198 -49517 -36902
rect -49473 -36928 -49177 -36902
rect -49473 -37172 -49447 -36928
rect -49447 -37172 -49203 -36928
rect -49203 -37172 -49177 -36928
rect -49473 -37198 -49177 -37172
rect -49133 -37198 -48837 -36902
rect -74473 -37858 -74177 -37242
rect -73473 -37858 -73177 -37242
rect -72473 -37858 -72177 -37242
rect -71473 -37858 -71177 -37242
rect -70473 -37858 -70177 -37242
rect -69473 -37858 -69177 -37242
rect -68473 -37858 -68177 -37242
rect -67473 -37858 -67177 -37242
rect -66473 -37858 -66177 -37242
rect -65473 -37858 -65177 -37242
rect -64473 -37858 -64177 -37242
rect -63473 -37858 -63177 -37242
rect -62473 -37858 -62177 -37242
rect -61473 -37858 -61177 -37242
rect -60473 -37858 -60177 -37242
rect -59473 -37858 -59177 -37242
rect -58473 -37858 -58177 -37242
rect -57473 -37858 -57177 -37242
rect -56473 -37858 -56177 -37242
rect -55473 -37858 -55177 -37242
rect -54473 -37858 -54177 -37242
rect -53473 -37858 -53177 -37242
rect -52473 -37858 -52177 -37242
rect -51473 -37858 -51177 -37242
rect -50473 -37858 -50177 -37242
rect -49473 -37858 -49177 -37242
rect -74813 -38198 -74517 -37902
rect -74473 -37928 -74177 -37902
rect -74473 -38172 -74447 -37928
rect -74447 -38172 -74203 -37928
rect -74203 -38172 -74177 -37928
rect -74473 -38198 -74177 -38172
rect -74133 -38198 -73517 -37902
rect -73473 -37928 -73177 -37902
rect -73473 -38172 -73447 -37928
rect -73447 -38172 -73203 -37928
rect -73203 -38172 -73177 -37928
rect -73473 -38198 -73177 -38172
rect -73133 -38198 -72517 -37902
rect -72473 -37928 -72177 -37902
rect -72473 -38172 -72447 -37928
rect -72447 -38172 -72203 -37928
rect -72203 -38172 -72177 -37928
rect -72473 -38198 -72177 -38172
rect -72133 -38198 -71517 -37902
rect -71473 -37928 -71177 -37902
rect -71473 -38172 -71447 -37928
rect -71447 -38172 -71203 -37928
rect -71203 -38172 -71177 -37928
rect -71473 -38198 -71177 -38172
rect -71133 -38198 -70517 -37902
rect -70473 -37928 -70177 -37902
rect -70473 -38172 -70447 -37928
rect -70447 -38172 -70203 -37928
rect -70203 -38172 -70177 -37928
rect -70473 -38198 -70177 -38172
rect -70133 -38198 -69517 -37902
rect -69473 -37928 -69177 -37902
rect -69473 -38172 -69447 -37928
rect -69447 -38172 -69203 -37928
rect -69203 -38172 -69177 -37928
rect -69473 -38198 -69177 -38172
rect -69133 -38198 -68517 -37902
rect -68473 -37928 -68177 -37902
rect -68473 -38172 -68447 -37928
rect -68447 -38172 -68203 -37928
rect -68203 -38172 -68177 -37928
rect -68473 -38198 -68177 -38172
rect -68133 -38198 -67517 -37902
rect -67473 -37928 -67177 -37902
rect -67473 -38172 -67447 -37928
rect -67447 -38172 -67203 -37928
rect -67203 -38172 -67177 -37928
rect -67473 -38198 -67177 -38172
rect -67133 -38198 -66517 -37902
rect -66473 -37928 -66177 -37902
rect -66473 -38172 -66447 -37928
rect -66447 -38172 -66203 -37928
rect -66203 -38172 -66177 -37928
rect -66473 -38198 -66177 -38172
rect -66133 -38198 -65517 -37902
rect -65473 -37928 -65177 -37902
rect -65473 -38172 -65447 -37928
rect -65447 -38172 -65203 -37928
rect -65203 -38172 -65177 -37928
rect -65473 -38198 -65177 -38172
rect -65133 -38198 -64517 -37902
rect -64473 -37928 -64177 -37902
rect -64473 -38172 -64447 -37928
rect -64447 -38172 -64203 -37928
rect -64203 -38172 -64177 -37928
rect -64473 -38198 -64177 -38172
rect -64133 -38198 -63517 -37902
rect -63473 -37928 -63177 -37902
rect -63473 -38172 -63447 -37928
rect -63447 -38172 -63203 -37928
rect -63203 -38172 -63177 -37928
rect -63473 -38198 -63177 -38172
rect -63133 -38198 -62517 -37902
rect -62473 -37928 -62177 -37902
rect -62473 -38172 -62447 -37928
rect -62447 -38172 -62203 -37928
rect -62203 -38172 -62177 -37928
rect -62473 -38198 -62177 -38172
rect -62133 -38198 -61517 -37902
rect -61473 -37928 -61177 -37902
rect -61473 -38172 -61447 -37928
rect -61447 -38172 -61203 -37928
rect -61203 -38172 -61177 -37928
rect -61473 -38198 -61177 -38172
rect -61133 -38198 -60517 -37902
rect -60473 -37928 -60177 -37902
rect -60473 -38172 -60447 -37928
rect -60447 -38172 -60203 -37928
rect -60203 -38172 -60177 -37928
rect -60473 -38198 -60177 -38172
rect -60133 -38198 -59517 -37902
rect -59473 -37928 -59177 -37902
rect -59473 -38172 -59447 -37928
rect -59447 -38172 -59203 -37928
rect -59203 -38172 -59177 -37928
rect -59473 -38198 -59177 -38172
rect -59133 -38198 -58517 -37902
rect -58473 -37928 -58177 -37902
rect -58473 -38172 -58447 -37928
rect -58447 -38172 -58203 -37928
rect -58203 -38172 -58177 -37928
rect -58473 -38198 -58177 -38172
rect -58133 -38198 -57517 -37902
rect -57473 -37928 -57177 -37902
rect -57473 -38172 -57447 -37928
rect -57447 -38172 -57203 -37928
rect -57203 -38172 -57177 -37928
rect -57473 -38198 -57177 -38172
rect -57133 -38198 -56517 -37902
rect -56473 -37928 -56177 -37902
rect -56473 -38172 -56447 -37928
rect -56447 -38172 -56203 -37928
rect -56203 -38172 -56177 -37928
rect -56473 -38198 -56177 -38172
rect -56133 -38198 -55517 -37902
rect -55473 -37928 -55177 -37902
rect -55473 -38172 -55447 -37928
rect -55447 -38172 -55203 -37928
rect -55203 -38172 -55177 -37928
rect -55473 -38198 -55177 -38172
rect -55133 -38198 -54517 -37902
rect -54473 -37928 -54177 -37902
rect -54473 -38172 -54447 -37928
rect -54447 -38172 -54203 -37928
rect -54203 -38172 -54177 -37928
rect -54473 -38198 -54177 -38172
rect -54133 -38198 -53517 -37902
rect -53473 -37928 -53177 -37902
rect -53473 -38172 -53447 -37928
rect -53447 -38172 -53203 -37928
rect -53203 -38172 -53177 -37928
rect -53473 -38198 -53177 -38172
rect -53133 -38198 -52517 -37902
rect -52473 -37928 -52177 -37902
rect -52473 -38172 -52447 -37928
rect -52447 -38172 -52203 -37928
rect -52203 -38172 -52177 -37928
rect -52473 -38198 -52177 -38172
rect -52133 -38198 -51517 -37902
rect -51473 -37928 -51177 -37902
rect -51473 -38172 -51447 -37928
rect -51447 -38172 -51203 -37928
rect -51203 -38172 -51177 -37928
rect -51473 -38198 -51177 -38172
rect -51133 -38198 -50517 -37902
rect -50473 -37928 -50177 -37902
rect -50473 -38172 -50447 -37928
rect -50447 -38172 -50203 -37928
rect -50203 -38172 -50177 -37928
rect -50473 -38198 -50177 -38172
rect -50133 -38198 -49517 -37902
rect -49473 -37928 -49177 -37902
rect -49473 -38172 -49447 -37928
rect -49447 -38172 -49203 -37928
rect -49203 -38172 -49177 -37928
rect -49473 -38198 -49177 -38172
rect -49133 -38198 -48837 -37902
rect -74473 -38858 -74177 -38242
rect -73473 -38858 -73177 -38242
rect -72473 -38858 -72177 -38242
rect -71473 -38858 -71177 -38242
rect -70473 -38858 -70177 -38242
rect -69473 -38858 -69177 -38242
rect -68473 -38858 -68177 -38242
rect -67473 -38858 -67177 -38242
rect -66473 -38858 -66177 -38242
rect -65473 -38858 -65177 -38242
rect -64473 -38858 -64177 -38242
rect -63473 -38858 -63177 -38242
rect -62473 -38858 -62177 -38242
rect -61473 -38858 -61177 -38242
rect -60473 -38858 -60177 -38242
rect -59473 -38858 -59177 -38242
rect -58473 -38858 -58177 -38242
rect -57473 -38858 -57177 -38242
rect -56473 -38858 -56177 -38242
rect -55473 -38858 -55177 -38242
rect -54473 -38858 -54177 -38242
rect -53473 -38858 -53177 -38242
rect -52473 -38858 -52177 -38242
rect -51473 -38858 -51177 -38242
rect -50473 -38858 -50177 -38242
rect -49473 -38858 -49177 -38242
rect -74813 -39198 -74517 -38902
rect -74473 -38928 -74177 -38902
rect -74473 -39172 -74447 -38928
rect -74447 -39172 -74203 -38928
rect -74203 -39172 -74177 -38928
rect -74473 -39198 -74177 -39172
rect -74133 -39198 -73517 -38902
rect -73473 -38928 -73177 -38902
rect -73473 -39172 -73447 -38928
rect -73447 -39172 -73203 -38928
rect -73203 -39172 -73177 -38928
rect -73473 -39198 -73177 -39172
rect -73133 -39198 -72517 -38902
rect -72473 -38928 -72177 -38902
rect -72473 -39172 -72447 -38928
rect -72447 -39172 -72203 -38928
rect -72203 -39172 -72177 -38928
rect -72473 -39198 -72177 -39172
rect -72133 -39198 -71517 -38902
rect -71473 -38928 -71177 -38902
rect -71473 -39172 -71447 -38928
rect -71447 -39172 -71203 -38928
rect -71203 -39172 -71177 -38928
rect -71473 -39198 -71177 -39172
rect -71133 -39198 -70517 -38902
rect -70473 -38928 -70177 -38902
rect -70473 -39172 -70447 -38928
rect -70447 -39172 -70203 -38928
rect -70203 -39172 -70177 -38928
rect -70473 -39198 -70177 -39172
rect -70133 -39198 -69517 -38902
rect -69473 -38928 -69177 -38902
rect -69473 -39172 -69447 -38928
rect -69447 -39172 -69203 -38928
rect -69203 -39172 -69177 -38928
rect -69473 -39198 -69177 -39172
rect -69133 -39198 -68517 -38902
rect -68473 -38928 -68177 -38902
rect -68473 -39172 -68447 -38928
rect -68447 -39172 -68203 -38928
rect -68203 -39172 -68177 -38928
rect -68473 -39198 -68177 -39172
rect -68133 -39198 -67517 -38902
rect -67473 -38928 -67177 -38902
rect -67473 -39172 -67447 -38928
rect -67447 -39172 -67203 -38928
rect -67203 -39172 -67177 -38928
rect -67473 -39198 -67177 -39172
rect -67133 -39198 -66517 -38902
rect -66473 -38928 -66177 -38902
rect -66473 -39172 -66447 -38928
rect -66447 -39172 -66203 -38928
rect -66203 -39172 -66177 -38928
rect -66473 -39198 -66177 -39172
rect -66133 -39198 -65517 -38902
rect -65473 -38928 -65177 -38902
rect -65473 -39172 -65447 -38928
rect -65447 -39172 -65203 -38928
rect -65203 -39172 -65177 -38928
rect -65473 -39198 -65177 -39172
rect -65133 -39198 -64517 -38902
rect -64473 -38928 -64177 -38902
rect -64473 -39172 -64447 -38928
rect -64447 -39172 -64203 -38928
rect -64203 -39172 -64177 -38928
rect -64473 -39198 -64177 -39172
rect -64133 -39198 -63517 -38902
rect -63473 -38928 -63177 -38902
rect -63473 -39172 -63447 -38928
rect -63447 -39172 -63203 -38928
rect -63203 -39172 -63177 -38928
rect -63473 -39198 -63177 -39172
rect -63133 -39198 -62517 -38902
rect -62473 -38928 -62177 -38902
rect -62473 -39172 -62447 -38928
rect -62447 -39172 -62203 -38928
rect -62203 -39172 -62177 -38928
rect -62473 -39198 -62177 -39172
rect -62133 -39198 -61517 -38902
rect -61473 -38928 -61177 -38902
rect -61473 -39172 -61447 -38928
rect -61447 -39172 -61203 -38928
rect -61203 -39172 -61177 -38928
rect -61473 -39198 -61177 -39172
rect -61133 -39198 -60517 -38902
rect -60473 -38928 -60177 -38902
rect -60473 -39172 -60447 -38928
rect -60447 -39172 -60203 -38928
rect -60203 -39172 -60177 -38928
rect -60473 -39198 -60177 -39172
rect -60133 -39198 -59517 -38902
rect -59473 -38928 -59177 -38902
rect -59473 -39172 -59447 -38928
rect -59447 -39172 -59203 -38928
rect -59203 -39172 -59177 -38928
rect -59473 -39198 -59177 -39172
rect -59133 -39198 -58517 -38902
rect -58473 -38928 -58177 -38902
rect -58473 -39172 -58447 -38928
rect -58447 -39172 -58203 -38928
rect -58203 -39172 -58177 -38928
rect -58473 -39198 -58177 -39172
rect -58133 -39198 -57517 -38902
rect -57473 -38928 -57177 -38902
rect -57473 -39172 -57447 -38928
rect -57447 -39172 -57203 -38928
rect -57203 -39172 -57177 -38928
rect -57473 -39198 -57177 -39172
rect -57133 -39198 -56517 -38902
rect -56473 -38928 -56177 -38902
rect -56473 -39172 -56447 -38928
rect -56447 -39172 -56203 -38928
rect -56203 -39172 -56177 -38928
rect -56473 -39198 -56177 -39172
rect -56133 -39198 -55517 -38902
rect -55473 -38928 -55177 -38902
rect -55473 -39172 -55447 -38928
rect -55447 -39172 -55203 -38928
rect -55203 -39172 -55177 -38928
rect -55473 -39198 -55177 -39172
rect -55133 -39198 -54517 -38902
rect -54473 -38928 -54177 -38902
rect -54473 -39172 -54447 -38928
rect -54447 -39172 -54203 -38928
rect -54203 -39172 -54177 -38928
rect -54473 -39198 -54177 -39172
rect -54133 -39198 -53517 -38902
rect -53473 -38928 -53177 -38902
rect -53473 -39172 -53447 -38928
rect -53447 -39172 -53203 -38928
rect -53203 -39172 -53177 -38928
rect -53473 -39198 -53177 -39172
rect -53133 -39198 -52517 -38902
rect -52473 -38928 -52177 -38902
rect -52473 -39172 -52447 -38928
rect -52447 -39172 -52203 -38928
rect -52203 -39172 -52177 -38928
rect -52473 -39198 -52177 -39172
rect -52133 -39198 -51517 -38902
rect -51473 -38928 -51177 -38902
rect -51473 -39172 -51447 -38928
rect -51447 -39172 -51203 -38928
rect -51203 -39172 -51177 -38928
rect -51473 -39198 -51177 -39172
rect -51133 -39198 -50517 -38902
rect -50473 -38928 -50177 -38902
rect -50473 -39172 -50447 -38928
rect -50447 -39172 -50203 -38928
rect -50203 -39172 -50177 -38928
rect -50473 -39198 -50177 -39172
rect -50133 -39198 -49517 -38902
rect -49473 -38928 -49177 -38902
rect -49473 -39172 -49447 -38928
rect -49447 -39172 -49203 -38928
rect -49203 -39172 -49177 -38928
rect -49473 -39198 -49177 -39172
rect -49133 -39198 -48837 -38902
rect -74473 -39858 -74177 -39242
rect -73473 -39858 -73177 -39242
rect -72473 -39858 -72177 -39242
rect -71473 -39858 -71177 -39242
rect -70473 -39858 -70177 -39242
rect -69473 -39858 -69177 -39242
rect -68473 -39858 -68177 -39242
rect -67473 -39858 -67177 -39242
rect -66473 -39858 -66177 -39242
rect -65473 -39858 -65177 -39242
rect -64473 -39858 -64177 -39242
rect -63473 -39858 -63177 -39242
rect -62473 -39858 -62177 -39242
rect -61473 -39858 -61177 -39242
rect -60473 -39858 -60177 -39242
rect -59473 -39858 -59177 -39242
rect -58473 -39858 -58177 -39242
rect -57473 -39858 -57177 -39242
rect -56473 -39858 -56177 -39242
rect -55473 -39858 -55177 -39242
rect -54473 -39858 -54177 -39242
rect -53473 -39858 -53177 -39242
rect -52473 -39858 -52177 -39242
rect -51473 -39858 -51177 -39242
rect -50473 -39858 -50177 -39242
rect -49473 -39858 -49177 -39242
rect -74813 -40198 -74517 -39902
rect -74473 -39928 -74177 -39902
rect -74473 -40172 -74447 -39928
rect -74447 -40172 -74203 -39928
rect -74203 -40172 -74177 -39928
rect -74473 -40198 -74177 -40172
rect -74133 -40198 -73517 -39902
rect -73473 -39928 -73177 -39902
rect -73473 -40172 -73447 -39928
rect -73447 -40172 -73203 -39928
rect -73203 -40172 -73177 -39928
rect -73473 -40198 -73177 -40172
rect -73133 -40198 -72517 -39902
rect -72473 -39928 -72177 -39902
rect -72473 -40172 -72447 -39928
rect -72447 -40172 -72203 -39928
rect -72203 -40172 -72177 -39928
rect -72473 -40198 -72177 -40172
rect -72133 -40198 -71517 -39902
rect -71473 -39928 -71177 -39902
rect -71473 -40172 -71447 -39928
rect -71447 -40172 -71203 -39928
rect -71203 -40172 -71177 -39928
rect -71473 -40198 -71177 -40172
rect -71133 -40198 -70517 -39902
rect -70473 -39928 -70177 -39902
rect -70473 -40172 -70447 -39928
rect -70447 -40172 -70203 -39928
rect -70203 -40172 -70177 -39928
rect -70473 -40198 -70177 -40172
rect -70133 -40198 -69517 -39902
rect -69473 -39928 -69177 -39902
rect -69473 -40172 -69447 -39928
rect -69447 -40172 -69203 -39928
rect -69203 -40172 -69177 -39928
rect -69473 -40198 -69177 -40172
rect -69133 -40198 -68517 -39902
rect -68473 -39928 -68177 -39902
rect -68473 -40172 -68447 -39928
rect -68447 -40172 -68203 -39928
rect -68203 -40172 -68177 -39928
rect -68473 -40198 -68177 -40172
rect -68133 -40198 -67517 -39902
rect -67473 -39928 -67177 -39902
rect -67473 -40172 -67447 -39928
rect -67447 -40172 -67203 -39928
rect -67203 -40172 -67177 -39928
rect -67473 -40198 -67177 -40172
rect -67133 -40198 -66517 -39902
rect -66473 -39928 -66177 -39902
rect -66473 -40172 -66447 -39928
rect -66447 -40172 -66203 -39928
rect -66203 -40172 -66177 -39928
rect -66473 -40198 -66177 -40172
rect -66133 -40198 -65517 -39902
rect -65473 -39928 -65177 -39902
rect -65473 -40172 -65447 -39928
rect -65447 -40172 -65203 -39928
rect -65203 -40172 -65177 -39928
rect -65473 -40198 -65177 -40172
rect -65133 -40198 -64517 -39902
rect -64473 -39928 -64177 -39902
rect -64473 -40172 -64447 -39928
rect -64447 -40172 -64203 -39928
rect -64203 -40172 -64177 -39928
rect -64473 -40198 -64177 -40172
rect -64133 -40198 -63517 -39902
rect -63473 -39928 -63177 -39902
rect -63473 -40172 -63447 -39928
rect -63447 -40172 -63203 -39928
rect -63203 -40172 -63177 -39928
rect -63473 -40198 -63177 -40172
rect -63133 -40198 -62517 -39902
rect -62473 -39928 -62177 -39902
rect -62473 -40172 -62447 -39928
rect -62447 -40172 -62203 -39928
rect -62203 -40172 -62177 -39928
rect -62473 -40198 -62177 -40172
rect -62133 -40198 -61517 -39902
rect -61473 -39928 -61177 -39902
rect -61473 -40172 -61447 -39928
rect -61447 -40172 -61203 -39928
rect -61203 -40172 -61177 -39928
rect -61473 -40198 -61177 -40172
rect -61133 -40198 -60517 -39902
rect -60473 -39928 -60177 -39902
rect -60473 -40172 -60447 -39928
rect -60447 -40172 -60203 -39928
rect -60203 -40172 -60177 -39928
rect -60473 -40198 -60177 -40172
rect -60133 -40198 -59517 -39902
rect -59473 -39928 -59177 -39902
rect -59473 -40172 -59447 -39928
rect -59447 -40172 -59203 -39928
rect -59203 -40172 -59177 -39928
rect -59473 -40198 -59177 -40172
rect -59133 -40198 -58517 -39902
rect -58473 -39928 -58177 -39902
rect -58473 -40172 -58447 -39928
rect -58447 -40172 -58203 -39928
rect -58203 -40172 -58177 -39928
rect -58473 -40198 -58177 -40172
rect -58133 -40198 -57517 -39902
rect -57473 -39928 -57177 -39902
rect -57473 -40172 -57447 -39928
rect -57447 -40172 -57203 -39928
rect -57203 -40172 -57177 -39928
rect -57473 -40198 -57177 -40172
rect -57133 -40198 -56517 -39902
rect -56473 -39928 -56177 -39902
rect -56473 -40172 -56447 -39928
rect -56447 -40172 -56203 -39928
rect -56203 -40172 -56177 -39928
rect -56473 -40198 -56177 -40172
rect -56133 -40198 -55517 -39902
rect -55473 -39928 -55177 -39902
rect -55473 -40172 -55447 -39928
rect -55447 -40172 -55203 -39928
rect -55203 -40172 -55177 -39928
rect -55473 -40198 -55177 -40172
rect -55133 -40198 -54517 -39902
rect -54473 -39928 -54177 -39902
rect -54473 -40172 -54447 -39928
rect -54447 -40172 -54203 -39928
rect -54203 -40172 -54177 -39928
rect -54473 -40198 -54177 -40172
rect -54133 -40198 -53517 -39902
rect -53473 -39928 -53177 -39902
rect -53473 -40172 -53447 -39928
rect -53447 -40172 -53203 -39928
rect -53203 -40172 -53177 -39928
rect -53473 -40198 -53177 -40172
rect -53133 -40198 -52517 -39902
rect -52473 -39928 -52177 -39902
rect -52473 -40172 -52447 -39928
rect -52447 -40172 -52203 -39928
rect -52203 -40172 -52177 -39928
rect -52473 -40198 -52177 -40172
rect -52133 -40198 -51517 -39902
rect -51473 -39928 -51177 -39902
rect -51473 -40172 -51447 -39928
rect -51447 -40172 -51203 -39928
rect -51203 -40172 -51177 -39928
rect -51473 -40198 -51177 -40172
rect -51133 -40198 -50517 -39902
rect -50473 -39928 -50177 -39902
rect -50473 -40172 -50447 -39928
rect -50447 -40172 -50203 -39928
rect -50203 -40172 -50177 -39928
rect -50473 -40198 -50177 -40172
rect -50133 -40198 -49517 -39902
rect -49473 -39928 -49177 -39902
rect -49473 -40172 -49447 -39928
rect -49447 -40172 -49203 -39928
rect -49203 -40172 -49177 -39928
rect -49473 -40198 -49177 -40172
rect -49133 -40198 -48837 -39902
rect -74473 -40858 -74177 -40242
rect -73473 -40858 -73177 -40242
rect -72473 -40858 -72177 -40242
rect -71473 -40858 -71177 -40242
rect -70473 -40858 -70177 -40242
rect -69473 -40858 -69177 -40242
rect -68473 -40858 -68177 -40242
rect -67473 -40858 -67177 -40242
rect -66473 -40858 -66177 -40242
rect -65473 -40858 -65177 -40242
rect -64473 -40858 -64177 -40242
rect -63473 -40858 -63177 -40242
rect -62473 -40858 -62177 -40242
rect -61473 -40858 -61177 -40242
rect -60473 -40858 -60177 -40242
rect -59473 -40858 -59177 -40242
rect -58473 -40858 -58177 -40242
rect -57473 -40858 -57177 -40242
rect -56473 -40858 -56177 -40242
rect -55473 -40858 -55177 -40242
rect -54473 -40858 -54177 -40242
rect -53473 -40858 -53177 -40242
rect -52473 -40858 -52177 -40242
rect -51473 -40858 -51177 -40242
rect -50473 -40858 -50177 -40242
rect -49473 -40858 -49177 -40242
rect -74813 -41198 -74517 -40902
rect -74473 -40928 -74177 -40902
rect -74473 -41172 -74447 -40928
rect -74447 -41172 -74203 -40928
rect -74203 -41172 -74177 -40928
rect -74473 -41198 -74177 -41172
rect -74133 -41198 -73517 -40902
rect -73473 -40928 -73177 -40902
rect -73473 -41172 -73447 -40928
rect -73447 -41172 -73203 -40928
rect -73203 -41172 -73177 -40928
rect -73473 -41198 -73177 -41172
rect -73133 -41198 -72517 -40902
rect -72473 -40928 -72177 -40902
rect -72473 -41172 -72447 -40928
rect -72447 -41172 -72203 -40928
rect -72203 -41172 -72177 -40928
rect -72473 -41198 -72177 -41172
rect -72133 -41198 -71517 -40902
rect -71473 -40928 -71177 -40902
rect -71473 -41172 -71447 -40928
rect -71447 -41172 -71203 -40928
rect -71203 -41172 -71177 -40928
rect -71473 -41198 -71177 -41172
rect -71133 -41198 -70517 -40902
rect -70473 -40928 -70177 -40902
rect -70473 -41172 -70447 -40928
rect -70447 -41172 -70203 -40928
rect -70203 -41172 -70177 -40928
rect -70473 -41198 -70177 -41172
rect -70133 -41198 -69517 -40902
rect -69473 -40928 -69177 -40902
rect -69473 -41172 -69447 -40928
rect -69447 -41172 -69203 -40928
rect -69203 -41172 -69177 -40928
rect -69473 -41198 -69177 -41172
rect -69133 -41198 -68517 -40902
rect -68473 -40928 -68177 -40902
rect -68473 -41172 -68447 -40928
rect -68447 -41172 -68203 -40928
rect -68203 -41172 -68177 -40928
rect -68473 -41198 -68177 -41172
rect -68133 -41198 -67517 -40902
rect -67473 -40928 -67177 -40902
rect -67473 -41172 -67447 -40928
rect -67447 -41172 -67203 -40928
rect -67203 -41172 -67177 -40928
rect -67473 -41198 -67177 -41172
rect -67133 -41198 -66517 -40902
rect -66473 -40928 -66177 -40902
rect -66473 -41172 -66447 -40928
rect -66447 -41172 -66203 -40928
rect -66203 -41172 -66177 -40928
rect -66473 -41198 -66177 -41172
rect -66133 -41198 -65517 -40902
rect -65473 -40928 -65177 -40902
rect -65473 -41172 -65447 -40928
rect -65447 -41172 -65203 -40928
rect -65203 -41172 -65177 -40928
rect -65473 -41198 -65177 -41172
rect -65133 -41198 -64517 -40902
rect -64473 -40928 -64177 -40902
rect -64473 -41172 -64447 -40928
rect -64447 -41172 -64203 -40928
rect -64203 -41172 -64177 -40928
rect -64473 -41198 -64177 -41172
rect -64133 -41198 -63517 -40902
rect -63473 -40928 -63177 -40902
rect -63473 -41172 -63447 -40928
rect -63447 -41172 -63203 -40928
rect -63203 -41172 -63177 -40928
rect -63473 -41198 -63177 -41172
rect -63133 -41198 -62517 -40902
rect -62473 -40928 -62177 -40902
rect -62473 -41172 -62447 -40928
rect -62447 -41172 -62203 -40928
rect -62203 -41172 -62177 -40928
rect -62473 -41198 -62177 -41172
rect -62133 -41198 -61517 -40902
rect -61473 -40928 -61177 -40902
rect -61473 -41172 -61447 -40928
rect -61447 -41172 -61203 -40928
rect -61203 -41172 -61177 -40928
rect -61473 -41198 -61177 -41172
rect -61133 -41198 -60517 -40902
rect -60473 -40928 -60177 -40902
rect -60473 -41172 -60447 -40928
rect -60447 -41172 -60203 -40928
rect -60203 -41172 -60177 -40928
rect -60473 -41198 -60177 -41172
rect -60133 -41198 -59517 -40902
rect -59473 -40928 -59177 -40902
rect -59473 -41172 -59447 -40928
rect -59447 -41172 -59203 -40928
rect -59203 -41172 -59177 -40928
rect -59473 -41198 -59177 -41172
rect -59133 -41198 -58517 -40902
rect -58473 -40928 -58177 -40902
rect -58473 -41172 -58447 -40928
rect -58447 -41172 -58203 -40928
rect -58203 -41172 -58177 -40928
rect -58473 -41198 -58177 -41172
rect -58133 -41198 -57517 -40902
rect -57473 -40928 -57177 -40902
rect -57473 -41172 -57447 -40928
rect -57447 -41172 -57203 -40928
rect -57203 -41172 -57177 -40928
rect -57473 -41198 -57177 -41172
rect -57133 -41198 -56517 -40902
rect -56473 -40928 -56177 -40902
rect -56473 -41172 -56447 -40928
rect -56447 -41172 -56203 -40928
rect -56203 -41172 -56177 -40928
rect -56473 -41198 -56177 -41172
rect -56133 -41198 -55517 -40902
rect -55473 -40928 -55177 -40902
rect -55473 -41172 -55447 -40928
rect -55447 -41172 -55203 -40928
rect -55203 -41172 -55177 -40928
rect -55473 -41198 -55177 -41172
rect -55133 -41198 -54517 -40902
rect -54473 -40928 -54177 -40902
rect -54473 -41172 -54447 -40928
rect -54447 -41172 -54203 -40928
rect -54203 -41172 -54177 -40928
rect -54473 -41198 -54177 -41172
rect -54133 -41198 -53517 -40902
rect -53473 -40928 -53177 -40902
rect -53473 -41172 -53447 -40928
rect -53447 -41172 -53203 -40928
rect -53203 -41172 -53177 -40928
rect -53473 -41198 -53177 -41172
rect -53133 -41198 -52517 -40902
rect -52473 -40928 -52177 -40902
rect -52473 -41172 -52447 -40928
rect -52447 -41172 -52203 -40928
rect -52203 -41172 -52177 -40928
rect -52473 -41198 -52177 -41172
rect -52133 -41198 -51517 -40902
rect -51473 -40928 -51177 -40902
rect -51473 -41172 -51447 -40928
rect -51447 -41172 -51203 -40928
rect -51203 -41172 -51177 -40928
rect -51473 -41198 -51177 -41172
rect -51133 -41198 -50517 -40902
rect -50473 -40928 -50177 -40902
rect -50473 -41172 -50447 -40928
rect -50447 -41172 -50203 -40928
rect -50203 -41172 -50177 -40928
rect -50473 -41198 -50177 -41172
rect -50133 -41198 -49517 -40902
rect -49473 -40928 -49177 -40902
rect -49473 -41172 -49447 -40928
rect -49447 -41172 -49203 -40928
rect -49203 -41172 -49177 -40928
rect -49473 -41198 -49177 -41172
rect -49133 -41198 -48837 -40902
rect -74473 -41858 -74177 -41242
rect -73473 -41858 -73177 -41242
rect -72473 -41858 -72177 -41242
rect -71473 -41858 -71177 -41242
rect -70473 -41858 -70177 -41242
rect -69473 -41858 -69177 -41242
rect -68473 -41858 -68177 -41242
rect -67473 -41858 -67177 -41242
rect -66473 -41858 -66177 -41242
rect -65473 -41858 -65177 -41242
rect -64473 -41858 -64177 -41242
rect -63473 -41858 -63177 -41242
rect -62473 -41858 -62177 -41242
rect -61473 -41858 -61177 -41242
rect -60473 -41858 -60177 -41242
rect -59473 -41858 -59177 -41242
rect -58473 -41858 -58177 -41242
rect -57473 -41858 -57177 -41242
rect -56473 -41858 -56177 -41242
rect -55473 -41858 -55177 -41242
rect -54473 -41858 -54177 -41242
rect -53473 -41858 -53177 -41242
rect -52473 -41858 -52177 -41242
rect -51473 -41858 -51177 -41242
rect -50473 -41858 -50177 -41242
rect -49473 -41858 -49177 -41242
rect -74813 -42198 -74517 -41902
rect -74473 -41928 -74177 -41902
rect -74473 -42172 -74447 -41928
rect -74447 -42172 -74203 -41928
rect -74203 -42172 -74177 -41928
rect -74473 -42198 -74177 -42172
rect -74133 -42198 -73517 -41902
rect -73473 -41928 -73177 -41902
rect -73473 -42172 -73447 -41928
rect -73447 -42172 -73203 -41928
rect -73203 -42172 -73177 -41928
rect -73473 -42198 -73177 -42172
rect -73133 -42198 -72517 -41902
rect -72473 -41928 -72177 -41902
rect -72473 -42172 -72447 -41928
rect -72447 -42172 -72203 -41928
rect -72203 -42172 -72177 -41928
rect -72473 -42198 -72177 -42172
rect -72133 -42198 -71517 -41902
rect -71473 -41928 -71177 -41902
rect -71473 -42172 -71447 -41928
rect -71447 -42172 -71203 -41928
rect -71203 -42172 -71177 -41928
rect -71473 -42198 -71177 -42172
rect -71133 -42198 -70517 -41902
rect -70473 -41928 -70177 -41902
rect -70473 -42172 -70447 -41928
rect -70447 -42172 -70203 -41928
rect -70203 -42172 -70177 -41928
rect -70473 -42198 -70177 -42172
rect -70133 -42198 -69517 -41902
rect -69473 -41928 -69177 -41902
rect -69473 -42172 -69447 -41928
rect -69447 -42172 -69203 -41928
rect -69203 -42172 -69177 -41928
rect -69473 -42198 -69177 -42172
rect -69133 -42198 -68517 -41902
rect -68473 -41928 -68177 -41902
rect -68473 -42172 -68447 -41928
rect -68447 -42172 -68203 -41928
rect -68203 -42172 -68177 -41928
rect -68473 -42198 -68177 -42172
rect -68133 -42198 -67517 -41902
rect -67473 -41928 -67177 -41902
rect -67473 -42172 -67447 -41928
rect -67447 -42172 -67203 -41928
rect -67203 -42172 -67177 -41928
rect -67473 -42198 -67177 -42172
rect -67133 -42198 -66517 -41902
rect -66473 -41928 -66177 -41902
rect -66473 -42172 -66447 -41928
rect -66447 -42172 -66203 -41928
rect -66203 -42172 -66177 -41928
rect -66473 -42198 -66177 -42172
rect -66133 -42198 -65517 -41902
rect -65473 -41928 -65177 -41902
rect -65473 -42172 -65447 -41928
rect -65447 -42172 -65203 -41928
rect -65203 -42172 -65177 -41928
rect -65473 -42198 -65177 -42172
rect -65133 -42198 -64517 -41902
rect -64473 -41928 -64177 -41902
rect -64473 -42172 -64447 -41928
rect -64447 -42172 -64203 -41928
rect -64203 -42172 -64177 -41928
rect -64473 -42198 -64177 -42172
rect -64133 -42198 -63517 -41902
rect -63473 -41928 -63177 -41902
rect -63473 -42172 -63447 -41928
rect -63447 -42172 -63203 -41928
rect -63203 -42172 -63177 -41928
rect -63473 -42198 -63177 -42172
rect -63133 -42198 -62517 -41902
rect -62473 -41928 -62177 -41902
rect -62473 -42172 -62447 -41928
rect -62447 -42172 -62203 -41928
rect -62203 -42172 -62177 -41928
rect -62473 -42198 -62177 -42172
rect -62133 -42198 -61517 -41902
rect -61473 -41928 -61177 -41902
rect -61473 -42172 -61447 -41928
rect -61447 -42172 -61203 -41928
rect -61203 -42172 -61177 -41928
rect -61473 -42198 -61177 -42172
rect -61133 -42198 -60517 -41902
rect -60473 -41928 -60177 -41902
rect -60473 -42172 -60447 -41928
rect -60447 -42172 -60203 -41928
rect -60203 -42172 -60177 -41928
rect -60473 -42198 -60177 -42172
rect -60133 -42198 -59517 -41902
rect -59473 -41928 -59177 -41902
rect -59473 -42172 -59447 -41928
rect -59447 -42172 -59203 -41928
rect -59203 -42172 -59177 -41928
rect -59473 -42198 -59177 -42172
rect -59133 -42198 -58517 -41902
rect -58473 -41928 -58177 -41902
rect -58473 -42172 -58447 -41928
rect -58447 -42172 -58203 -41928
rect -58203 -42172 -58177 -41928
rect -58473 -42198 -58177 -42172
rect -58133 -42198 -57517 -41902
rect -57473 -41928 -57177 -41902
rect -57473 -42172 -57447 -41928
rect -57447 -42172 -57203 -41928
rect -57203 -42172 -57177 -41928
rect -57473 -42198 -57177 -42172
rect -57133 -42198 -56517 -41902
rect -56473 -41928 -56177 -41902
rect -56473 -42172 -56447 -41928
rect -56447 -42172 -56203 -41928
rect -56203 -42172 -56177 -41928
rect -56473 -42198 -56177 -42172
rect -56133 -42198 -55517 -41902
rect -55473 -41928 -55177 -41902
rect -55473 -42172 -55447 -41928
rect -55447 -42172 -55203 -41928
rect -55203 -42172 -55177 -41928
rect -55473 -42198 -55177 -42172
rect -55133 -42198 -54517 -41902
rect -54473 -41928 -54177 -41902
rect -54473 -42172 -54447 -41928
rect -54447 -42172 -54203 -41928
rect -54203 -42172 -54177 -41928
rect -54473 -42198 -54177 -42172
rect -54133 -42198 -53517 -41902
rect -53473 -41928 -53177 -41902
rect -53473 -42172 -53447 -41928
rect -53447 -42172 -53203 -41928
rect -53203 -42172 -53177 -41928
rect -53473 -42198 -53177 -42172
rect -53133 -42198 -52517 -41902
rect -52473 -41928 -52177 -41902
rect -52473 -42172 -52447 -41928
rect -52447 -42172 -52203 -41928
rect -52203 -42172 -52177 -41928
rect -52473 -42198 -52177 -42172
rect -52133 -42198 -51517 -41902
rect -51473 -41928 -51177 -41902
rect -51473 -42172 -51447 -41928
rect -51447 -42172 -51203 -41928
rect -51203 -42172 -51177 -41928
rect -51473 -42198 -51177 -42172
rect -51133 -42198 -50517 -41902
rect -50473 -41928 -50177 -41902
rect -50473 -42172 -50447 -41928
rect -50447 -42172 -50203 -41928
rect -50203 -42172 -50177 -41928
rect -50473 -42198 -50177 -42172
rect -50133 -42198 -49517 -41902
rect -49473 -41928 -49177 -41902
rect -49473 -42172 -49447 -41928
rect -49447 -42172 -49203 -41928
rect -49203 -42172 -49177 -41928
rect -49473 -42198 -49177 -42172
rect -49133 -42198 -48837 -41902
rect -74473 -42858 -74177 -42242
rect -73473 -42858 -73177 -42242
rect -72473 -42858 -72177 -42242
rect -71473 -42858 -71177 -42242
rect -70473 -42858 -70177 -42242
rect -69473 -42858 -69177 -42242
rect -68473 -42858 -68177 -42242
rect -67473 -42858 -67177 -42242
rect -66473 -42858 -66177 -42242
rect -65473 -42858 -65177 -42242
rect -64473 -42858 -64177 -42242
rect -63473 -42858 -63177 -42242
rect -62473 -42858 -62177 -42242
rect -61473 -42858 -61177 -42242
rect -60473 -42858 -60177 -42242
rect -59473 -42858 -59177 -42242
rect -58473 -42858 -58177 -42242
rect -57473 -42858 -57177 -42242
rect -56473 -42858 -56177 -42242
rect -55473 -42858 -55177 -42242
rect -54473 -42858 -54177 -42242
rect -53473 -42858 -53177 -42242
rect -52473 -42858 -52177 -42242
rect -51473 -42858 -51177 -42242
rect -50473 -42858 -50177 -42242
rect -49473 -42858 -49177 -42242
rect -74813 -43198 -74517 -42902
rect -74473 -42928 -74177 -42902
rect -74473 -43172 -74447 -42928
rect -74447 -43172 -74203 -42928
rect -74203 -43172 -74177 -42928
rect -74473 -43198 -74177 -43172
rect -74133 -43198 -73517 -42902
rect -73473 -42928 -73177 -42902
rect -73473 -43172 -73447 -42928
rect -73447 -43172 -73203 -42928
rect -73203 -43172 -73177 -42928
rect -73473 -43198 -73177 -43172
rect -73133 -43198 -72517 -42902
rect -72473 -42928 -72177 -42902
rect -72473 -43172 -72447 -42928
rect -72447 -43172 -72203 -42928
rect -72203 -43172 -72177 -42928
rect -72473 -43198 -72177 -43172
rect -72133 -43198 -71517 -42902
rect -71473 -42928 -71177 -42902
rect -71473 -43172 -71447 -42928
rect -71447 -43172 -71203 -42928
rect -71203 -43172 -71177 -42928
rect -71473 -43198 -71177 -43172
rect -71133 -43198 -70517 -42902
rect -70473 -42928 -70177 -42902
rect -70473 -43172 -70447 -42928
rect -70447 -43172 -70203 -42928
rect -70203 -43172 -70177 -42928
rect -70473 -43198 -70177 -43172
rect -70133 -43198 -69517 -42902
rect -69473 -42928 -69177 -42902
rect -69473 -43172 -69447 -42928
rect -69447 -43172 -69203 -42928
rect -69203 -43172 -69177 -42928
rect -69473 -43198 -69177 -43172
rect -69133 -43198 -68517 -42902
rect -68473 -42928 -68177 -42902
rect -68473 -43172 -68447 -42928
rect -68447 -43172 -68203 -42928
rect -68203 -43172 -68177 -42928
rect -68473 -43198 -68177 -43172
rect -68133 -43198 -67517 -42902
rect -67473 -42928 -67177 -42902
rect -67473 -43172 -67447 -42928
rect -67447 -43172 -67203 -42928
rect -67203 -43172 -67177 -42928
rect -67473 -43198 -67177 -43172
rect -67133 -43198 -66517 -42902
rect -66473 -42928 -66177 -42902
rect -66473 -43172 -66447 -42928
rect -66447 -43172 -66203 -42928
rect -66203 -43172 -66177 -42928
rect -66473 -43198 -66177 -43172
rect -66133 -43198 -65517 -42902
rect -65473 -42928 -65177 -42902
rect -65473 -43172 -65447 -42928
rect -65447 -43172 -65203 -42928
rect -65203 -43172 -65177 -42928
rect -65473 -43198 -65177 -43172
rect -65133 -43198 -64517 -42902
rect -64473 -42928 -64177 -42902
rect -64473 -43172 -64447 -42928
rect -64447 -43172 -64203 -42928
rect -64203 -43172 -64177 -42928
rect -64473 -43198 -64177 -43172
rect -64133 -43198 -63517 -42902
rect -63473 -42928 -63177 -42902
rect -63473 -43172 -63447 -42928
rect -63447 -43172 -63203 -42928
rect -63203 -43172 -63177 -42928
rect -63473 -43198 -63177 -43172
rect -63133 -43198 -62517 -42902
rect -62473 -42928 -62177 -42902
rect -62473 -43172 -62447 -42928
rect -62447 -43172 -62203 -42928
rect -62203 -43172 -62177 -42928
rect -62473 -43198 -62177 -43172
rect -62133 -43198 -61517 -42902
rect -61473 -42928 -61177 -42902
rect -61473 -43172 -61447 -42928
rect -61447 -43172 -61203 -42928
rect -61203 -43172 -61177 -42928
rect -61473 -43198 -61177 -43172
rect -61133 -43198 -60517 -42902
rect -60473 -42928 -60177 -42902
rect -60473 -43172 -60447 -42928
rect -60447 -43172 -60203 -42928
rect -60203 -43172 -60177 -42928
rect -60473 -43198 -60177 -43172
rect -60133 -43198 -59517 -42902
rect -59473 -42928 -59177 -42902
rect -59473 -43172 -59447 -42928
rect -59447 -43172 -59203 -42928
rect -59203 -43172 -59177 -42928
rect -59473 -43198 -59177 -43172
rect -59133 -43198 -58517 -42902
rect -58473 -42928 -58177 -42902
rect -58473 -43172 -58447 -42928
rect -58447 -43172 -58203 -42928
rect -58203 -43172 -58177 -42928
rect -58473 -43198 -58177 -43172
rect -58133 -43198 -57517 -42902
rect -57473 -42928 -57177 -42902
rect -57473 -43172 -57447 -42928
rect -57447 -43172 -57203 -42928
rect -57203 -43172 -57177 -42928
rect -57473 -43198 -57177 -43172
rect -57133 -43198 -56517 -42902
rect -56473 -42928 -56177 -42902
rect -56473 -43172 -56447 -42928
rect -56447 -43172 -56203 -42928
rect -56203 -43172 -56177 -42928
rect -56473 -43198 -56177 -43172
rect -56133 -43198 -55517 -42902
rect -55473 -42928 -55177 -42902
rect -55473 -43172 -55447 -42928
rect -55447 -43172 -55203 -42928
rect -55203 -43172 -55177 -42928
rect -55473 -43198 -55177 -43172
rect -55133 -43198 -54517 -42902
rect -54473 -42928 -54177 -42902
rect -54473 -43172 -54447 -42928
rect -54447 -43172 -54203 -42928
rect -54203 -43172 -54177 -42928
rect -54473 -43198 -54177 -43172
rect -54133 -43198 -53517 -42902
rect -53473 -42928 -53177 -42902
rect -53473 -43172 -53447 -42928
rect -53447 -43172 -53203 -42928
rect -53203 -43172 -53177 -42928
rect -53473 -43198 -53177 -43172
rect -53133 -43198 -52517 -42902
rect -52473 -42928 -52177 -42902
rect -52473 -43172 -52447 -42928
rect -52447 -43172 -52203 -42928
rect -52203 -43172 -52177 -42928
rect -52473 -43198 -52177 -43172
rect -52133 -43198 -51517 -42902
rect -51473 -42928 -51177 -42902
rect -51473 -43172 -51447 -42928
rect -51447 -43172 -51203 -42928
rect -51203 -43172 -51177 -42928
rect -51473 -43198 -51177 -43172
rect -51133 -43198 -50517 -42902
rect -50473 -42928 -50177 -42902
rect -50473 -43172 -50447 -42928
rect -50447 -43172 -50203 -42928
rect -50203 -43172 -50177 -42928
rect -50473 -43198 -50177 -43172
rect -50133 -43198 -49517 -42902
rect -49473 -42928 -49177 -42902
rect -49473 -43172 -49447 -42928
rect -49447 -43172 -49203 -42928
rect -49203 -43172 -49177 -42928
rect -49473 -43198 -49177 -43172
rect -49133 -43198 -48837 -42902
rect -74473 -43858 -74177 -43242
rect -73473 -43858 -73177 -43242
rect -72473 -43858 -72177 -43242
rect -71473 -43858 -71177 -43242
rect -70473 -43858 -70177 -43242
rect -69473 -43858 -69177 -43242
rect -68473 -43858 -68177 -43242
rect -67473 -43858 -67177 -43242
rect -66473 -43858 -66177 -43242
rect -65473 -43858 -65177 -43242
rect -64473 -43858 -64177 -43242
rect -63473 -43858 -63177 -43242
rect -62473 -43858 -62177 -43242
rect -61473 -43858 -61177 -43242
rect -60473 -43858 -60177 -43242
rect -59473 -43858 -59177 -43242
rect -58473 -43858 -58177 -43242
rect -57473 -43858 -57177 -43242
rect -56473 -43858 -56177 -43242
rect -55473 -43858 -55177 -43242
rect -54473 -43858 -54177 -43242
rect -53473 -43858 -53177 -43242
rect -52473 -43858 -52177 -43242
rect -51473 -43858 -51177 -43242
rect -50473 -43858 -50177 -43242
rect -49473 -43858 -49177 -43242
rect -74813 -44198 -74517 -43902
rect -74473 -43928 -74177 -43902
rect -74473 -44172 -74447 -43928
rect -74447 -44172 -74203 -43928
rect -74203 -44172 -74177 -43928
rect -74473 -44198 -74177 -44172
rect -74133 -44198 -73517 -43902
rect -73473 -43928 -73177 -43902
rect -73473 -44172 -73447 -43928
rect -73447 -44172 -73203 -43928
rect -73203 -44172 -73177 -43928
rect -73473 -44198 -73177 -44172
rect -73133 -44198 -72517 -43902
rect -72473 -43928 -72177 -43902
rect -72473 -44172 -72447 -43928
rect -72447 -44172 -72203 -43928
rect -72203 -44172 -72177 -43928
rect -72473 -44198 -72177 -44172
rect -72133 -44198 -71517 -43902
rect -71473 -43928 -71177 -43902
rect -71473 -44172 -71447 -43928
rect -71447 -44172 -71203 -43928
rect -71203 -44172 -71177 -43928
rect -71473 -44198 -71177 -44172
rect -71133 -44198 -70517 -43902
rect -70473 -43928 -70177 -43902
rect -70473 -44172 -70447 -43928
rect -70447 -44172 -70203 -43928
rect -70203 -44172 -70177 -43928
rect -70473 -44198 -70177 -44172
rect -70133 -44198 -69517 -43902
rect -69473 -43928 -69177 -43902
rect -69473 -44172 -69447 -43928
rect -69447 -44172 -69203 -43928
rect -69203 -44172 -69177 -43928
rect -69473 -44198 -69177 -44172
rect -69133 -44198 -68517 -43902
rect -68473 -43928 -68177 -43902
rect -68473 -44172 -68447 -43928
rect -68447 -44172 -68203 -43928
rect -68203 -44172 -68177 -43928
rect -68473 -44198 -68177 -44172
rect -68133 -44198 -67517 -43902
rect -67473 -43928 -67177 -43902
rect -67473 -44172 -67447 -43928
rect -67447 -44172 -67203 -43928
rect -67203 -44172 -67177 -43928
rect -67473 -44198 -67177 -44172
rect -67133 -44198 -66517 -43902
rect -66473 -43928 -66177 -43902
rect -66473 -44172 -66447 -43928
rect -66447 -44172 -66203 -43928
rect -66203 -44172 -66177 -43928
rect -66473 -44198 -66177 -44172
rect -66133 -44198 -65517 -43902
rect -65473 -43928 -65177 -43902
rect -65473 -44172 -65447 -43928
rect -65447 -44172 -65203 -43928
rect -65203 -44172 -65177 -43928
rect -65473 -44198 -65177 -44172
rect -65133 -44198 -64517 -43902
rect -64473 -43928 -64177 -43902
rect -64473 -44172 -64447 -43928
rect -64447 -44172 -64203 -43928
rect -64203 -44172 -64177 -43928
rect -64473 -44198 -64177 -44172
rect -64133 -44198 -63517 -43902
rect -63473 -43928 -63177 -43902
rect -63473 -44172 -63447 -43928
rect -63447 -44172 -63203 -43928
rect -63203 -44172 -63177 -43928
rect -63473 -44198 -63177 -44172
rect -63133 -44198 -62517 -43902
rect -62473 -43928 -62177 -43902
rect -62473 -44172 -62447 -43928
rect -62447 -44172 -62203 -43928
rect -62203 -44172 -62177 -43928
rect -62473 -44198 -62177 -44172
rect -62133 -44198 -61517 -43902
rect -61473 -43928 -61177 -43902
rect -61473 -44172 -61447 -43928
rect -61447 -44172 -61203 -43928
rect -61203 -44172 -61177 -43928
rect -61473 -44198 -61177 -44172
rect -61133 -44198 -60517 -43902
rect -60473 -43928 -60177 -43902
rect -60473 -44172 -60447 -43928
rect -60447 -44172 -60203 -43928
rect -60203 -44172 -60177 -43928
rect -60473 -44198 -60177 -44172
rect -60133 -44198 -59517 -43902
rect -59473 -43928 -59177 -43902
rect -59473 -44172 -59447 -43928
rect -59447 -44172 -59203 -43928
rect -59203 -44172 -59177 -43928
rect -59473 -44198 -59177 -44172
rect -59133 -44198 -58517 -43902
rect -58473 -43928 -58177 -43902
rect -58473 -44172 -58447 -43928
rect -58447 -44172 -58203 -43928
rect -58203 -44172 -58177 -43928
rect -58473 -44198 -58177 -44172
rect -58133 -44198 -57517 -43902
rect -57473 -43928 -57177 -43902
rect -57473 -44172 -57447 -43928
rect -57447 -44172 -57203 -43928
rect -57203 -44172 -57177 -43928
rect -57473 -44198 -57177 -44172
rect -57133 -44198 -56517 -43902
rect -56473 -43928 -56177 -43902
rect -56473 -44172 -56447 -43928
rect -56447 -44172 -56203 -43928
rect -56203 -44172 -56177 -43928
rect -56473 -44198 -56177 -44172
rect -56133 -44198 -55517 -43902
rect -55473 -43928 -55177 -43902
rect -55473 -44172 -55447 -43928
rect -55447 -44172 -55203 -43928
rect -55203 -44172 -55177 -43928
rect -55473 -44198 -55177 -44172
rect -55133 -44198 -54517 -43902
rect -54473 -43928 -54177 -43902
rect -54473 -44172 -54447 -43928
rect -54447 -44172 -54203 -43928
rect -54203 -44172 -54177 -43928
rect -54473 -44198 -54177 -44172
rect -54133 -44198 -53517 -43902
rect -53473 -43928 -53177 -43902
rect -53473 -44172 -53447 -43928
rect -53447 -44172 -53203 -43928
rect -53203 -44172 -53177 -43928
rect -53473 -44198 -53177 -44172
rect -53133 -44198 -52517 -43902
rect -52473 -43928 -52177 -43902
rect -52473 -44172 -52447 -43928
rect -52447 -44172 -52203 -43928
rect -52203 -44172 -52177 -43928
rect -52473 -44198 -52177 -44172
rect -52133 -44198 -51517 -43902
rect -51473 -43928 -51177 -43902
rect -51473 -44172 -51447 -43928
rect -51447 -44172 -51203 -43928
rect -51203 -44172 -51177 -43928
rect -51473 -44198 -51177 -44172
rect -51133 -44198 -50517 -43902
rect -50473 -43928 -50177 -43902
rect -50473 -44172 -50447 -43928
rect -50447 -44172 -50203 -43928
rect -50203 -44172 -50177 -43928
rect -50473 -44198 -50177 -44172
rect -50133 -44198 -49517 -43902
rect -49473 -43928 -49177 -43902
rect -49473 -44172 -49447 -43928
rect -49447 -44172 -49203 -43928
rect -49203 -44172 -49177 -43928
rect -49473 -44198 -49177 -44172
rect -49133 -44198 -48837 -43902
rect -74473 -44858 -74177 -44242
rect -73473 -44858 -73177 -44242
rect -72473 -44858 -72177 -44242
rect -71473 -44858 -71177 -44242
rect -70473 -44858 -70177 -44242
rect -69473 -44858 -69177 -44242
rect -68473 -44858 -68177 -44242
rect -67473 -44858 -67177 -44242
rect -66473 -44858 -66177 -44242
rect -65473 -44858 -65177 -44242
rect -64473 -44858 -64177 -44242
rect -63473 -44858 -63177 -44242
rect -62473 -44858 -62177 -44242
rect -61473 -44858 -61177 -44242
rect -60473 -44858 -60177 -44242
rect -59473 -44858 -59177 -44242
rect -58473 -44858 -58177 -44242
rect -57473 -44858 -57177 -44242
rect -56473 -44858 -56177 -44242
rect -55473 -44858 -55177 -44242
rect -54473 -44858 -54177 -44242
rect -53473 -44858 -53177 -44242
rect -52473 -44858 -52177 -44242
rect -51473 -44858 -51177 -44242
rect -50473 -44858 -50177 -44242
rect -49473 -44858 -49177 -44242
rect -46228 -44496 -36332 -32604
rect -46228 -44498 -36332 -44496
rect -4228 -32604 5668 -32602
rect -4228 -44496 5668 -32604
rect 8627 -32858 8923 -32242
rect 9627 -32858 9923 -32242
rect 10627 -32858 10923 -32242
rect 11627 -32858 11923 -32242
rect 12627 -32858 12923 -32242
rect 13627 -32858 13923 -32242
rect 14627 -32858 14923 -32242
rect 15627 -32858 15923 -32242
rect 16627 -32858 16923 -32242
rect 17627 -32858 17923 -32242
rect 18627 -32858 18923 -32242
rect 19627 -32858 19923 -32242
rect 20627 -32858 20923 -32242
rect 21627 -32858 21923 -32242
rect 22627 -32858 22923 -32242
rect 23627 -32858 23923 -32242
rect 24627 -32858 24923 -32242
rect 25627 -32858 25923 -32242
rect 26627 -32858 26923 -32242
rect 27627 -32858 27923 -32242
rect 28627 -32858 28923 -32242
rect 29627 -32858 29923 -32242
rect 30627 -32858 30923 -32242
rect 31627 -32858 31923 -32242
rect 32627 -32858 32923 -32242
rect 33627 -32858 33923 -32242
rect 8287 -33198 8583 -32902
rect 8627 -32928 8923 -32902
rect 8627 -33172 8653 -32928
rect 8653 -33172 8897 -32928
rect 8897 -33172 8923 -32928
rect 8627 -33198 8923 -33172
rect 8967 -33198 9583 -32902
rect 9627 -32928 9923 -32902
rect 9627 -33172 9653 -32928
rect 9653 -33172 9897 -32928
rect 9897 -33172 9923 -32928
rect 9627 -33198 9923 -33172
rect 9967 -33198 10583 -32902
rect 10627 -32928 10923 -32902
rect 10627 -33172 10653 -32928
rect 10653 -33172 10897 -32928
rect 10897 -33172 10923 -32928
rect 10627 -33198 10923 -33172
rect 10967 -33198 11583 -32902
rect 11627 -32928 11923 -32902
rect 11627 -33172 11653 -32928
rect 11653 -33172 11897 -32928
rect 11897 -33172 11923 -32928
rect 11627 -33198 11923 -33172
rect 11967 -33198 12583 -32902
rect 12627 -32928 12923 -32902
rect 12627 -33172 12653 -32928
rect 12653 -33172 12897 -32928
rect 12897 -33172 12923 -32928
rect 12627 -33198 12923 -33172
rect 12967 -33198 13583 -32902
rect 13627 -32928 13923 -32902
rect 13627 -33172 13653 -32928
rect 13653 -33172 13897 -32928
rect 13897 -33172 13923 -32928
rect 13627 -33198 13923 -33172
rect 13967 -33198 14583 -32902
rect 14627 -32928 14923 -32902
rect 14627 -33172 14653 -32928
rect 14653 -33172 14897 -32928
rect 14897 -33172 14923 -32928
rect 14627 -33198 14923 -33172
rect 14967 -33198 15583 -32902
rect 15627 -32928 15923 -32902
rect 15627 -33172 15653 -32928
rect 15653 -33172 15897 -32928
rect 15897 -33172 15923 -32928
rect 15627 -33198 15923 -33172
rect 15967 -33198 16583 -32902
rect 16627 -32928 16923 -32902
rect 16627 -33172 16653 -32928
rect 16653 -33172 16897 -32928
rect 16897 -33172 16923 -32928
rect 16627 -33198 16923 -33172
rect 16967 -33198 17583 -32902
rect 17627 -32928 17923 -32902
rect 17627 -33172 17653 -32928
rect 17653 -33172 17897 -32928
rect 17897 -33172 17923 -32928
rect 17627 -33198 17923 -33172
rect 17967 -33198 18583 -32902
rect 18627 -32928 18923 -32902
rect 18627 -33172 18653 -32928
rect 18653 -33172 18897 -32928
rect 18897 -33172 18923 -32928
rect 18627 -33198 18923 -33172
rect 18967 -33198 19583 -32902
rect 19627 -32928 19923 -32902
rect 19627 -33172 19653 -32928
rect 19653 -33172 19897 -32928
rect 19897 -33172 19923 -32928
rect 19627 -33198 19923 -33172
rect 19967 -33198 20583 -32902
rect 20627 -32928 20923 -32902
rect 20627 -33172 20653 -32928
rect 20653 -33172 20897 -32928
rect 20897 -33172 20923 -32928
rect 20627 -33198 20923 -33172
rect 20967 -33198 21583 -32902
rect 21627 -32928 21923 -32902
rect 21627 -33172 21653 -32928
rect 21653 -33172 21897 -32928
rect 21897 -33172 21923 -32928
rect 21627 -33198 21923 -33172
rect 21967 -33198 22583 -32902
rect 22627 -32928 22923 -32902
rect 22627 -33172 22653 -32928
rect 22653 -33172 22897 -32928
rect 22897 -33172 22923 -32928
rect 22627 -33198 22923 -33172
rect 22967 -33198 23583 -32902
rect 23627 -32928 23923 -32902
rect 23627 -33172 23653 -32928
rect 23653 -33172 23897 -32928
rect 23897 -33172 23923 -32928
rect 23627 -33198 23923 -33172
rect 23967 -33198 24583 -32902
rect 24627 -32928 24923 -32902
rect 24627 -33172 24653 -32928
rect 24653 -33172 24897 -32928
rect 24897 -33172 24923 -32928
rect 24627 -33198 24923 -33172
rect 24967 -33198 25583 -32902
rect 25627 -32928 25923 -32902
rect 25627 -33172 25653 -32928
rect 25653 -33172 25897 -32928
rect 25897 -33172 25923 -32928
rect 25627 -33198 25923 -33172
rect 25967 -33198 26583 -32902
rect 26627 -32928 26923 -32902
rect 26627 -33172 26653 -32928
rect 26653 -33172 26897 -32928
rect 26897 -33172 26923 -32928
rect 26627 -33198 26923 -33172
rect 26967 -33198 27583 -32902
rect 27627 -32928 27923 -32902
rect 27627 -33172 27653 -32928
rect 27653 -33172 27897 -32928
rect 27897 -33172 27923 -32928
rect 27627 -33198 27923 -33172
rect 27967 -33198 28583 -32902
rect 28627 -32928 28923 -32902
rect 28627 -33172 28653 -32928
rect 28653 -33172 28897 -32928
rect 28897 -33172 28923 -32928
rect 28627 -33198 28923 -33172
rect 28967 -33198 29583 -32902
rect 29627 -32928 29923 -32902
rect 29627 -33172 29653 -32928
rect 29653 -33172 29897 -32928
rect 29897 -33172 29923 -32928
rect 29627 -33198 29923 -33172
rect 29967 -33198 30583 -32902
rect 30627 -32928 30923 -32902
rect 30627 -33172 30653 -32928
rect 30653 -33172 30897 -32928
rect 30897 -33172 30923 -32928
rect 30627 -33198 30923 -33172
rect 30967 -33198 31583 -32902
rect 31627 -32928 31923 -32902
rect 31627 -33172 31653 -32928
rect 31653 -33172 31897 -32928
rect 31897 -33172 31923 -32928
rect 31627 -33198 31923 -33172
rect 31967 -33198 32583 -32902
rect 32627 -32928 32923 -32902
rect 32627 -33172 32653 -32928
rect 32653 -33172 32897 -32928
rect 32897 -33172 32923 -32928
rect 32627 -33198 32923 -33172
rect 32967 -33198 33583 -32902
rect 33627 -32928 33923 -32902
rect 33627 -33172 33653 -32928
rect 33653 -33172 33897 -32928
rect 33897 -33172 33923 -32928
rect 33627 -33198 33923 -33172
rect 33967 -33198 34263 -32902
rect 8627 -33858 8923 -33242
rect 9627 -33858 9923 -33242
rect 10627 -33858 10923 -33242
rect 11627 -33858 11923 -33242
rect 12627 -33858 12923 -33242
rect 13627 -33858 13923 -33242
rect 14627 -33858 14923 -33242
rect 15627 -33858 15923 -33242
rect 16627 -33858 16923 -33242
rect 17627 -33858 17923 -33242
rect 18627 -33858 18923 -33242
rect 19627 -33858 19923 -33242
rect 20627 -33858 20923 -33242
rect 21627 -33858 21923 -33242
rect 22627 -33858 22923 -33242
rect 23627 -33858 23923 -33242
rect 24627 -33858 24923 -33242
rect 25627 -33858 25923 -33242
rect 26627 -33858 26923 -33242
rect 27627 -33858 27923 -33242
rect 28627 -33858 28923 -33242
rect 29627 -33858 29923 -33242
rect 30627 -33858 30923 -33242
rect 31627 -33858 31923 -33242
rect 32627 -33858 32923 -33242
rect 33627 -33858 33923 -33242
rect 8287 -34198 8583 -33902
rect 8627 -33928 8923 -33902
rect 8627 -34172 8653 -33928
rect 8653 -34172 8897 -33928
rect 8897 -34172 8923 -33928
rect 8627 -34198 8923 -34172
rect 8967 -34198 9583 -33902
rect 9627 -33928 9923 -33902
rect 9627 -34172 9653 -33928
rect 9653 -34172 9897 -33928
rect 9897 -34172 9923 -33928
rect 9627 -34198 9923 -34172
rect 9967 -34198 10583 -33902
rect 10627 -33928 10923 -33902
rect 10627 -34172 10653 -33928
rect 10653 -34172 10897 -33928
rect 10897 -34172 10923 -33928
rect 10627 -34198 10923 -34172
rect 10967 -34198 11583 -33902
rect 11627 -33928 11923 -33902
rect 11627 -34172 11653 -33928
rect 11653 -34172 11897 -33928
rect 11897 -34172 11923 -33928
rect 11627 -34198 11923 -34172
rect 11967 -34198 12583 -33902
rect 12627 -33928 12923 -33902
rect 12627 -34172 12653 -33928
rect 12653 -34172 12897 -33928
rect 12897 -34172 12923 -33928
rect 12627 -34198 12923 -34172
rect 12967 -34198 13583 -33902
rect 13627 -33928 13923 -33902
rect 13627 -34172 13653 -33928
rect 13653 -34172 13897 -33928
rect 13897 -34172 13923 -33928
rect 13627 -34198 13923 -34172
rect 13967 -34198 14583 -33902
rect 14627 -33928 14923 -33902
rect 14627 -34172 14653 -33928
rect 14653 -34172 14897 -33928
rect 14897 -34172 14923 -33928
rect 14627 -34198 14923 -34172
rect 14967 -34198 15583 -33902
rect 15627 -33928 15923 -33902
rect 15627 -34172 15653 -33928
rect 15653 -34172 15897 -33928
rect 15897 -34172 15923 -33928
rect 15627 -34198 15923 -34172
rect 15967 -34198 16583 -33902
rect 16627 -33928 16923 -33902
rect 16627 -34172 16653 -33928
rect 16653 -34172 16897 -33928
rect 16897 -34172 16923 -33928
rect 16627 -34198 16923 -34172
rect 16967 -34198 17583 -33902
rect 17627 -33928 17923 -33902
rect 17627 -34172 17653 -33928
rect 17653 -34172 17897 -33928
rect 17897 -34172 17923 -33928
rect 17627 -34198 17923 -34172
rect 17967 -34198 18583 -33902
rect 18627 -33928 18923 -33902
rect 18627 -34172 18653 -33928
rect 18653 -34172 18897 -33928
rect 18897 -34172 18923 -33928
rect 18627 -34198 18923 -34172
rect 18967 -34198 19583 -33902
rect 19627 -33928 19923 -33902
rect 19627 -34172 19653 -33928
rect 19653 -34172 19897 -33928
rect 19897 -34172 19923 -33928
rect 19627 -34198 19923 -34172
rect 19967 -34198 20583 -33902
rect 20627 -33928 20923 -33902
rect 20627 -34172 20653 -33928
rect 20653 -34172 20897 -33928
rect 20897 -34172 20923 -33928
rect 20627 -34198 20923 -34172
rect 20967 -34198 21583 -33902
rect 21627 -33928 21923 -33902
rect 21627 -34172 21653 -33928
rect 21653 -34172 21897 -33928
rect 21897 -34172 21923 -33928
rect 21627 -34198 21923 -34172
rect 21967 -34198 22583 -33902
rect 22627 -33928 22923 -33902
rect 22627 -34172 22653 -33928
rect 22653 -34172 22897 -33928
rect 22897 -34172 22923 -33928
rect 22627 -34198 22923 -34172
rect 22967 -34198 23583 -33902
rect 23627 -33928 23923 -33902
rect 23627 -34172 23653 -33928
rect 23653 -34172 23897 -33928
rect 23897 -34172 23923 -33928
rect 23627 -34198 23923 -34172
rect 23967 -34198 24583 -33902
rect 24627 -33928 24923 -33902
rect 24627 -34172 24653 -33928
rect 24653 -34172 24897 -33928
rect 24897 -34172 24923 -33928
rect 24627 -34198 24923 -34172
rect 24967 -34198 25583 -33902
rect 25627 -33928 25923 -33902
rect 25627 -34172 25653 -33928
rect 25653 -34172 25897 -33928
rect 25897 -34172 25923 -33928
rect 25627 -34198 25923 -34172
rect 25967 -34198 26583 -33902
rect 26627 -33928 26923 -33902
rect 26627 -34172 26653 -33928
rect 26653 -34172 26897 -33928
rect 26897 -34172 26923 -33928
rect 26627 -34198 26923 -34172
rect 26967 -34198 27583 -33902
rect 27627 -33928 27923 -33902
rect 27627 -34172 27653 -33928
rect 27653 -34172 27897 -33928
rect 27897 -34172 27923 -33928
rect 27627 -34198 27923 -34172
rect 27967 -34198 28583 -33902
rect 28627 -33928 28923 -33902
rect 28627 -34172 28653 -33928
rect 28653 -34172 28897 -33928
rect 28897 -34172 28923 -33928
rect 28627 -34198 28923 -34172
rect 28967 -34198 29583 -33902
rect 29627 -33928 29923 -33902
rect 29627 -34172 29653 -33928
rect 29653 -34172 29897 -33928
rect 29897 -34172 29923 -33928
rect 29627 -34198 29923 -34172
rect 29967 -34198 30583 -33902
rect 30627 -33928 30923 -33902
rect 30627 -34172 30653 -33928
rect 30653 -34172 30897 -33928
rect 30897 -34172 30923 -33928
rect 30627 -34198 30923 -34172
rect 30967 -34198 31583 -33902
rect 31627 -33928 31923 -33902
rect 31627 -34172 31653 -33928
rect 31653 -34172 31897 -33928
rect 31897 -34172 31923 -33928
rect 31627 -34198 31923 -34172
rect 31967 -34198 32583 -33902
rect 32627 -33928 32923 -33902
rect 32627 -34172 32653 -33928
rect 32653 -34172 32897 -33928
rect 32897 -34172 32923 -33928
rect 32627 -34198 32923 -34172
rect 32967 -34198 33583 -33902
rect 33627 -33928 33923 -33902
rect 33627 -34172 33653 -33928
rect 33653 -34172 33897 -33928
rect 33897 -34172 33923 -33928
rect 33627 -34198 33923 -34172
rect 33967 -34198 34263 -33902
rect 8627 -34858 8923 -34242
rect 9627 -34858 9923 -34242
rect 10627 -34858 10923 -34242
rect 11627 -34858 11923 -34242
rect 12627 -34858 12923 -34242
rect 13627 -34858 13923 -34242
rect 14627 -34858 14923 -34242
rect 15627 -34858 15923 -34242
rect 16627 -34858 16923 -34242
rect 17627 -34858 17923 -34242
rect 18627 -34858 18923 -34242
rect 19627 -34858 19923 -34242
rect 20627 -34858 20923 -34242
rect 21627 -34858 21923 -34242
rect 22627 -34858 22923 -34242
rect 23627 -34858 23923 -34242
rect 24627 -34858 24923 -34242
rect 25627 -34858 25923 -34242
rect 26627 -34858 26923 -34242
rect 27627 -34858 27923 -34242
rect 28627 -34858 28923 -34242
rect 29627 -34858 29923 -34242
rect 30627 -34858 30923 -34242
rect 31627 -34858 31923 -34242
rect 32627 -34858 32923 -34242
rect 33627 -34858 33923 -34242
rect 8287 -35198 8583 -34902
rect 8627 -34928 8923 -34902
rect 8627 -35172 8653 -34928
rect 8653 -35172 8897 -34928
rect 8897 -35172 8923 -34928
rect 8627 -35198 8923 -35172
rect 8967 -35198 9583 -34902
rect 9627 -34928 9923 -34902
rect 9627 -35172 9653 -34928
rect 9653 -35172 9897 -34928
rect 9897 -35172 9923 -34928
rect 9627 -35198 9923 -35172
rect 9967 -35198 10583 -34902
rect 10627 -34928 10923 -34902
rect 10627 -35172 10653 -34928
rect 10653 -35172 10897 -34928
rect 10897 -35172 10923 -34928
rect 10627 -35198 10923 -35172
rect 10967 -35198 11583 -34902
rect 11627 -34928 11923 -34902
rect 11627 -35172 11653 -34928
rect 11653 -35172 11897 -34928
rect 11897 -35172 11923 -34928
rect 11627 -35198 11923 -35172
rect 11967 -35198 12583 -34902
rect 12627 -34928 12923 -34902
rect 12627 -35172 12653 -34928
rect 12653 -35172 12897 -34928
rect 12897 -35172 12923 -34928
rect 12627 -35198 12923 -35172
rect 12967 -35198 13583 -34902
rect 13627 -34928 13923 -34902
rect 13627 -35172 13653 -34928
rect 13653 -35172 13897 -34928
rect 13897 -35172 13923 -34928
rect 13627 -35198 13923 -35172
rect 13967 -35198 14583 -34902
rect 14627 -34928 14923 -34902
rect 14627 -35172 14653 -34928
rect 14653 -35172 14897 -34928
rect 14897 -35172 14923 -34928
rect 14627 -35198 14923 -35172
rect 14967 -35198 15583 -34902
rect 15627 -34928 15923 -34902
rect 15627 -35172 15653 -34928
rect 15653 -35172 15897 -34928
rect 15897 -35172 15923 -34928
rect 15627 -35198 15923 -35172
rect 15967 -35198 16583 -34902
rect 16627 -34928 16923 -34902
rect 16627 -35172 16653 -34928
rect 16653 -35172 16897 -34928
rect 16897 -35172 16923 -34928
rect 16627 -35198 16923 -35172
rect 16967 -35198 17583 -34902
rect 17627 -34928 17923 -34902
rect 17627 -35172 17653 -34928
rect 17653 -35172 17897 -34928
rect 17897 -35172 17923 -34928
rect 17627 -35198 17923 -35172
rect 17967 -35198 18583 -34902
rect 18627 -34928 18923 -34902
rect 18627 -35172 18653 -34928
rect 18653 -35172 18897 -34928
rect 18897 -35172 18923 -34928
rect 18627 -35198 18923 -35172
rect 18967 -35198 19583 -34902
rect 19627 -34928 19923 -34902
rect 19627 -35172 19653 -34928
rect 19653 -35172 19897 -34928
rect 19897 -35172 19923 -34928
rect 19627 -35198 19923 -35172
rect 19967 -35198 20583 -34902
rect 20627 -34928 20923 -34902
rect 20627 -35172 20653 -34928
rect 20653 -35172 20897 -34928
rect 20897 -35172 20923 -34928
rect 20627 -35198 20923 -35172
rect 20967 -35198 21583 -34902
rect 21627 -34928 21923 -34902
rect 21627 -35172 21653 -34928
rect 21653 -35172 21897 -34928
rect 21897 -35172 21923 -34928
rect 21627 -35198 21923 -35172
rect 21967 -35198 22583 -34902
rect 22627 -34928 22923 -34902
rect 22627 -35172 22653 -34928
rect 22653 -35172 22897 -34928
rect 22897 -35172 22923 -34928
rect 22627 -35198 22923 -35172
rect 22967 -35198 23583 -34902
rect 23627 -34928 23923 -34902
rect 23627 -35172 23653 -34928
rect 23653 -35172 23897 -34928
rect 23897 -35172 23923 -34928
rect 23627 -35198 23923 -35172
rect 23967 -35198 24583 -34902
rect 24627 -34928 24923 -34902
rect 24627 -35172 24653 -34928
rect 24653 -35172 24897 -34928
rect 24897 -35172 24923 -34928
rect 24627 -35198 24923 -35172
rect 24967 -35198 25583 -34902
rect 25627 -34928 25923 -34902
rect 25627 -35172 25653 -34928
rect 25653 -35172 25897 -34928
rect 25897 -35172 25923 -34928
rect 25627 -35198 25923 -35172
rect 25967 -35198 26583 -34902
rect 26627 -34928 26923 -34902
rect 26627 -35172 26653 -34928
rect 26653 -35172 26897 -34928
rect 26897 -35172 26923 -34928
rect 26627 -35198 26923 -35172
rect 26967 -35198 27583 -34902
rect 27627 -34928 27923 -34902
rect 27627 -35172 27653 -34928
rect 27653 -35172 27897 -34928
rect 27897 -35172 27923 -34928
rect 27627 -35198 27923 -35172
rect 27967 -35198 28583 -34902
rect 28627 -34928 28923 -34902
rect 28627 -35172 28653 -34928
rect 28653 -35172 28897 -34928
rect 28897 -35172 28923 -34928
rect 28627 -35198 28923 -35172
rect 28967 -35198 29583 -34902
rect 29627 -34928 29923 -34902
rect 29627 -35172 29653 -34928
rect 29653 -35172 29897 -34928
rect 29897 -35172 29923 -34928
rect 29627 -35198 29923 -35172
rect 29967 -35198 30583 -34902
rect 30627 -34928 30923 -34902
rect 30627 -35172 30653 -34928
rect 30653 -35172 30897 -34928
rect 30897 -35172 30923 -34928
rect 30627 -35198 30923 -35172
rect 30967 -35198 31583 -34902
rect 31627 -34928 31923 -34902
rect 31627 -35172 31653 -34928
rect 31653 -35172 31897 -34928
rect 31897 -35172 31923 -34928
rect 31627 -35198 31923 -35172
rect 31967 -35198 32583 -34902
rect 32627 -34928 32923 -34902
rect 32627 -35172 32653 -34928
rect 32653 -35172 32897 -34928
rect 32897 -35172 32923 -34928
rect 32627 -35198 32923 -35172
rect 32967 -35198 33583 -34902
rect 33627 -34928 33923 -34902
rect 33627 -35172 33653 -34928
rect 33653 -35172 33897 -34928
rect 33897 -35172 33923 -34928
rect 33627 -35198 33923 -35172
rect 33967 -35198 34263 -34902
rect 8627 -35858 8923 -35242
rect 9627 -35858 9923 -35242
rect 10627 -35858 10923 -35242
rect 11627 -35858 11923 -35242
rect 12627 -35858 12923 -35242
rect 13627 -35858 13923 -35242
rect 14627 -35858 14923 -35242
rect 15627 -35858 15923 -35242
rect 16627 -35858 16923 -35242
rect 17627 -35858 17923 -35242
rect 18627 -35858 18923 -35242
rect 19627 -35858 19923 -35242
rect 20627 -35858 20923 -35242
rect 21627 -35858 21923 -35242
rect 22627 -35858 22923 -35242
rect 23627 -35858 23923 -35242
rect 24627 -35858 24923 -35242
rect 25627 -35858 25923 -35242
rect 26627 -35858 26923 -35242
rect 27627 -35858 27923 -35242
rect 28627 -35858 28923 -35242
rect 29627 -35858 29923 -35242
rect 30627 -35858 30923 -35242
rect 31627 -35858 31923 -35242
rect 32627 -35858 32923 -35242
rect 33627 -35858 33923 -35242
rect 8287 -36198 8583 -35902
rect 8627 -35928 8923 -35902
rect 8627 -36172 8653 -35928
rect 8653 -36172 8897 -35928
rect 8897 -36172 8923 -35928
rect 8627 -36198 8923 -36172
rect 8967 -36198 9583 -35902
rect 9627 -35928 9923 -35902
rect 9627 -36172 9653 -35928
rect 9653 -36172 9897 -35928
rect 9897 -36172 9923 -35928
rect 9627 -36198 9923 -36172
rect 9967 -36198 10583 -35902
rect 10627 -35928 10923 -35902
rect 10627 -36172 10653 -35928
rect 10653 -36172 10897 -35928
rect 10897 -36172 10923 -35928
rect 10627 -36198 10923 -36172
rect 10967 -36198 11583 -35902
rect 11627 -35928 11923 -35902
rect 11627 -36172 11653 -35928
rect 11653 -36172 11897 -35928
rect 11897 -36172 11923 -35928
rect 11627 -36198 11923 -36172
rect 11967 -36198 12583 -35902
rect 12627 -35928 12923 -35902
rect 12627 -36172 12653 -35928
rect 12653 -36172 12897 -35928
rect 12897 -36172 12923 -35928
rect 12627 -36198 12923 -36172
rect 12967 -36198 13583 -35902
rect 13627 -35928 13923 -35902
rect 13627 -36172 13653 -35928
rect 13653 -36172 13897 -35928
rect 13897 -36172 13923 -35928
rect 13627 -36198 13923 -36172
rect 13967 -36198 14583 -35902
rect 14627 -35928 14923 -35902
rect 14627 -36172 14653 -35928
rect 14653 -36172 14897 -35928
rect 14897 -36172 14923 -35928
rect 14627 -36198 14923 -36172
rect 14967 -36198 15583 -35902
rect 15627 -35928 15923 -35902
rect 15627 -36172 15653 -35928
rect 15653 -36172 15897 -35928
rect 15897 -36172 15923 -35928
rect 15627 -36198 15923 -36172
rect 15967 -36198 16583 -35902
rect 16627 -35928 16923 -35902
rect 16627 -36172 16653 -35928
rect 16653 -36172 16897 -35928
rect 16897 -36172 16923 -35928
rect 16627 -36198 16923 -36172
rect 16967 -36198 17583 -35902
rect 17627 -35928 17923 -35902
rect 17627 -36172 17653 -35928
rect 17653 -36172 17897 -35928
rect 17897 -36172 17923 -35928
rect 17627 -36198 17923 -36172
rect 17967 -36198 18583 -35902
rect 18627 -35928 18923 -35902
rect 18627 -36172 18653 -35928
rect 18653 -36172 18897 -35928
rect 18897 -36172 18923 -35928
rect 18627 -36198 18923 -36172
rect 18967 -36198 19583 -35902
rect 19627 -35928 19923 -35902
rect 19627 -36172 19653 -35928
rect 19653 -36172 19897 -35928
rect 19897 -36172 19923 -35928
rect 19627 -36198 19923 -36172
rect 19967 -36198 20583 -35902
rect 20627 -35928 20923 -35902
rect 20627 -36172 20653 -35928
rect 20653 -36172 20897 -35928
rect 20897 -36172 20923 -35928
rect 20627 -36198 20923 -36172
rect 20967 -36198 21583 -35902
rect 21627 -35928 21923 -35902
rect 21627 -36172 21653 -35928
rect 21653 -36172 21897 -35928
rect 21897 -36172 21923 -35928
rect 21627 -36198 21923 -36172
rect 21967 -36198 22583 -35902
rect 22627 -35928 22923 -35902
rect 22627 -36172 22653 -35928
rect 22653 -36172 22897 -35928
rect 22897 -36172 22923 -35928
rect 22627 -36198 22923 -36172
rect 22967 -36198 23583 -35902
rect 23627 -35928 23923 -35902
rect 23627 -36172 23653 -35928
rect 23653 -36172 23897 -35928
rect 23897 -36172 23923 -35928
rect 23627 -36198 23923 -36172
rect 23967 -36198 24583 -35902
rect 24627 -35928 24923 -35902
rect 24627 -36172 24653 -35928
rect 24653 -36172 24897 -35928
rect 24897 -36172 24923 -35928
rect 24627 -36198 24923 -36172
rect 24967 -36198 25583 -35902
rect 25627 -35928 25923 -35902
rect 25627 -36172 25653 -35928
rect 25653 -36172 25897 -35928
rect 25897 -36172 25923 -35928
rect 25627 -36198 25923 -36172
rect 25967 -36198 26583 -35902
rect 26627 -35928 26923 -35902
rect 26627 -36172 26653 -35928
rect 26653 -36172 26897 -35928
rect 26897 -36172 26923 -35928
rect 26627 -36198 26923 -36172
rect 26967 -36198 27583 -35902
rect 27627 -35928 27923 -35902
rect 27627 -36172 27653 -35928
rect 27653 -36172 27897 -35928
rect 27897 -36172 27923 -35928
rect 27627 -36198 27923 -36172
rect 27967 -36198 28583 -35902
rect 28627 -35928 28923 -35902
rect 28627 -36172 28653 -35928
rect 28653 -36172 28897 -35928
rect 28897 -36172 28923 -35928
rect 28627 -36198 28923 -36172
rect 28967 -36198 29583 -35902
rect 29627 -35928 29923 -35902
rect 29627 -36172 29653 -35928
rect 29653 -36172 29897 -35928
rect 29897 -36172 29923 -35928
rect 29627 -36198 29923 -36172
rect 29967 -36198 30583 -35902
rect 30627 -35928 30923 -35902
rect 30627 -36172 30653 -35928
rect 30653 -36172 30897 -35928
rect 30897 -36172 30923 -35928
rect 30627 -36198 30923 -36172
rect 30967 -36198 31583 -35902
rect 31627 -35928 31923 -35902
rect 31627 -36172 31653 -35928
rect 31653 -36172 31897 -35928
rect 31897 -36172 31923 -35928
rect 31627 -36198 31923 -36172
rect 31967 -36198 32583 -35902
rect 32627 -35928 32923 -35902
rect 32627 -36172 32653 -35928
rect 32653 -36172 32897 -35928
rect 32897 -36172 32923 -35928
rect 32627 -36198 32923 -36172
rect 32967 -36198 33583 -35902
rect 33627 -35928 33923 -35902
rect 33627 -36172 33653 -35928
rect 33653 -36172 33897 -35928
rect 33897 -36172 33923 -35928
rect 33627 -36198 33923 -36172
rect 33967 -36198 34263 -35902
rect 8627 -36858 8923 -36242
rect 9627 -36858 9923 -36242
rect 10627 -36858 10923 -36242
rect 11627 -36858 11923 -36242
rect 12627 -36858 12923 -36242
rect 13627 -36858 13923 -36242
rect 14627 -36858 14923 -36242
rect 15627 -36858 15923 -36242
rect 16627 -36858 16923 -36242
rect 17627 -36858 17923 -36242
rect 18627 -36858 18923 -36242
rect 19627 -36858 19923 -36242
rect 20627 -36858 20923 -36242
rect 21627 -36858 21923 -36242
rect 22627 -36858 22923 -36242
rect 23627 -36858 23923 -36242
rect 24627 -36858 24923 -36242
rect 25627 -36858 25923 -36242
rect 26627 -36858 26923 -36242
rect 27627 -36858 27923 -36242
rect 28627 -36858 28923 -36242
rect 29627 -36858 29923 -36242
rect 30627 -36858 30923 -36242
rect 31627 -36858 31923 -36242
rect 32627 -36858 32923 -36242
rect 33627 -36858 33923 -36242
rect 8287 -37198 8583 -36902
rect 8627 -36928 8923 -36902
rect 8627 -37172 8653 -36928
rect 8653 -37172 8897 -36928
rect 8897 -37172 8923 -36928
rect 8627 -37198 8923 -37172
rect 8967 -37198 9583 -36902
rect 9627 -36928 9923 -36902
rect 9627 -37172 9653 -36928
rect 9653 -37172 9897 -36928
rect 9897 -37172 9923 -36928
rect 9627 -37198 9923 -37172
rect 9967 -37198 10583 -36902
rect 10627 -36928 10923 -36902
rect 10627 -37172 10653 -36928
rect 10653 -37172 10897 -36928
rect 10897 -37172 10923 -36928
rect 10627 -37198 10923 -37172
rect 10967 -37198 11583 -36902
rect 11627 -36928 11923 -36902
rect 11627 -37172 11653 -36928
rect 11653 -37172 11897 -36928
rect 11897 -37172 11923 -36928
rect 11627 -37198 11923 -37172
rect 11967 -37198 12583 -36902
rect 12627 -36928 12923 -36902
rect 12627 -37172 12653 -36928
rect 12653 -37172 12897 -36928
rect 12897 -37172 12923 -36928
rect 12627 -37198 12923 -37172
rect 12967 -37198 13583 -36902
rect 13627 -36928 13923 -36902
rect 13627 -37172 13653 -36928
rect 13653 -37172 13897 -36928
rect 13897 -37172 13923 -36928
rect 13627 -37198 13923 -37172
rect 13967 -37198 14583 -36902
rect 14627 -36928 14923 -36902
rect 14627 -37172 14653 -36928
rect 14653 -37172 14897 -36928
rect 14897 -37172 14923 -36928
rect 14627 -37198 14923 -37172
rect 14967 -37198 15583 -36902
rect 15627 -36928 15923 -36902
rect 15627 -37172 15653 -36928
rect 15653 -37172 15897 -36928
rect 15897 -37172 15923 -36928
rect 15627 -37198 15923 -37172
rect 15967 -37198 16583 -36902
rect 16627 -36928 16923 -36902
rect 16627 -37172 16653 -36928
rect 16653 -37172 16897 -36928
rect 16897 -37172 16923 -36928
rect 16627 -37198 16923 -37172
rect 16967 -37198 17583 -36902
rect 17627 -36928 17923 -36902
rect 17627 -37172 17653 -36928
rect 17653 -37172 17897 -36928
rect 17897 -37172 17923 -36928
rect 17627 -37198 17923 -37172
rect 17967 -37198 18583 -36902
rect 18627 -36928 18923 -36902
rect 18627 -37172 18653 -36928
rect 18653 -37172 18897 -36928
rect 18897 -37172 18923 -36928
rect 18627 -37198 18923 -37172
rect 18967 -37198 19583 -36902
rect 19627 -36928 19923 -36902
rect 19627 -37172 19653 -36928
rect 19653 -37172 19897 -36928
rect 19897 -37172 19923 -36928
rect 19627 -37198 19923 -37172
rect 19967 -37198 20583 -36902
rect 20627 -36928 20923 -36902
rect 20627 -37172 20653 -36928
rect 20653 -37172 20897 -36928
rect 20897 -37172 20923 -36928
rect 20627 -37198 20923 -37172
rect 20967 -37198 21583 -36902
rect 21627 -36928 21923 -36902
rect 21627 -37172 21653 -36928
rect 21653 -37172 21897 -36928
rect 21897 -37172 21923 -36928
rect 21627 -37198 21923 -37172
rect 21967 -37198 22583 -36902
rect 22627 -36928 22923 -36902
rect 22627 -37172 22653 -36928
rect 22653 -37172 22897 -36928
rect 22897 -37172 22923 -36928
rect 22627 -37198 22923 -37172
rect 22967 -37198 23583 -36902
rect 23627 -36928 23923 -36902
rect 23627 -37172 23653 -36928
rect 23653 -37172 23897 -36928
rect 23897 -37172 23923 -36928
rect 23627 -37198 23923 -37172
rect 23967 -37198 24583 -36902
rect 24627 -36928 24923 -36902
rect 24627 -37172 24653 -36928
rect 24653 -37172 24897 -36928
rect 24897 -37172 24923 -36928
rect 24627 -37198 24923 -37172
rect 24967 -37198 25583 -36902
rect 25627 -36928 25923 -36902
rect 25627 -37172 25653 -36928
rect 25653 -37172 25897 -36928
rect 25897 -37172 25923 -36928
rect 25627 -37198 25923 -37172
rect 25967 -37198 26583 -36902
rect 26627 -36928 26923 -36902
rect 26627 -37172 26653 -36928
rect 26653 -37172 26897 -36928
rect 26897 -37172 26923 -36928
rect 26627 -37198 26923 -37172
rect 26967 -37198 27583 -36902
rect 27627 -36928 27923 -36902
rect 27627 -37172 27653 -36928
rect 27653 -37172 27897 -36928
rect 27897 -37172 27923 -36928
rect 27627 -37198 27923 -37172
rect 27967 -37198 28583 -36902
rect 28627 -36928 28923 -36902
rect 28627 -37172 28653 -36928
rect 28653 -37172 28897 -36928
rect 28897 -37172 28923 -36928
rect 28627 -37198 28923 -37172
rect 28967 -37198 29583 -36902
rect 29627 -36928 29923 -36902
rect 29627 -37172 29653 -36928
rect 29653 -37172 29897 -36928
rect 29897 -37172 29923 -36928
rect 29627 -37198 29923 -37172
rect 29967 -37198 30583 -36902
rect 30627 -36928 30923 -36902
rect 30627 -37172 30653 -36928
rect 30653 -37172 30897 -36928
rect 30897 -37172 30923 -36928
rect 30627 -37198 30923 -37172
rect 30967 -37198 31583 -36902
rect 31627 -36928 31923 -36902
rect 31627 -37172 31653 -36928
rect 31653 -37172 31897 -36928
rect 31897 -37172 31923 -36928
rect 31627 -37198 31923 -37172
rect 31967 -37198 32583 -36902
rect 32627 -36928 32923 -36902
rect 32627 -37172 32653 -36928
rect 32653 -37172 32897 -36928
rect 32897 -37172 32923 -36928
rect 32627 -37198 32923 -37172
rect 32967 -37198 33583 -36902
rect 33627 -36928 33923 -36902
rect 33627 -37172 33653 -36928
rect 33653 -37172 33897 -36928
rect 33897 -37172 33923 -36928
rect 33627 -37198 33923 -37172
rect 33967 -37198 34263 -36902
rect 8627 -37858 8923 -37242
rect 9627 -37858 9923 -37242
rect 10627 -37858 10923 -37242
rect 11627 -37858 11923 -37242
rect 12627 -37858 12923 -37242
rect 13627 -37858 13923 -37242
rect 14627 -37858 14923 -37242
rect 15627 -37858 15923 -37242
rect 16627 -37858 16923 -37242
rect 17627 -37858 17923 -37242
rect 18627 -37858 18923 -37242
rect 19627 -37858 19923 -37242
rect 20627 -37858 20923 -37242
rect 21627 -37858 21923 -37242
rect 22627 -37858 22923 -37242
rect 23627 -37858 23923 -37242
rect 24627 -37858 24923 -37242
rect 25627 -37858 25923 -37242
rect 26627 -37858 26923 -37242
rect 27627 -37858 27923 -37242
rect 28627 -37858 28923 -37242
rect 29627 -37858 29923 -37242
rect 30627 -37858 30923 -37242
rect 31627 -37858 31923 -37242
rect 32627 -37858 32923 -37242
rect 33627 -37858 33923 -37242
rect 8287 -38198 8583 -37902
rect 8627 -37928 8923 -37902
rect 8627 -38172 8653 -37928
rect 8653 -38172 8897 -37928
rect 8897 -38172 8923 -37928
rect 8627 -38198 8923 -38172
rect 8967 -38198 9583 -37902
rect 9627 -37928 9923 -37902
rect 9627 -38172 9653 -37928
rect 9653 -38172 9897 -37928
rect 9897 -38172 9923 -37928
rect 9627 -38198 9923 -38172
rect 9967 -38198 10583 -37902
rect 10627 -37928 10923 -37902
rect 10627 -38172 10653 -37928
rect 10653 -38172 10897 -37928
rect 10897 -38172 10923 -37928
rect 10627 -38198 10923 -38172
rect 10967 -38198 11583 -37902
rect 11627 -37928 11923 -37902
rect 11627 -38172 11653 -37928
rect 11653 -38172 11897 -37928
rect 11897 -38172 11923 -37928
rect 11627 -38198 11923 -38172
rect 11967 -38198 12583 -37902
rect 12627 -37928 12923 -37902
rect 12627 -38172 12653 -37928
rect 12653 -38172 12897 -37928
rect 12897 -38172 12923 -37928
rect 12627 -38198 12923 -38172
rect 12967 -38198 13583 -37902
rect 13627 -37928 13923 -37902
rect 13627 -38172 13653 -37928
rect 13653 -38172 13897 -37928
rect 13897 -38172 13923 -37928
rect 13627 -38198 13923 -38172
rect 13967 -38198 14583 -37902
rect 14627 -37928 14923 -37902
rect 14627 -38172 14653 -37928
rect 14653 -38172 14897 -37928
rect 14897 -38172 14923 -37928
rect 14627 -38198 14923 -38172
rect 14967 -38198 15583 -37902
rect 15627 -37928 15923 -37902
rect 15627 -38172 15653 -37928
rect 15653 -38172 15897 -37928
rect 15897 -38172 15923 -37928
rect 15627 -38198 15923 -38172
rect 15967 -38198 16583 -37902
rect 16627 -37928 16923 -37902
rect 16627 -38172 16653 -37928
rect 16653 -38172 16897 -37928
rect 16897 -38172 16923 -37928
rect 16627 -38198 16923 -38172
rect 16967 -38198 17583 -37902
rect 17627 -37928 17923 -37902
rect 17627 -38172 17653 -37928
rect 17653 -38172 17897 -37928
rect 17897 -38172 17923 -37928
rect 17627 -38198 17923 -38172
rect 17967 -38198 18583 -37902
rect 18627 -37928 18923 -37902
rect 18627 -38172 18653 -37928
rect 18653 -38172 18897 -37928
rect 18897 -38172 18923 -37928
rect 18627 -38198 18923 -38172
rect 18967 -38198 19583 -37902
rect 19627 -37928 19923 -37902
rect 19627 -38172 19653 -37928
rect 19653 -38172 19897 -37928
rect 19897 -38172 19923 -37928
rect 19627 -38198 19923 -38172
rect 19967 -38198 20583 -37902
rect 20627 -37928 20923 -37902
rect 20627 -38172 20653 -37928
rect 20653 -38172 20897 -37928
rect 20897 -38172 20923 -37928
rect 20627 -38198 20923 -38172
rect 20967 -38198 21583 -37902
rect 21627 -37928 21923 -37902
rect 21627 -38172 21653 -37928
rect 21653 -38172 21897 -37928
rect 21897 -38172 21923 -37928
rect 21627 -38198 21923 -38172
rect 21967 -38198 22583 -37902
rect 22627 -37928 22923 -37902
rect 22627 -38172 22653 -37928
rect 22653 -38172 22897 -37928
rect 22897 -38172 22923 -37928
rect 22627 -38198 22923 -38172
rect 22967 -38198 23583 -37902
rect 23627 -37928 23923 -37902
rect 23627 -38172 23653 -37928
rect 23653 -38172 23897 -37928
rect 23897 -38172 23923 -37928
rect 23627 -38198 23923 -38172
rect 23967 -38198 24583 -37902
rect 24627 -37928 24923 -37902
rect 24627 -38172 24653 -37928
rect 24653 -38172 24897 -37928
rect 24897 -38172 24923 -37928
rect 24627 -38198 24923 -38172
rect 24967 -38198 25583 -37902
rect 25627 -37928 25923 -37902
rect 25627 -38172 25653 -37928
rect 25653 -38172 25897 -37928
rect 25897 -38172 25923 -37928
rect 25627 -38198 25923 -38172
rect 25967 -38198 26583 -37902
rect 26627 -37928 26923 -37902
rect 26627 -38172 26653 -37928
rect 26653 -38172 26897 -37928
rect 26897 -38172 26923 -37928
rect 26627 -38198 26923 -38172
rect 26967 -38198 27583 -37902
rect 27627 -37928 27923 -37902
rect 27627 -38172 27653 -37928
rect 27653 -38172 27897 -37928
rect 27897 -38172 27923 -37928
rect 27627 -38198 27923 -38172
rect 27967 -38198 28583 -37902
rect 28627 -37928 28923 -37902
rect 28627 -38172 28653 -37928
rect 28653 -38172 28897 -37928
rect 28897 -38172 28923 -37928
rect 28627 -38198 28923 -38172
rect 28967 -38198 29583 -37902
rect 29627 -37928 29923 -37902
rect 29627 -38172 29653 -37928
rect 29653 -38172 29897 -37928
rect 29897 -38172 29923 -37928
rect 29627 -38198 29923 -38172
rect 29967 -38198 30583 -37902
rect 30627 -37928 30923 -37902
rect 30627 -38172 30653 -37928
rect 30653 -38172 30897 -37928
rect 30897 -38172 30923 -37928
rect 30627 -38198 30923 -38172
rect 30967 -38198 31583 -37902
rect 31627 -37928 31923 -37902
rect 31627 -38172 31653 -37928
rect 31653 -38172 31897 -37928
rect 31897 -38172 31923 -37928
rect 31627 -38198 31923 -38172
rect 31967 -38198 32583 -37902
rect 32627 -37928 32923 -37902
rect 32627 -38172 32653 -37928
rect 32653 -38172 32897 -37928
rect 32897 -38172 32923 -37928
rect 32627 -38198 32923 -38172
rect 32967 -38198 33583 -37902
rect 33627 -37928 33923 -37902
rect 33627 -38172 33653 -37928
rect 33653 -38172 33897 -37928
rect 33897 -38172 33923 -37928
rect 33627 -38198 33923 -38172
rect 33967 -38198 34263 -37902
rect 8627 -38858 8923 -38242
rect 9627 -38858 9923 -38242
rect 10627 -38858 10923 -38242
rect 11627 -38858 11923 -38242
rect 12627 -38858 12923 -38242
rect 13627 -38858 13923 -38242
rect 14627 -38858 14923 -38242
rect 15627 -38858 15923 -38242
rect 16627 -38858 16923 -38242
rect 17627 -38858 17923 -38242
rect 18627 -38858 18923 -38242
rect 19627 -38858 19923 -38242
rect 20627 -38858 20923 -38242
rect 21627 -38858 21923 -38242
rect 22627 -38858 22923 -38242
rect 23627 -38858 23923 -38242
rect 24627 -38858 24923 -38242
rect 25627 -38858 25923 -38242
rect 26627 -38858 26923 -38242
rect 27627 -38858 27923 -38242
rect 28627 -38858 28923 -38242
rect 29627 -38858 29923 -38242
rect 30627 -38858 30923 -38242
rect 31627 -38858 31923 -38242
rect 32627 -38858 32923 -38242
rect 33627 -38858 33923 -38242
rect 8287 -39198 8583 -38902
rect 8627 -38928 8923 -38902
rect 8627 -39172 8653 -38928
rect 8653 -39172 8897 -38928
rect 8897 -39172 8923 -38928
rect 8627 -39198 8923 -39172
rect 8967 -39198 9583 -38902
rect 9627 -38928 9923 -38902
rect 9627 -39172 9653 -38928
rect 9653 -39172 9897 -38928
rect 9897 -39172 9923 -38928
rect 9627 -39198 9923 -39172
rect 9967 -39198 10583 -38902
rect 10627 -38928 10923 -38902
rect 10627 -39172 10653 -38928
rect 10653 -39172 10897 -38928
rect 10897 -39172 10923 -38928
rect 10627 -39198 10923 -39172
rect 10967 -39198 11583 -38902
rect 11627 -38928 11923 -38902
rect 11627 -39172 11653 -38928
rect 11653 -39172 11897 -38928
rect 11897 -39172 11923 -38928
rect 11627 -39198 11923 -39172
rect 11967 -39198 12583 -38902
rect 12627 -38928 12923 -38902
rect 12627 -39172 12653 -38928
rect 12653 -39172 12897 -38928
rect 12897 -39172 12923 -38928
rect 12627 -39198 12923 -39172
rect 12967 -39198 13583 -38902
rect 13627 -38928 13923 -38902
rect 13627 -39172 13653 -38928
rect 13653 -39172 13897 -38928
rect 13897 -39172 13923 -38928
rect 13627 -39198 13923 -39172
rect 13967 -39198 14583 -38902
rect 14627 -38928 14923 -38902
rect 14627 -39172 14653 -38928
rect 14653 -39172 14897 -38928
rect 14897 -39172 14923 -38928
rect 14627 -39198 14923 -39172
rect 14967 -39198 15583 -38902
rect 15627 -38928 15923 -38902
rect 15627 -39172 15653 -38928
rect 15653 -39172 15897 -38928
rect 15897 -39172 15923 -38928
rect 15627 -39198 15923 -39172
rect 15967 -39198 16583 -38902
rect 16627 -38928 16923 -38902
rect 16627 -39172 16653 -38928
rect 16653 -39172 16897 -38928
rect 16897 -39172 16923 -38928
rect 16627 -39198 16923 -39172
rect 16967 -39198 17583 -38902
rect 17627 -38928 17923 -38902
rect 17627 -39172 17653 -38928
rect 17653 -39172 17897 -38928
rect 17897 -39172 17923 -38928
rect 17627 -39198 17923 -39172
rect 17967 -39198 18583 -38902
rect 18627 -38928 18923 -38902
rect 18627 -39172 18653 -38928
rect 18653 -39172 18897 -38928
rect 18897 -39172 18923 -38928
rect 18627 -39198 18923 -39172
rect 18967 -39198 19583 -38902
rect 19627 -38928 19923 -38902
rect 19627 -39172 19653 -38928
rect 19653 -39172 19897 -38928
rect 19897 -39172 19923 -38928
rect 19627 -39198 19923 -39172
rect 19967 -39198 20583 -38902
rect 20627 -38928 20923 -38902
rect 20627 -39172 20653 -38928
rect 20653 -39172 20897 -38928
rect 20897 -39172 20923 -38928
rect 20627 -39198 20923 -39172
rect 20967 -39198 21583 -38902
rect 21627 -38928 21923 -38902
rect 21627 -39172 21653 -38928
rect 21653 -39172 21897 -38928
rect 21897 -39172 21923 -38928
rect 21627 -39198 21923 -39172
rect 21967 -39198 22583 -38902
rect 22627 -38928 22923 -38902
rect 22627 -39172 22653 -38928
rect 22653 -39172 22897 -38928
rect 22897 -39172 22923 -38928
rect 22627 -39198 22923 -39172
rect 22967 -39198 23583 -38902
rect 23627 -38928 23923 -38902
rect 23627 -39172 23653 -38928
rect 23653 -39172 23897 -38928
rect 23897 -39172 23923 -38928
rect 23627 -39198 23923 -39172
rect 23967 -39198 24583 -38902
rect 24627 -38928 24923 -38902
rect 24627 -39172 24653 -38928
rect 24653 -39172 24897 -38928
rect 24897 -39172 24923 -38928
rect 24627 -39198 24923 -39172
rect 24967 -39198 25583 -38902
rect 25627 -38928 25923 -38902
rect 25627 -39172 25653 -38928
rect 25653 -39172 25897 -38928
rect 25897 -39172 25923 -38928
rect 25627 -39198 25923 -39172
rect 25967 -39198 26583 -38902
rect 26627 -38928 26923 -38902
rect 26627 -39172 26653 -38928
rect 26653 -39172 26897 -38928
rect 26897 -39172 26923 -38928
rect 26627 -39198 26923 -39172
rect 26967 -39198 27583 -38902
rect 27627 -38928 27923 -38902
rect 27627 -39172 27653 -38928
rect 27653 -39172 27897 -38928
rect 27897 -39172 27923 -38928
rect 27627 -39198 27923 -39172
rect 27967 -39198 28583 -38902
rect 28627 -38928 28923 -38902
rect 28627 -39172 28653 -38928
rect 28653 -39172 28897 -38928
rect 28897 -39172 28923 -38928
rect 28627 -39198 28923 -39172
rect 28967 -39198 29583 -38902
rect 29627 -38928 29923 -38902
rect 29627 -39172 29653 -38928
rect 29653 -39172 29897 -38928
rect 29897 -39172 29923 -38928
rect 29627 -39198 29923 -39172
rect 29967 -39198 30583 -38902
rect 30627 -38928 30923 -38902
rect 30627 -39172 30653 -38928
rect 30653 -39172 30897 -38928
rect 30897 -39172 30923 -38928
rect 30627 -39198 30923 -39172
rect 30967 -39198 31583 -38902
rect 31627 -38928 31923 -38902
rect 31627 -39172 31653 -38928
rect 31653 -39172 31897 -38928
rect 31897 -39172 31923 -38928
rect 31627 -39198 31923 -39172
rect 31967 -39198 32583 -38902
rect 32627 -38928 32923 -38902
rect 32627 -39172 32653 -38928
rect 32653 -39172 32897 -38928
rect 32897 -39172 32923 -38928
rect 32627 -39198 32923 -39172
rect 32967 -39198 33583 -38902
rect 33627 -38928 33923 -38902
rect 33627 -39172 33653 -38928
rect 33653 -39172 33897 -38928
rect 33897 -39172 33923 -38928
rect 33627 -39198 33923 -39172
rect 33967 -39198 34263 -38902
rect 8627 -39858 8923 -39242
rect 9627 -39858 9923 -39242
rect 10627 -39858 10923 -39242
rect 11627 -39858 11923 -39242
rect 12627 -39858 12923 -39242
rect 13627 -39858 13923 -39242
rect 14627 -39858 14923 -39242
rect 15627 -39858 15923 -39242
rect 16627 -39858 16923 -39242
rect 17627 -39858 17923 -39242
rect 18627 -39858 18923 -39242
rect 19627 -39858 19923 -39242
rect 20627 -39858 20923 -39242
rect 21627 -39858 21923 -39242
rect 22627 -39858 22923 -39242
rect 23627 -39858 23923 -39242
rect 24627 -39858 24923 -39242
rect 25627 -39858 25923 -39242
rect 26627 -39858 26923 -39242
rect 27627 -39858 27923 -39242
rect 28627 -39858 28923 -39242
rect 29627 -39858 29923 -39242
rect 30627 -39858 30923 -39242
rect 31627 -39858 31923 -39242
rect 32627 -39858 32923 -39242
rect 33627 -39858 33923 -39242
rect 8287 -40198 8583 -39902
rect 8627 -39928 8923 -39902
rect 8627 -40172 8653 -39928
rect 8653 -40172 8897 -39928
rect 8897 -40172 8923 -39928
rect 8627 -40198 8923 -40172
rect 8967 -40198 9583 -39902
rect 9627 -39928 9923 -39902
rect 9627 -40172 9653 -39928
rect 9653 -40172 9897 -39928
rect 9897 -40172 9923 -39928
rect 9627 -40198 9923 -40172
rect 9967 -40198 10583 -39902
rect 10627 -39928 10923 -39902
rect 10627 -40172 10653 -39928
rect 10653 -40172 10897 -39928
rect 10897 -40172 10923 -39928
rect 10627 -40198 10923 -40172
rect 10967 -40198 11583 -39902
rect 11627 -39928 11923 -39902
rect 11627 -40172 11653 -39928
rect 11653 -40172 11897 -39928
rect 11897 -40172 11923 -39928
rect 11627 -40198 11923 -40172
rect 11967 -40198 12583 -39902
rect 12627 -39928 12923 -39902
rect 12627 -40172 12653 -39928
rect 12653 -40172 12897 -39928
rect 12897 -40172 12923 -39928
rect 12627 -40198 12923 -40172
rect 12967 -40198 13583 -39902
rect 13627 -39928 13923 -39902
rect 13627 -40172 13653 -39928
rect 13653 -40172 13897 -39928
rect 13897 -40172 13923 -39928
rect 13627 -40198 13923 -40172
rect 13967 -40198 14583 -39902
rect 14627 -39928 14923 -39902
rect 14627 -40172 14653 -39928
rect 14653 -40172 14897 -39928
rect 14897 -40172 14923 -39928
rect 14627 -40198 14923 -40172
rect 14967 -40198 15583 -39902
rect 15627 -39928 15923 -39902
rect 15627 -40172 15653 -39928
rect 15653 -40172 15897 -39928
rect 15897 -40172 15923 -39928
rect 15627 -40198 15923 -40172
rect 15967 -40198 16583 -39902
rect 16627 -39928 16923 -39902
rect 16627 -40172 16653 -39928
rect 16653 -40172 16897 -39928
rect 16897 -40172 16923 -39928
rect 16627 -40198 16923 -40172
rect 16967 -40198 17583 -39902
rect 17627 -39928 17923 -39902
rect 17627 -40172 17653 -39928
rect 17653 -40172 17897 -39928
rect 17897 -40172 17923 -39928
rect 17627 -40198 17923 -40172
rect 17967 -40198 18583 -39902
rect 18627 -39928 18923 -39902
rect 18627 -40172 18653 -39928
rect 18653 -40172 18897 -39928
rect 18897 -40172 18923 -39928
rect 18627 -40198 18923 -40172
rect 18967 -40198 19583 -39902
rect 19627 -39928 19923 -39902
rect 19627 -40172 19653 -39928
rect 19653 -40172 19897 -39928
rect 19897 -40172 19923 -39928
rect 19627 -40198 19923 -40172
rect 19967 -40198 20583 -39902
rect 20627 -39928 20923 -39902
rect 20627 -40172 20653 -39928
rect 20653 -40172 20897 -39928
rect 20897 -40172 20923 -39928
rect 20627 -40198 20923 -40172
rect 20967 -40198 21583 -39902
rect 21627 -39928 21923 -39902
rect 21627 -40172 21653 -39928
rect 21653 -40172 21897 -39928
rect 21897 -40172 21923 -39928
rect 21627 -40198 21923 -40172
rect 21967 -40198 22583 -39902
rect 22627 -39928 22923 -39902
rect 22627 -40172 22653 -39928
rect 22653 -40172 22897 -39928
rect 22897 -40172 22923 -39928
rect 22627 -40198 22923 -40172
rect 22967 -40198 23583 -39902
rect 23627 -39928 23923 -39902
rect 23627 -40172 23653 -39928
rect 23653 -40172 23897 -39928
rect 23897 -40172 23923 -39928
rect 23627 -40198 23923 -40172
rect 23967 -40198 24583 -39902
rect 24627 -39928 24923 -39902
rect 24627 -40172 24653 -39928
rect 24653 -40172 24897 -39928
rect 24897 -40172 24923 -39928
rect 24627 -40198 24923 -40172
rect 24967 -40198 25583 -39902
rect 25627 -39928 25923 -39902
rect 25627 -40172 25653 -39928
rect 25653 -40172 25897 -39928
rect 25897 -40172 25923 -39928
rect 25627 -40198 25923 -40172
rect 25967 -40198 26583 -39902
rect 26627 -39928 26923 -39902
rect 26627 -40172 26653 -39928
rect 26653 -40172 26897 -39928
rect 26897 -40172 26923 -39928
rect 26627 -40198 26923 -40172
rect 26967 -40198 27583 -39902
rect 27627 -39928 27923 -39902
rect 27627 -40172 27653 -39928
rect 27653 -40172 27897 -39928
rect 27897 -40172 27923 -39928
rect 27627 -40198 27923 -40172
rect 27967 -40198 28583 -39902
rect 28627 -39928 28923 -39902
rect 28627 -40172 28653 -39928
rect 28653 -40172 28897 -39928
rect 28897 -40172 28923 -39928
rect 28627 -40198 28923 -40172
rect 28967 -40198 29583 -39902
rect 29627 -39928 29923 -39902
rect 29627 -40172 29653 -39928
rect 29653 -40172 29897 -39928
rect 29897 -40172 29923 -39928
rect 29627 -40198 29923 -40172
rect 29967 -40198 30583 -39902
rect 30627 -39928 30923 -39902
rect 30627 -40172 30653 -39928
rect 30653 -40172 30897 -39928
rect 30897 -40172 30923 -39928
rect 30627 -40198 30923 -40172
rect 30967 -40198 31583 -39902
rect 31627 -39928 31923 -39902
rect 31627 -40172 31653 -39928
rect 31653 -40172 31897 -39928
rect 31897 -40172 31923 -39928
rect 31627 -40198 31923 -40172
rect 31967 -40198 32583 -39902
rect 32627 -39928 32923 -39902
rect 32627 -40172 32653 -39928
rect 32653 -40172 32897 -39928
rect 32897 -40172 32923 -39928
rect 32627 -40198 32923 -40172
rect 32967 -40198 33583 -39902
rect 33627 -39928 33923 -39902
rect 33627 -40172 33653 -39928
rect 33653 -40172 33897 -39928
rect 33897 -40172 33923 -39928
rect 33627 -40198 33923 -40172
rect 33967 -40198 34263 -39902
rect 8627 -40858 8923 -40242
rect 9627 -40858 9923 -40242
rect 10627 -40858 10923 -40242
rect 11627 -40858 11923 -40242
rect 12627 -40858 12923 -40242
rect 13627 -40858 13923 -40242
rect 14627 -40858 14923 -40242
rect 15627 -40858 15923 -40242
rect 16627 -40858 16923 -40242
rect 17627 -40858 17923 -40242
rect 18627 -40858 18923 -40242
rect 19627 -40858 19923 -40242
rect 20627 -40858 20923 -40242
rect 21627 -40858 21923 -40242
rect 22627 -40858 22923 -40242
rect 23627 -40858 23923 -40242
rect 24627 -40858 24923 -40242
rect 25627 -40858 25923 -40242
rect 26627 -40858 26923 -40242
rect 27627 -40858 27923 -40242
rect 28627 -40858 28923 -40242
rect 29627 -40858 29923 -40242
rect 30627 -40858 30923 -40242
rect 31627 -40858 31923 -40242
rect 32627 -40858 32923 -40242
rect 33627 -40858 33923 -40242
rect 8287 -41198 8583 -40902
rect 8627 -40928 8923 -40902
rect 8627 -41172 8653 -40928
rect 8653 -41172 8897 -40928
rect 8897 -41172 8923 -40928
rect 8627 -41198 8923 -41172
rect 8967 -41198 9583 -40902
rect 9627 -40928 9923 -40902
rect 9627 -41172 9653 -40928
rect 9653 -41172 9897 -40928
rect 9897 -41172 9923 -40928
rect 9627 -41198 9923 -41172
rect 9967 -41198 10583 -40902
rect 10627 -40928 10923 -40902
rect 10627 -41172 10653 -40928
rect 10653 -41172 10897 -40928
rect 10897 -41172 10923 -40928
rect 10627 -41198 10923 -41172
rect 10967 -41198 11583 -40902
rect 11627 -40928 11923 -40902
rect 11627 -41172 11653 -40928
rect 11653 -41172 11897 -40928
rect 11897 -41172 11923 -40928
rect 11627 -41198 11923 -41172
rect 11967 -41198 12583 -40902
rect 12627 -40928 12923 -40902
rect 12627 -41172 12653 -40928
rect 12653 -41172 12897 -40928
rect 12897 -41172 12923 -40928
rect 12627 -41198 12923 -41172
rect 12967 -41198 13583 -40902
rect 13627 -40928 13923 -40902
rect 13627 -41172 13653 -40928
rect 13653 -41172 13897 -40928
rect 13897 -41172 13923 -40928
rect 13627 -41198 13923 -41172
rect 13967 -41198 14583 -40902
rect 14627 -40928 14923 -40902
rect 14627 -41172 14653 -40928
rect 14653 -41172 14897 -40928
rect 14897 -41172 14923 -40928
rect 14627 -41198 14923 -41172
rect 14967 -41198 15583 -40902
rect 15627 -40928 15923 -40902
rect 15627 -41172 15653 -40928
rect 15653 -41172 15897 -40928
rect 15897 -41172 15923 -40928
rect 15627 -41198 15923 -41172
rect 15967 -41198 16583 -40902
rect 16627 -40928 16923 -40902
rect 16627 -41172 16653 -40928
rect 16653 -41172 16897 -40928
rect 16897 -41172 16923 -40928
rect 16627 -41198 16923 -41172
rect 16967 -41198 17583 -40902
rect 17627 -40928 17923 -40902
rect 17627 -41172 17653 -40928
rect 17653 -41172 17897 -40928
rect 17897 -41172 17923 -40928
rect 17627 -41198 17923 -41172
rect 17967 -41198 18583 -40902
rect 18627 -40928 18923 -40902
rect 18627 -41172 18653 -40928
rect 18653 -41172 18897 -40928
rect 18897 -41172 18923 -40928
rect 18627 -41198 18923 -41172
rect 18967 -41198 19583 -40902
rect 19627 -40928 19923 -40902
rect 19627 -41172 19653 -40928
rect 19653 -41172 19897 -40928
rect 19897 -41172 19923 -40928
rect 19627 -41198 19923 -41172
rect 19967 -41198 20583 -40902
rect 20627 -40928 20923 -40902
rect 20627 -41172 20653 -40928
rect 20653 -41172 20897 -40928
rect 20897 -41172 20923 -40928
rect 20627 -41198 20923 -41172
rect 20967 -41198 21583 -40902
rect 21627 -40928 21923 -40902
rect 21627 -41172 21653 -40928
rect 21653 -41172 21897 -40928
rect 21897 -41172 21923 -40928
rect 21627 -41198 21923 -41172
rect 21967 -41198 22583 -40902
rect 22627 -40928 22923 -40902
rect 22627 -41172 22653 -40928
rect 22653 -41172 22897 -40928
rect 22897 -41172 22923 -40928
rect 22627 -41198 22923 -41172
rect 22967 -41198 23583 -40902
rect 23627 -40928 23923 -40902
rect 23627 -41172 23653 -40928
rect 23653 -41172 23897 -40928
rect 23897 -41172 23923 -40928
rect 23627 -41198 23923 -41172
rect 23967 -41198 24583 -40902
rect 24627 -40928 24923 -40902
rect 24627 -41172 24653 -40928
rect 24653 -41172 24897 -40928
rect 24897 -41172 24923 -40928
rect 24627 -41198 24923 -41172
rect 24967 -41198 25583 -40902
rect 25627 -40928 25923 -40902
rect 25627 -41172 25653 -40928
rect 25653 -41172 25897 -40928
rect 25897 -41172 25923 -40928
rect 25627 -41198 25923 -41172
rect 25967 -41198 26583 -40902
rect 26627 -40928 26923 -40902
rect 26627 -41172 26653 -40928
rect 26653 -41172 26897 -40928
rect 26897 -41172 26923 -40928
rect 26627 -41198 26923 -41172
rect 26967 -41198 27583 -40902
rect 27627 -40928 27923 -40902
rect 27627 -41172 27653 -40928
rect 27653 -41172 27897 -40928
rect 27897 -41172 27923 -40928
rect 27627 -41198 27923 -41172
rect 27967 -41198 28583 -40902
rect 28627 -40928 28923 -40902
rect 28627 -41172 28653 -40928
rect 28653 -41172 28897 -40928
rect 28897 -41172 28923 -40928
rect 28627 -41198 28923 -41172
rect 28967 -41198 29583 -40902
rect 29627 -40928 29923 -40902
rect 29627 -41172 29653 -40928
rect 29653 -41172 29897 -40928
rect 29897 -41172 29923 -40928
rect 29627 -41198 29923 -41172
rect 29967 -41198 30583 -40902
rect 30627 -40928 30923 -40902
rect 30627 -41172 30653 -40928
rect 30653 -41172 30897 -40928
rect 30897 -41172 30923 -40928
rect 30627 -41198 30923 -41172
rect 30967 -41198 31583 -40902
rect 31627 -40928 31923 -40902
rect 31627 -41172 31653 -40928
rect 31653 -41172 31897 -40928
rect 31897 -41172 31923 -40928
rect 31627 -41198 31923 -41172
rect 31967 -41198 32583 -40902
rect 32627 -40928 32923 -40902
rect 32627 -41172 32653 -40928
rect 32653 -41172 32897 -40928
rect 32897 -41172 32923 -40928
rect 32627 -41198 32923 -41172
rect 32967 -41198 33583 -40902
rect 33627 -40928 33923 -40902
rect 33627 -41172 33653 -40928
rect 33653 -41172 33897 -40928
rect 33897 -41172 33923 -40928
rect 33627 -41198 33923 -41172
rect 33967 -41198 34263 -40902
rect 8627 -41858 8923 -41242
rect 9627 -41858 9923 -41242
rect 10627 -41858 10923 -41242
rect 11627 -41858 11923 -41242
rect 12627 -41858 12923 -41242
rect 13627 -41858 13923 -41242
rect 14627 -41858 14923 -41242
rect 15627 -41858 15923 -41242
rect 16627 -41858 16923 -41242
rect 17627 -41858 17923 -41242
rect 18627 -41858 18923 -41242
rect 19627 -41858 19923 -41242
rect 20627 -41858 20923 -41242
rect 21627 -41858 21923 -41242
rect 22627 -41858 22923 -41242
rect 23627 -41858 23923 -41242
rect 24627 -41858 24923 -41242
rect 25627 -41858 25923 -41242
rect 26627 -41858 26923 -41242
rect 27627 -41858 27923 -41242
rect 28627 -41858 28923 -41242
rect 29627 -41858 29923 -41242
rect 30627 -41858 30923 -41242
rect 31627 -41858 31923 -41242
rect 32627 -41858 32923 -41242
rect 33627 -41858 33923 -41242
rect 8287 -42198 8583 -41902
rect 8627 -41928 8923 -41902
rect 8627 -42172 8653 -41928
rect 8653 -42172 8897 -41928
rect 8897 -42172 8923 -41928
rect 8627 -42198 8923 -42172
rect 8967 -42198 9583 -41902
rect 9627 -41928 9923 -41902
rect 9627 -42172 9653 -41928
rect 9653 -42172 9897 -41928
rect 9897 -42172 9923 -41928
rect 9627 -42198 9923 -42172
rect 9967 -42198 10583 -41902
rect 10627 -41928 10923 -41902
rect 10627 -42172 10653 -41928
rect 10653 -42172 10897 -41928
rect 10897 -42172 10923 -41928
rect 10627 -42198 10923 -42172
rect 10967 -42198 11583 -41902
rect 11627 -41928 11923 -41902
rect 11627 -42172 11653 -41928
rect 11653 -42172 11897 -41928
rect 11897 -42172 11923 -41928
rect 11627 -42198 11923 -42172
rect 11967 -42198 12583 -41902
rect 12627 -41928 12923 -41902
rect 12627 -42172 12653 -41928
rect 12653 -42172 12897 -41928
rect 12897 -42172 12923 -41928
rect 12627 -42198 12923 -42172
rect 12967 -42198 13583 -41902
rect 13627 -41928 13923 -41902
rect 13627 -42172 13653 -41928
rect 13653 -42172 13897 -41928
rect 13897 -42172 13923 -41928
rect 13627 -42198 13923 -42172
rect 13967 -42198 14583 -41902
rect 14627 -41928 14923 -41902
rect 14627 -42172 14653 -41928
rect 14653 -42172 14897 -41928
rect 14897 -42172 14923 -41928
rect 14627 -42198 14923 -42172
rect 14967 -42198 15583 -41902
rect 15627 -41928 15923 -41902
rect 15627 -42172 15653 -41928
rect 15653 -42172 15897 -41928
rect 15897 -42172 15923 -41928
rect 15627 -42198 15923 -42172
rect 15967 -42198 16583 -41902
rect 16627 -41928 16923 -41902
rect 16627 -42172 16653 -41928
rect 16653 -42172 16897 -41928
rect 16897 -42172 16923 -41928
rect 16627 -42198 16923 -42172
rect 16967 -42198 17583 -41902
rect 17627 -41928 17923 -41902
rect 17627 -42172 17653 -41928
rect 17653 -42172 17897 -41928
rect 17897 -42172 17923 -41928
rect 17627 -42198 17923 -42172
rect 17967 -42198 18583 -41902
rect 18627 -41928 18923 -41902
rect 18627 -42172 18653 -41928
rect 18653 -42172 18897 -41928
rect 18897 -42172 18923 -41928
rect 18627 -42198 18923 -42172
rect 18967 -42198 19583 -41902
rect 19627 -41928 19923 -41902
rect 19627 -42172 19653 -41928
rect 19653 -42172 19897 -41928
rect 19897 -42172 19923 -41928
rect 19627 -42198 19923 -42172
rect 19967 -42198 20583 -41902
rect 20627 -41928 20923 -41902
rect 20627 -42172 20653 -41928
rect 20653 -42172 20897 -41928
rect 20897 -42172 20923 -41928
rect 20627 -42198 20923 -42172
rect 20967 -42198 21583 -41902
rect 21627 -41928 21923 -41902
rect 21627 -42172 21653 -41928
rect 21653 -42172 21897 -41928
rect 21897 -42172 21923 -41928
rect 21627 -42198 21923 -42172
rect 21967 -42198 22583 -41902
rect 22627 -41928 22923 -41902
rect 22627 -42172 22653 -41928
rect 22653 -42172 22897 -41928
rect 22897 -42172 22923 -41928
rect 22627 -42198 22923 -42172
rect 22967 -42198 23583 -41902
rect 23627 -41928 23923 -41902
rect 23627 -42172 23653 -41928
rect 23653 -42172 23897 -41928
rect 23897 -42172 23923 -41928
rect 23627 -42198 23923 -42172
rect 23967 -42198 24583 -41902
rect 24627 -41928 24923 -41902
rect 24627 -42172 24653 -41928
rect 24653 -42172 24897 -41928
rect 24897 -42172 24923 -41928
rect 24627 -42198 24923 -42172
rect 24967 -42198 25583 -41902
rect 25627 -41928 25923 -41902
rect 25627 -42172 25653 -41928
rect 25653 -42172 25897 -41928
rect 25897 -42172 25923 -41928
rect 25627 -42198 25923 -42172
rect 25967 -42198 26583 -41902
rect 26627 -41928 26923 -41902
rect 26627 -42172 26653 -41928
rect 26653 -42172 26897 -41928
rect 26897 -42172 26923 -41928
rect 26627 -42198 26923 -42172
rect 26967 -42198 27583 -41902
rect 27627 -41928 27923 -41902
rect 27627 -42172 27653 -41928
rect 27653 -42172 27897 -41928
rect 27897 -42172 27923 -41928
rect 27627 -42198 27923 -42172
rect 27967 -42198 28583 -41902
rect 28627 -41928 28923 -41902
rect 28627 -42172 28653 -41928
rect 28653 -42172 28897 -41928
rect 28897 -42172 28923 -41928
rect 28627 -42198 28923 -42172
rect 28967 -42198 29583 -41902
rect 29627 -41928 29923 -41902
rect 29627 -42172 29653 -41928
rect 29653 -42172 29897 -41928
rect 29897 -42172 29923 -41928
rect 29627 -42198 29923 -42172
rect 29967 -42198 30583 -41902
rect 30627 -41928 30923 -41902
rect 30627 -42172 30653 -41928
rect 30653 -42172 30897 -41928
rect 30897 -42172 30923 -41928
rect 30627 -42198 30923 -42172
rect 30967 -42198 31583 -41902
rect 31627 -41928 31923 -41902
rect 31627 -42172 31653 -41928
rect 31653 -42172 31897 -41928
rect 31897 -42172 31923 -41928
rect 31627 -42198 31923 -42172
rect 31967 -42198 32583 -41902
rect 32627 -41928 32923 -41902
rect 32627 -42172 32653 -41928
rect 32653 -42172 32897 -41928
rect 32897 -42172 32923 -41928
rect 32627 -42198 32923 -42172
rect 32967 -42198 33583 -41902
rect 33627 -41928 33923 -41902
rect 33627 -42172 33653 -41928
rect 33653 -42172 33897 -41928
rect 33897 -42172 33923 -41928
rect 33627 -42198 33923 -42172
rect 33967 -42198 34263 -41902
rect 8627 -42858 8923 -42242
rect 9627 -42858 9923 -42242
rect 10627 -42858 10923 -42242
rect 11627 -42858 11923 -42242
rect 12627 -42858 12923 -42242
rect 13627 -42858 13923 -42242
rect 14627 -42858 14923 -42242
rect 15627 -42858 15923 -42242
rect 16627 -42858 16923 -42242
rect 17627 -42858 17923 -42242
rect 18627 -42858 18923 -42242
rect 19627 -42858 19923 -42242
rect 20627 -42858 20923 -42242
rect 21627 -42858 21923 -42242
rect 22627 -42858 22923 -42242
rect 23627 -42858 23923 -42242
rect 24627 -42858 24923 -42242
rect 25627 -42858 25923 -42242
rect 26627 -42858 26923 -42242
rect 27627 -42858 27923 -42242
rect 28627 -42858 28923 -42242
rect 29627 -42858 29923 -42242
rect 30627 -42858 30923 -42242
rect 31627 -42858 31923 -42242
rect 32627 -42858 32923 -42242
rect 33627 -42858 33923 -42242
rect 8287 -43198 8583 -42902
rect 8627 -42928 8923 -42902
rect 8627 -43172 8653 -42928
rect 8653 -43172 8897 -42928
rect 8897 -43172 8923 -42928
rect 8627 -43198 8923 -43172
rect 8967 -43198 9583 -42902
rect 9627 -42928 9923 -42902
rect 9627 -43172 9653 -42928
rect 9653 -43172 9897 -42928
rect 9897 -43172 9923 -42928
rect 9627 -43198 9923 -43172
rect 9967 -43198 10583 -42902
rect 10627 -42928 10923 -42902
rect 10627 -43172 10653 -42928
rect 10653 -43172 10897 -42928
rect 10897 -43172 10923 -42928
rect 10627 -43198 10923 -43172
rect 10967 -43198 11583 -42902
rect 11627 -42928 11923 -42902
rect 11627 -43172 11653 -42928
rect 11653 -43172 11897 -42928
rect 11897 -43172 11923 -42928
rect 11627 -43198 11923 -43172
rect 11967 -43198 12583 -42902
rect 12627 -42928 12923 -42902
rect 12627 -43172 12653 -42928
rect 12653 -43172 12897 -42928
rect 12897 -43172 12923 -42928
rect 12627 -43198 12923 -43172
rect 12967 -43198 13583 -42902
rect 13627 -42928 13923 -42902
rect 13627 -43172 13653 -42928
rect 13653 -43172 13897 -42928
rect 13897 -43172 13923 -42928
rect 13627 -43198 13923 -43172
rect 13967 -43198 14583 -42902
rect 14627 -42928 14923 -42902
rect 14627 -43172 14653 -42928
rect 14653 -43172 14897 -42928
rect 14897 -43172 14923 -42928
rect 14627 -43198 14923 -43172
rect 14967 -43198 15583 -42902
rect 15627 -42928 15923 -42902
rect 15627 -43172 15653 -42928
rect 15653 -43172 15897 -42928
rect 15897 -43172 15923 -42928
rect 15627 -43198 15923 -43172
rect 15967 -43198 16583 -42902
rect 16627 -42928 16923 -42902
rect 16627 -43172 16653 -42928
rect 16653 -43172 16897 -42928
rect 16897 -43172 16923 -42928
rect 16627 -43198 16923 -43172
rect 16967 -43198 17583 -42902
rect 17627 -42928 17923 -42902
rect 17627 -43172 17653 -42928
rect 17653 -43172 17897 -42928
rect 17897 -43172 17923 -42928
rect 17627 -43198 17923 -43172
rect 17967 -43198 18583 -42902
rect 18627 -42928 18923 -42902
rect 18627 -43172 18653 -42928
rect 18653 -43172 18897 -42928
rect 18897 -43172 18923 -42928
rect 18627 -43198 18923 -43172
rect 18967 -43198 19583 -42902
rect 19627 -42928 19923 -42902
rect 19627 -43172 19653 -42928
rect 19653 -43172 19897 -42928
rect 19897 -43172 19923 -42928
rect 19627 -43198 19923 -43172
rect 19967 -43198 20583 -42902
rect 20627 -42928 20923 -42902
rect 20627 -43172 20653 -42928
rect 20653 -43172 20897 -42928
rect 20897 -43172 20923 -42928
rect 20627 -43198 20923 -43172
rect 20967 -43198 21583 -42902
rect 21627 -42928 21923 -42902
rect 21627 -43172 21653 -42928
rect 21653 -43172 21897 -42928
rect 21897 -43172 21923 -42928
rect 21627 -43198 21923 -43172
rect 21967 -43198 22583 -42902
rect 22627 -42928 22923 -42902
rect 22627 -43172 22653 -42928
rect 22653 -43172 22897 -42928
rect 22897 -43172 22923 -42928
rect 22627 -43198 22923 -43172
rect 22967 -43198 23583 -42902
rect 23627 -42928 23923 -42902
rect 23627 -43172 23653 -42928
rect 23653 -43172 23897 -42928
rect 23897 -43172 23923 -42928
rect 23627 -43198 23923 -43172
rect 23967 -43198 24583 -42902
rect 24627 -42928 24923 -42902
rect 24627 -43172 24653 -42928
rect 24653 -43172 24897 -42928
rect 24897 -43172 24923 -42928
rect 24627 -43198 24923 -43172
rect 24967 -43198 25583 -42902
rect 25627 -42928 25923 -42902
rect 25627 -43172 25653 -42928
rect 25653 -43172 25897 -42928
rect 25897 -43172 25923 -42928
rect 25627 -43198 25923 -43172
rect 25967 -43198 26583 -42902
rect 26627 -42928 26923 -42902
rect 26627 -43172 26653 -42928
rect 26653 -43172 26897 -42928
rect 26897 -43172 26923 -42928
rect 26627 -43198 26923 -43172
rect 26967 -43198 27583 -42902
rect 27627 -42928 27923 -42902
rect 27627 -43172 27653 -42928
rect 27653 -43172 27897 -42928
rect 27897 -43172 27923 -42928
rect 27627 -43198 27923 -43172
rect 27967 -43198 28583 -42902
rect 28627 -42928 28923 -42902
rect 28627 -43172 28653 -42928
rect 28653 -43172 28897 -42928
rect 28897 -43172 28923 -42928
rect 28627 -43198 28923 -43172
rect 28967 -43198 29583 -42902
rect 29627 -42928 29923 -42902
rect 29627 -43172 29653 -42928
rect 29653 -43172 29897 -42928
rect 29897 -43172 29923 -42928
rect 29627 -43198 29923 -43172
rect 29967 -43198 30583 -42902
rect 30627 -42928 30923 -42902
rect 30627 -43172 30653 -42928
rect 30653 -43172 30897 -42928
rect 30897 -43172 30923 -42928
rect 30627 -43198 30923 -43172
rect 30967 -43198 31583 -42902
rect 31627 -42928 31923 -42902
rect 31627 -43172 31653 -42928
rect 31653 -43172 31897 -42928
rect 31897 -43172 31923 -42928
rect 31627 -43198 31923 -43172
rect 31967 -43198 32583 -42902
rect 32627 -42928 32923 -42902
rect 32627 -43172 32653 -42928
rect 32653 -43172 32897 -42928
rect 32897 -43172 32923 -42928
rect 32627 -43198 32923 -43172
rect 32967 -43198 33583 -42902
rect 33627 -42928 33923 -42902
rect 33627 -43172 33653 -42928
rect 33653 -43172 33897 -42928
rect 33897 -43172 33923 -42928
rect 33627 -43198 33923 -43172
rect 33967 -43198 34263 -42902
rect 8627 -43858 8923 -43242
rect 9627 -43858 9923 -43242
rect 10627 -43858 10923 -43242
rect 11627 -43858 11923 -43242
rect 12627 -43858 12923 -43242
rect 13627 -43858 13923 -43242
rect 14627 -43858 14923 -43242
rect 15627 -43858 15923 -43242
rect 16627 -43858 16923 -43242
rect 17627 -43858 17923 -43242
rect 18627 -43858 18923 -43242
rect 19627 -43858 19923 -43242
rect 20627 -43858 20923 -43242
rect 21627 -43858 21923 -43242
rect 22627 -43858 22923 -43242
rect 23627 -43858 23923 -43242
rect 24627 -43858 24923 -43242
rect 25627 -43858 25923 -43242
rect 26627 -43858 26923 -43242
rect 27627 -43858 27923 -43242
rect 28627 -43858 28923 -43242
rect 29627 -43858 29923 -43242
rect 30627 -43858 30923 -43242
rect 31627 -43858 31923 -43242
rect 32627 -43858 32923 -43242
rect 33627 -43858 33923 -43242
rect 8287 -44198 8583 -43902
rect 8627 -43928 8923 -43902
rect 8627 -44172 8653 -43928
rect 8653 -44172 8897 -43928
rect 8897 -44172 8923 -43928
rect 8627 -44198 8923 -44172
rect 8967 -44198 9583 -43902
rect 9627 -43928 9923 -43902
rect 9627 -44172 9653 -43928
rect 9653 -44172 9897 -43928
rect 9897 -44172 9923 -43928
rect 9627 -44198 9923 -44172
rect 9967 -44198 10583 -43902
rect 10627 -43928 10923 -43902
rect 10627 -44172 10653 -43928
rect 10653 -44172 10897 -43928
rect 10897 -44172 10923 -43928
rect 10627 -44198 10923 -44172
rect 10967 -44198 11583 -43902
rect 11627 -43928 11923 -43902
rect 11627 -44172 11653 -43928
rect 11653 -44172 11897 -43928
rect 11897 -44172 11923 -43928
rect 11627 -44198 11923 -44172
rect 11967 -44198 12583 -43902
rect 12627 -43928 12923 -43902
rect 12627 -44172 12653 -43928
rect 12653 -44172 12897 -43928
rect 12897 -44172 12923 -43928
rect 12627 -44198 12923 -44172
rect 12967 -44198 13583 -43902
rect 13627 -43928 13923 -43902
rect 13627 -44172 13653 -43928
rect 13653 -44172 13897 -43928
rect 13897 -44172 13923 -43928
rect 13627 -44198 13923 -44172
rect 13967 -44198 14583 -43902
rect 14627 -43928 14923 -43902
rect 14627 -44172 14653 -43928
rect 14653 -44172 14897 -43928
rect 14897 -44172 14923 -43928
rect 14627 -44198 14923 -44172
rect 14967 -44198 15583 -43902
rect 15627 -43928 15923 -43902
rect 15627 -44172 15653 -43928
rect 15653 -44172 15897 -43928
rect 15897 -44172 15923 -43928
rect 15627 -44198 15923 -44172
rect 15967 -44198 16583 -43902
rect 16627 -43928 16923 -43902
rect 16627 -44172 16653 -43928
rect 16653 -44172 16897 -43928
rect 16897 -44172 16923 -43928
rect 16627 -44198 16923 -44172
rect 16967 -44198 17583 -43902
rect 17627 -43928 17923 -43902
rect 17627 -44172 17653 -43928
rect 17653 -44172 17897 -43928
rect 17897 -44172 17923 -43928
rect 17627 -44198 17923 -44172
rect 17967 -44198 18583 -43902
rect 18627 -43928 18923 -43902
rect 18627 -44172 18653 -43928
rect 18653 -44172 18897 -43928
rect 18897 -44172 18923 -43928
rect 18627 -44198 18923 -44172
rect 18967 -44198 19583 -43902
rect 19627 -43928 19923 -43902
rect 19627 -44172 19653 -43928
rect 19653 -44172 19897 -43928
rect 19897 -44172 19923 -43928
rect 19627 -44198 19923 -44172
rect 19967 -44198 20583 -43902
rect 20627 -43928 20923 -43902
rect 20627 -44172 20653 -43928
rect 20653 -44172 20897 -43928
rect 20897 -44172 20923 -43928
rect 20627 -44198 20923 -44172
rect 20967 -44198 21583 -43902
rect 21627 -43928 21923 -43902
rect 21627 -44172 21653 -43928
rect 21653 -44172 21897 -43928
rect 21897 -44172 21923 -43928
rect 21627 -44198 21923 -44172
rect 21967 -44198 22583 -43902
rect 22627 -43928 22923 -43902
rect 22627 -44172 22653 -43928
rect 22653 -44172 22897 -43928
rect 22897 -44172 22923 -43928
rect 22627 -44198 22923 -44172
rect 22967 -44198 23583 -43902
rect 23627 -43928 23923 -43902
rect 23627 -44172 23653 -43928
rect 23653 -44172 23897 -43928
rect 23897 -44172 23923 -43928
rect 23627 -44198 23923 -44172
rect 23967 -44198 24583 -43902
rect 24627 -43928 24923 -43902
rect 24627 -44172 24653 -43928
rect 24653 -44172 24897 -43928
rect 24897 -44172 24923 -43928
rect 24627 -44198 24923 -44172
rect 24967 -44198 25583 -43902
rect 25627 -43928 25923 -43902
rect 25627 -44172 25653 -43928
rect 25653 -44172 25897 -43928
rect 25897 -44172 25923 -43928
rect 25627 -44198 25923 -44172
rect 25967 -44198 26583 -43902
rect 26627 -43928 26923 -43902
rect 26627 -44172 26653 -43928
rect 26653 -44172 26897 -43928
rect 26897 -44172 26923 -43928
rect 26627 -44198 26923 -44172
rect 26967 -44198 27583 -43902
rect 27627 -43928 27923 -43902
rect 27627 -44172 27653 -43928
rect 27653 -44172 27897 -43928
rect 27897 -44172 27923 -43928
rect 27627 -44198 27923 -44172
rect 27967 -44198 28583 -43902
rect 28627 -43928 28923 -43902
rect 28627 -44172 28653 -43928
rect 28653 -44172 28897 -43928
rect 28897 -44172 28923 -43928
rect 28627 -44198 28923 -44172
rect 28967 -44198 29583 -43902
rect 29627 -43928 29923 -43902
rect 29627 -44172 29653 -43928
rect 29653 -44172 29897 -43928
rect 29897 -44172 29923 -43928
rect 29627 -44198 29923 -44172
rect 29967 -44198 30583 -43902
rect 30627 -43928 30923 -43902
rect 30627 -44172 30653 -43928
rect 30653 -44172 30897 -43928
rect 30897 -44172 30923 -43928
rect 30627 -44198 30923 -44172
rect 30967 -44198 31583 -43902
rect 31627 -43928 31923 -43902
rect 31627 -44172 31653 -43928
rect 31653 -44172 31897 -43928
rect 31897 -44172 31923 -43928
rect 31627 -44198 31923 -44172
rect 31967 -44198 32583 -43902
rect 32627 -43928 32923 -43902
rect 32627 -44172 32653 -43928
rect 32653 -44172 32897 -43928
rect 32897 -44172 32923 -43928
rect 32627 -44198 32923 -44172
rect 32967 -44198 33583 -43902
rect 33627 -43928 33923 -43902
rect 33627 -44172 33653 -43928
rect 33653 -44172 33897 -43928
rect 33897 -44172 33923 -43928
rect 33627 -44198 33923 -44172
rect 33967 -44198 34263 -43902
rect -4228 -44498 5668 -44496
rect 8627 -44858 8923 -44242
rect 9627 -44858 9923 -44242
rect 10627 -44858 10923 -44242
rect 11627 -44858 11923 -44242
rect 12627 -44858 12923 -44242
rect 13627 -44858 13923 -44242
rect 14627 -44858 14923 -44242
rect 15627 -44858 15923 -44242
rect 16627 -44858 16923 -44242
rect 17627 -44858 17923 -44242
rect 18627 -44858 18923 -44242
rect 19627 -44858 19923 -44242
rect 20627 -44858 20923 -44242
rect 21627 -44858 21923 -44242
rect 22627 -44858 22923 -44242
rect 23627 -44858 23923 -44242
rect 24627 -44858 24923 -44242
rect 25627 -44858 25923 -44242
rect 26627 -44858 26923 -44242
rect 27627 -44858 27923 -44242
rect 28627 -44858 28923 -44242
rect 29627 -44858 29923 -44242
rect 30627 -44858 30923 -44242
rect 31627 -44858 31923 -44242
rect 32627 -44858 32923 -44242
rect 33627 -44858 33923 -44242
rect -74813 -45198 -74517 -44902
rect -74473 -44928 -74177 -44902
rect -74473 -45172 -74447 -44928
rect -74447 -45172 -74203 -44928
rect -74203 -45172 -74177 -44928
rect -74473 -45198 -74177 -45172
rect -74133 -45198 -73517 -44902
rect -73473 -44928 -73177 -44902
rect -73473 -45172 -73447 -44928
rect -73447 -45172 -73203 -44928
rect -73203 -45172 -73177 -44928
rect -73473 -45198 -73177 -45172
rect -73133 -45198 -72517 -44902
rect -72473 -44928 -72177 -44902
rect -72473 -45172 -72447 -44928
rect -72447 -45172 -72203 -44928
rect -72203 -45172 -72177 -44928
rect -72473 -45198 -72177 -45172
rect -72133 -45198 -71517 -44902
rect -71473 -44928 -71177 -44902
rect -71473 -45172 -71447 -44928
rect -71447 -45172 -71203 -44928
rect -71203 -45172 -71177 -44928
rect -71473 -45198 -71177 -45172
rect -71133 -45198 -70517 -44902
rect -70473 -44928 -70177 -44902
rect -70473 -45172 -70447 -44928
rect -70447 -45172 -70203 -44928
rect -70203 -45172 -70177 -44928
rect -70473 -45198 -70177 -45172
rect -70133 -45198 -69517 -44902
rect -69473 -44928 -69177 -44902
rect -69473 -45172 -69447 -44928
rect -69447 -45172 -69203 -44928
rect -69203 -45172 -69177 -44928
rect -69473 -45198 -69177 -45172
rect -69133 -45198 -68517 -44902
rect -68473 -44928 -68177 -44902
rect -68473 -45172 -68447 -44928
rect -68447 -45172 -68203 -44928
rect -68203 -45172 -68177 -44928
rect -68473 -45198 -68177 -45172
rect -68133 -45198 -67517 -44902
rect -67473 -44928 -67177 -44902
rect -67473 -45172 -67447 -44928
rect -67447 -45172 -67203 -44928
rect -67203 -45172 -67177 -44928
rect -67473 -45198 -67177 -45172
rect -67133 -45198 -66517 -44902
rect -66473 -44928 -66177 -44902
rect -66473 -45172 -66447 -44928
rect -66447 -45172 -66203 -44928
rect -66203 -45172 -66177 -44928
rect -66473 -45198 -66177 -45172
rect -66133 -45198 -65517 -44902
rect -65473 -44928 -65177 -44902
rect -65473 -45172 -65447 -44928
rect -65447 -45172 -65203 -44928
rect -65203 -45172 -65177 -44928
rect -65473 -45198 -65177 -45172
rect -65133 -45198 -64517 -44902
rect -64473 -44928 -64177 -44902
rect -64473 -45172 -64447 -44928
rect -64447 -45172 -64203 -44928
rect -64203 -45172 -64177 -44928
rect -64473 -45198 -64177 -45172
rect -64133 -45198 -63517 -44902
rect -63473 -44928 -63177 -44902
rect -63473 -45172 -63447 -44928
rect -63447 -45172 -63203 -44928
rect -63203 -45172 -63177 -44928
rect -63473 -45198 -63177 -45172
rect -63133 -45198 -62517 -44902
rect -62473 -44928 -62177 -44902
rect -62473 -45172 -62447 -44928
rect -62447 -45172 -62203 -44928
rect -62203 -45172 -62177 -44928
rect -62473 -45198 -62177 -45172
rect -62133 -45198 -61517 -44902
rect -61473 -44928 -61177 -44902
rect -61473 -45172 -61447 -44928
rect -61447 -45172 -61203 -44928
rect -61203 -45172 -61177 -44928
rect -61473 -45198 -61177 -45172
rect -61133 -45198 -60517 -44902
rect -60473 -44928 -60177 -44902
rect -60473 -45172 -60447 -44928
rect -60447 -45172 -60203 -44928
rect -60203 -45172 -60177 -44928
rect -60473 -45198 -60177 -45172
rect -60133 -45198 -59517 -44902
rect -59473 -44928 -59177 -44902
rect -59473 -45172 -59447 -44928
rect -59447 -45172 -59203 -44928
rect -59203 -45172 -59177 -44928
rect -59473 -45198 -59177 -45172
rect -59133 -45198 -58517 -44902
rect -58473 -44928 -58177 -44902
rect -58473 -45172 -58447 -44928
rect -58447 -45172 -58203 -44928
rect -58203 -45172 -58177 -44928
rect -58473 -45198 -58177 -45172
rect -58133 -45198 -57517 -44902
rect -57473 -44928 -57177 -44902
rect -57473 -45172 -57447 -44928
rect -57447 -45172 -57203 -44928
rect -57203 -45172 -57177 -44928
rect -57473 -45198 -57177 -45172
rect -57133 -45198 -56517 -44902
rect -56473 -44928 -56177 -44902
rect -56473 -45172 -56447 -44928
rect -56447 -45172 -56203 -44928
rect -56203 -45172 -56177 -44928
rect -56473 -45198 -56177 -45172
rect -56133 -45198 -55517 -44902
rect -55473 -44928 -55177 -44902
rect -55473 -45172 -55447 -44928
rect -55447 -45172 -55203 -44928
rect -55203 -45172 -55177 -44928
rect -55473 -45198 -55177 -45172
rect -55133 -45198 -54517 -44902
rect -54473 -44928 -54177 -44902
rect -54473 -45172 -54447 -44928
rect -54447 -45172 -54203 -44928
rect -54203 -45172 -54177 -44928
rect -54473 -45198 -54177 -45172
rect -54133 -45198 -53517 -44902
rect -53473 -44928 -53177 -44902
rect -53473 -45172 -53447 -44928
rect -53447 -45172 -53203 -44928
rect -53203 -45172 -53177 -44928
rect -53473 -45198 -53177 -45172
rect -53133 -45198 -52517 -44902
rect -52473 -44928 -52177 -44902
rect -52473 -45172 -52447 -44928
rect -52447 -45172 -52203 -44928
rect -52203 -45172 -52177 -44928
rect -52473 -45198 -52177 -45172
rect -52133 -45198 -51517 -44902
rect -51473 -44928 -51177 -44902
rect -51473 -45172 -51447 -44928
rect -51447 -45172 -51203 -44928
rect -51203 -45172 -51177 -44928
rect -51473 -45198 -51177 -45172
rect -51133 -45198 -50517 -44902
rect -50473 -44928 -50177 -44902
rect -50473 -45172 -50447 -44928
rect -50447 -45172 -50203 -44928
rect -50203 -45172 -50177 -44928
rect -50473 -45198 -50177 -45172
rect -50133 -45198 -49517 -44902
rect -49473 -44928 -49177 -44902
rect -49473 -45172 -49447 -44928
rect -49447 -45172 -49203 -44928
rect -49203 -45172 -49177 -44928
rect -49473 -45198 -49177 -45172
rect -49133 -45198 -48837 -44902
rect 8287 -45198 8583 -44902
rect 8627 -44928 8923 -44902
rect 8627 -45172 8653 -44928
rect 8653 -45172 8897 -44928
rect 8897 -45172 8923 -44928
rect 8627 -45198 8923 -45172
rect 8967 -45198 9583 -44902
rect 9627 -44928 9923 -44902
rect 9627 -45172 9653 -44928
rect 9653 -45172 9897 -44928
rect 9897 -45172 9923 -44928
rect 9627 -45198 9923 -45172
rect 9967 -45198 10583 -44902
rect 10627 -44928 10923 -44902
rect 10627 -45172 10653 -44928
rect 10653 -45172 10897 -44928
rect 10897 -45172 10923 -44928
rect 10627 -45198 10923 -45172
rect 10967 -45198 11583 -44902
rect 11627 -44928 11923 -44902
rect 11627 -45172 11653 -44928
rect 11653 -45172 11897 -44928
rect 11897 -45172 11923 -44928
rect 11627 -45198 11923 -45172
rect 11967 -45198 12583 -44902
rect 12627 -44928 12923 -44902
rect 12627 -45172 12653 -44928
rect 12653 -45172 12897 -44928
rect 12897 -45172 12923 -44928
rect 12627 -45198 12923 -45172
rect 12967 -45198 13583 -44902
rect 13627 -44928 13923 -44902
rect 13627 -45172 13653 -44928
rect 13653 -45172 13897 -44928
rect 13897 -45172 13923 -44928
rect 13627 -45198 13923 -45172
rect 13967 -45198 14583 -44902
rect 14627 -44928 14923 -44902
rect 14627 -45172 14653 -44928
rect 14653 -45172 14897 -44928
rect 14897 -45172 14923 -44928
rect 14627 -45198 14923 -45172
rect 14967 -45198 15583 -44902
rect 15627 -44928 15923 -44902
rect 15627 -45172 15653 -44928
rect 15653 -45172 15897 -44928
rect 15897 -45172 15923 -44928
rect 15627 -45198 15923 -45172
rect 15967 -45198 16583 -44902
rect 16627 -44928 16923 -44902
rect 16627 -45172 16653 -44928
rect 16653 -45172 16897 -44928
rect 16897 -45172 16923 -44928
rect 16627 -45198 16923 -45172
rect 16967 -45198 17583 -44902
rect 17627 -44928 17923 -44902
rect 17627 -45172 17653 -44928
rect 17653 -45172 17897 -44928
rect 17897 -45172 17923 -44928
rect 17627 -45198 17923 -45172
rect 17967 -45198 18583 -44902
rect 18627 -44928 18923 -44902
rect 18627 -45172 18653 -44928
rect 18653 -45172 18897 -44928
rect 18897 -45172 18923 -44928
rect 18627 -45198 18923 -45172
rect 18967 -45198 19583 -44902
rect 19627 -44928 19923 -44902
rect 19627 -45172 19653 -44928
rect 19653 -45172 19897 -44928
rect 19897 -45172 19923 -44928
rect 19627 -45198 19923 -45172
rect 19967 -45198 20583 -44902
rect 20627 -44928 20923 -44902
rect 20627 -45172 20653 -44928
rect 20653 -45172 20897 -44928
rect 20897 -45172 20923 -44928
rect 20627 -45198 20923 -45172
rect 20967 -45198 21583 -44902
rect 21627 -44928 21923 -44902
rect 21627 -45172 21653 -44928
rect 21653 -45172 21897 -44928
rect 21897 -45172 21923 -44928
rect 21627 -45198 21923 -45172
rect 21967 -45198 22583 -44902
rect 22627 -44928 22923 -44902
rect 22627 -45172 22653 -44928
rect 22653 -45172 22897 -44928
rect 22897 -45172 22923 -44928
rect 22627 -45198 22923 -45172
rect 22967 -45198 23583 -44902
rect 23627 -44928 23923 -44902
rect 23627 -45172 23653 -44928
rect 23653 -45172 23897 -44928
rect 23897 -45172 23923 -44928
rect 23627 -45198 23923 -45172
rect 23967 -45198 24583 -44902
rect 24627 -44928 24923 -44902
rect 24627 -45172 24653 -44928
rect 24653 -45172 24897 -44928
rect 24897 -45172 24923 -44928
rect 24627 -45198 24923 -45172
rect 24967 -45198 25583 -44902
rect 25627 -44928 25923 -44902
rect 25627 -45172 25653 -44928
rect 25653 -45172 25897 -44928
rect 25897 -45172 25923 -44928
rect 25627 -45198 25923 -45172
rect 25967 -45198 26583 -44902
rect 26627 -44928 26923 -44902
rect 26627 -45172 26653 -44928
rect 26653 -45172 26897 -44928
rect 26897 -45172 26923 -44928
rect 26627 -45198 26923 -45172
rect 26967 -45198 27583 -44902
rect 27627 -44928 27923 -44902
rect 27627 -45172 27653 -44928
rect 27653 -45172 27897 -44928
rect 27897 -45172 27923 -44928
rect 27627 -45198 27923 -45172
rect 27967 -45198 28583 -44902
rect 28627 -44928 28923 -44902
rect 28627 -45172 28653 -44928
rect 28653 -45172 28897 -44928
rect 28897 -45172 28923 -44928
rect 28627 -45198 28923 -45172
rect 28967 -45198 29583 -44902
rect 29627 -44928 29923 -44902
rect 29627 -45172 29653 -44928
rect 29653 -45172 29897 -44928
rect 29897 -45172 29923 -44928
rect 29627 -45198 29923 -45172
rect 29967 -45198 30583 -44902
rect 30627 -44928 30923 -44902
rect 30627 -45172 30653 -44928
rect 30653 -45172 30897 -44928
rect 30897 -45172 30923 -44928
rect 30627 -45198 30923 -45172
rect 30967 -45198 31583 -44902
rect 31627 -44928 31923 -44902
rect 31627 -45172 31653 -44928
rect 31653 -45172 31897 -44928
rect 31897 -45172 31923 -44928
rect 31627 -45198 31923 -45172
rect 31967 -45198 32583 -44902
rect 32627 -44928 32923 -44902
rect 32627 -45172 32653 -44928
rect 32653 -45172 32897 -44928
rect 32897 -45172 32923 -44928
rect 32627 -45198 32923 -45172
rect 32967 -45198 33583 -44902
rect 33627 -44928 33923 -44902
rect 33627 -45172 33653 -44928
rect 33653 -45172 33897 -44928
rect 33897 -45172 33923 -44928
rect 33627 -45198 33923 -45172
rect 33967 -45198 34263 -44902
rect -74473 -45858 -74177 -45242
rect -73473 -45858 -73177 -45242
rect -72473 -45858 -72177 -45242
rect -71473 -45858 -71177 -45242
rect -70473 -45858 -70177 -45242
rect -69473 -45858 -69177 -45242
rect -68473 -45858 -68177 -45242
rect -67473 -45858 -67177 -45242
rect -66473 -45858 -66177 -45242
rect -65473 -45858 -65177 -45242
rect -64473 -45858 -64177 -45242
rect -63473 -45858 -63177 -45242
rect -62473 -45858 -62177 -45242
rect -61473 -45858 -61177 -45242
rect -60473 -45858 -60177 -45242
rect -59473 -45858 -59177 -45242
rect -58473 -45858 -58177 -45242
rect -57473 -45858 -57177 -45242
rect -56473 -45858 -56177 -45242
rect -55473 -45858 -55177 -45242
rect -54473 -45858 -54177 -45242
rect -53473 -45858 -53177 -45242
rect -52473 -45858 -52177 -45242
rect -51473 -45858 -51177 -45242
rect -50473 -45858 -50177 -45242
rect -49473 -45858 -49177 -45242
rect 8627 -45858 8923 -45242
rect 9627 -45858 9923 -45242
rect 10627 -45858 10923 -45242
rect 11627 -45858 11923 -45242
rect 12627 -45858 12923 -45242
rect 13627 -45858 13923 -45242
rect 14627 -45858 14923 -45242
rect 15627 -45858 15923 -45242
rect 16627 -45858 16923 -45242
rect 17627 -45858 17923 -45242
rect 18627 -45858 18923 -45242
rect 19627 -45858 19923 -45242
rect 20627 -45858 20923 -45242
rect 21627 -45858 21923 -45242
rect 22627 -45858 22923 -45242
rect 23627 -45858 23923 -45242
rect 24627 -45858 24923 -45242
rect 25627 -45858 25923 -45242
rect 26627 -45858 26923 -45242
rect 27627 -45858 27923 -45242
rect 28627 -45858 28923 -45242
rect 29627 -45858 29923 -45242
rect 30627 -45858 30923 -45242
rect 31627 -45858 31923 -45242
rect 32627 -45858 32923 -45242
rect 33627 -45858 33923 -45242
rect -74813 -46198 -74517 -45902
rect -74473 -45928 -74177 -45902
rect -74473 -46172 -74447 -45928
rect -74447 -46172 -74203 -45928
rect -74203 -46172 -74177 -45928
rect -74473 -46198 -74177 -46172
rect -74133 -46198 -73517 -45902
rect -73473 -45928 -73177 -45902
rect -73473 -46172 -73447 -45928
rect -73447 -46172 -73203 -45928
rect -73203 -46172 -73177 -45928
rect -73473 -46198 -73177 -46172
rect -73133 -46198 -72517 -45902
rect -72473 -45928 -72177 -45902
rect -72473 -46172 -72447 -45928
rect -72447 -46172 -72203 -45928
rect -72203 -46172 -72177 -45928
rect -72473 -46198 -72177 -46172
rect -72133 -46198 -71517 -45902
rect -71473 -45928 -71177 -45902
rect -71473 -46172 -71447 -45928
rect -71447 -46172 -71203 -45928
rect -71203 -46172 -71177 -45928
rect -71473 -46198 -71177 -46172
rect -71133 -46198 -70517 -45902
rect -70473 -45928 -70177 -45902
rect -70473 -46172 -70447 -45928
rect -70447 -46172 -70203 -45928
rect -70203 -46172 -70177 -45928
rect -70473 -46198 -70177 -46172
rect -70133 -46198 -69517 -45902
rect -69473 -45928 -69177 -45902
rect -69473 -46172 -69447 -45928
rect -69447 -46172 -69203 -45928
rect -69203 -46172 -69177 -45928
rect -69473 -46198 -69177 -46172
rect -69133 -46198 -68517 -45902
rect -68473 -45928 -68177 -45902
rect -68473 -46172 -68447 -45928
rect -68447 -46172 -68203 -45928
rect -68203 -46172 -68177 -45928
rect -68473 -46198 -68177 -46172
rect -68133 -46198 -67517 -45902
rect -67473 -45928 -67177 -45902
rect -67473 -46172 -67447 -45928
rect -67447 -46172 -67203 -45928
rect -67203 -46172 -67177 -45928
rect -67473 -46198 -67177 -46172
rect -67133 -46198 -66517 -45902
rect -66473 -45928 -66177 -45902
rect -66473 -46172 -66447 -45928
rect -66447 -46172 -66203 -45928
rect -66203 -46172 -66177 -45928
rect -66473 -46198 -66177 -46172
rect -66133 -46198 -65517 -45902
rect -65473 -45928 -65177 -45902
rect -65473 -46172 -65447 -45928
rect -65447 -46172 -65203 -45928
rect -65203 -46172 -65177 -45928
rect -65473 -46198 -65177 -46172
rect -65133 -46198 -64517 -45902
rect -64473 -45928 -64177 -45902
rect -64473 -46172 -64447 -45928
rect -64447 -46172 -64203 -45928
rect -64203 -46172 -64177 -45928
rect -64473 -46198 -64177 -46172
rect -64133 -46198 -63517 -45902
rect -63473 -45928 -63177 -45902
rect -63473 -46172 -63447 -45928
rect -63447 -46172 -63203 -45928
rect -63203 -46172 -63177 -45928
rect -63473 -46198 -63177 -46172
rect -63133 -46198 -62517 -45902
rect -62473 -45928 -62177 -45902
rect -62473 -46172 -62447 -45928
rect -62447 -46172 -62203 -45928
rect -62203 -46172 -62177 -45928
rect -62473 -46198 -62177 -46172
rect -62133 -46198 -61517 -45902
rect -61473 -45928 -61177 -45902
rect -61473 -46172 -61447 -45928
rect -61447 -46172 -61203 -45928
rect -61203 -46172 -61177 -45928
rect -61473 -46198 -61177 -46172
rect -61133 -46198 -60517 -45902
rect -60473 -45928 -60177 -45902
rect -60473 -46172 -60447 -45928
rect -60447 -46172 -60203 -45928
rect -60203 -46172 -60177 -45928
rect -60473 -46198 -60177 -46172
rect -60133 -46198 -59517 -45902
rect -59473 -45928 -59177 -45902
rect -59473 -46172 -59447 -45928
rect -59447 -46172 -59203 -45928
rect -59203 -46172 -59177 -45928
rect -59473 -46198 -59177 -46172
rect -59133 -46198 -58517 -45902
rect -58473 -45928 -58177 -45902
rect -58473 -46172 -58447 -45928
rect -58447 -46172 -58203 -45928
rect -58203 -46172 -58177 -45928
rect -58473 -46198 -58177 -46172
rect -58133 -46198 -57517 -45902
rect -57473 -45928 -57177 -45902
rect -57473 -46172 -57447 -45928
rect -57447 -46172 -57203 -45928
rect -57203 -46172 -57177 -45928
rect -57473 -46198 -57177 -46172
rect -57133 -46198 -56517 -45902
rect -56473 -45928 -56177 -45902
rect -56473 -46172 -56447 -45928
rect -56447 -46172 -56203 -45928
rect -56203 -46172 -56177 -45928
rect -56473 -46198 -56177 -46172
rect -56133 -46198 -55517 -45902
rect -55473 -45928 -55177 -45902
rect -55473 -46172 -55447 -45928
rect -55447 -46172 -55203 -45928
rect -55203 -46172 -55177 -45928
rect -55473 -46198 -55177 -46172
rect -55133 -46198 -54517 -45902
rect -54473 -45928 -54177 -45902
rect -54473 -46172 -54447 -45928
rect -54447 -46172 -54203 -45928
rect -54203 -46172 -54177 -45928
rect -54473 -46198 -54177 -46172
rect -54133 -46198 -53517 -45902
rect -53473 -45928 -53177 -45902
rect -53473 -46172 -53447 -45928
rect -53447 -46172 -53203 -45928
rect -53203 -46172 -53177 -45928
rect -53473 -46198 -53177 -46172
rect -53133 -46198 -52517 -45902
rect -52473 -45928 -52177 -45902
rect -52473 -46172 -52447 -45928
rect -52447 -46172 -52203 -45928
rect -52203 -46172 -52177 -45928
rect -52473 -46198 -52177 -46172
rect -52133 -46198 -51517 -45902
rect -51473 -45928 -51177 -45902
rect -51473 -46172 -51447 -45928
rect -51447 -46172 -51203 -45928
rect -51203 -46172 -51177 -45928
rect -51473 -46198 -51177 -46172
rect -51133 -46198 -50517 -45902
rect -50473 -45928 -50177 -45902
rect -50473 -46172 -50447 -45928
rect -50447 -46172 -50203 -45928
rect -50203 -46172 -50177 -45928
rect -50473 -46198 -50177 -46172
rect -50133 -46198 -49517 -45902
rect -49473 -45928 -49177 -45902
rect -49473 -46172 -49447 -45928
rect -49447 -46172 -49203 -45928
rect -49203 -46172 -49177 -45928
rect -49473 -46198 -49177 -46172
rect -49133 -46198 -48837 -45902
rect 8287 -46198 8583 -45902
rect 8627 -45928 8923 -45902
rect 8627 -46172 8653 -45928
rect 8653 -46172 8897 -45928
rect 8897 -46172 8923 -45928
rect 8627 -46198 8923 -46172
rect 8967 -46198 9583 -45902
rect 9627 -45928 9923 -45902
rect 9627 -46172 9653 -45928
rect 9653 -46172 9897 -45928
rect 9897 -46172 9923 -45928
rect 9627 -46198 9923 -46172
rect 9967 -46198 10583 -45902
rect 10627 -45928 10923 -45902
rect 10627 -46172 10653 -45928
rect 10653 -46172 10897 -45928
rect 10897 -46172 10923 -45928
rect 10627 -46198 10923 -46172
rect 10967 -46198 11583 -45902
rect 11627 -45928 11923 -45902
rect 11627 -46172 11653 -45928
rect 11653 -46172 11897 -45928
rect 11897 -46172 11923 -45928
rect 11627 -46198 11923 -46172
rect 11967 -46198 12583 -45902
rect 12627 -45928 12923 -45902
rect 12627 -46172 12653 -45928
rect 12653 -46172 12897 -45928
rect 12897 -46172 12923 -45928
rect 12627 -46198 12923 -46172
rect 12967 -46198 13583 -45902
rect 13627 -45928 13923 -45902
rect 13627 -46172 13653 -45928
rect 13653 -46172 13897 -45928
rect 13897 -46172 13923 -45928
rect 13627 -46198 13923 -46172
rect 13967 -46198 14583 -45902
rect 14627 -45928 14923 -45902
rect 14627 -46172 14653 -45928
rect 14653 -46172 14897 -45928
rect 14897 -46172 14923 -45928
rect 14627 -46198 14923 -46172
rect 14967 -46198 15583 -45902
rect 15627 -45928 15923 -45902
rect 15627 -46172 15653 -45928
rect 15653 -46172 15897 -45928
rect 15897 -46172 15923 -45928
rect 15627 -46198 15923 -46172
rect 15967 -46198 16583 -45902
rect 16627 -45928 16923 -45902
rect 16627 -46172 16653 -45928
rect 16653 -46172 16897 -45928
rect 16897 -46172 16923 -45928
rect 16627 -46198 16923 -46172
rect 16967 -46198 17583 -45902
rect 17627 -45928 17923 -45902
rect 17627 -46172 17653 -45928
rect 17653 -46172 17897 -45928
rect 17897 -46172 17923 -45928
rect 17627 -46198 17923 -46172
rect 17967 -46198 18583 -45902
rect 18627 -45928 18923 -45902
rect 18627 -46172 18653 -45928
rect 18653 -46172 18897 -45928
rect 18897 -46172 18923 -45928
rect 18627 -46198 18923 -46172
rect 18967 -46198 19583 -45902
rect 19627 -45928 19923 -45902
rect 19627 -46172 19653 -45928
rect 19653 -46172 19897 -45928
rect 19897 -46172 19923 -45928
rect 19627 -46198 19923 -46172
rect 19967 -46198 20583 -45902
rect 20627 -45928 20923 -45902
rect 20627 -46172 20653 -45928
rect 20653 -46172 20897 -45928
rect 20897 -46172 20923 -45928
rect 20627 -46198 20923 -46172
rect 20967 -46198 21583 -45902
rect 21627 -45928 21923 -45902
rect 21627 -46172 21653 -45928
rect 21653 -46172 21897 -45928
rect 21897 -46172 21923 -45928
rect 21627 -46198 21923 -46172
rect 21967 -46198 22583 -45902
rect 22627 -45928 22923 -45902
rect 22627 -46172 22653 -45928
rect 22653 -46172 22897 -45928
rect 22897 -46172 22923 -45928
rect 22627 -46198 22923 -46172
rect 22967 -46198 23583 -45902
rect 23627 -45928 23923 -45902
rect 23627 -46172 23653 -45928
rect 23653 -46172 23897 -45928
rect 23897 -46172 23923 -45928
rect 23627 -46198 23923 -46172
rect 23967 -46198 24583 -45902
rect 24627 -45928 24923 -45902
rect 24627 -46172 24653 -45928
rect 24653 -46172 24897 -45928
rect 24897 -46172 24923 -45928
rect 24627 -46198 24923 -46172
rect 24967 -46198 25583 -45902
rect 25627 -45928 25923 -45902
rect 25627 -46172 25653 -45928
rect 25653 -46172 25897 -45928
rect 25897 -46172 25923 -45928
rect 25627 -46198 25923 -46172
rect 25967 -46198 26583 -45902
rect 26627 -45928 26923 -45902
rect 26627 -46172 26653 -45928
rect 26653 -46172 26897 -45928
rect 26897 -46172 26923 -45928
rect 26627 -46198 26923 -46172
rect 26967 -46198 27583 -45902
rect 27627 -45928 27923 -45902
rect 27627 -46172 27653 -45928
rect 27653 -46172 27897 -45928
rect 27897 -46172 27923 -45928
rect 27627 -46198 27923 -46172
rect 27967 -46198 28583 -45902
rect 28627 -45928 28923 -45902
rect 28627 -46172 28653 -45928
rect 28653 -46172 28897 -45928
rect 28897 -46172 28923 -45928
rect 28627 -46198 28923 -46172
rect 28967 -46198 29583 -45902
rect 29627 -45928 29923 -45902
rect 29627 -46172 29653 -45928
rect 29653 -46172 29897 -45928
rect 29897 -46172 29923 -45928
rect 29627 -46198 29923 -46172
rect 29967 -46198 30583 -45902
rect 30627 -45928 30923 -45902
rect 30627 -46172 30653 -45928
rect 30653 -46172 30897 -45928
rect 30897 -46172 30923 -45928
rect 30627 -46198 30923 -46172
rect 30967 -46198 31583 -45902
rect 31627 -45928 31923 -45902
rect 31627 -46172 31653 -45928
rect 31653 -46172 31897 -45928
rect 31897 -46172 31923 -45928
rect 31627 -46198 31923 -46172
rect 31967 -46198 32583 -45902
rect 32627 -45928 32923 -45902
rect 32627 -46172 32653 -45928
rect 32653 -46172 32897 -45928
rect 32897 -46172 32923 -45928
rect 32627 -46198 32923 -46172
rect 32967 -46198 33583 -45902
rect 33627 -45928 33923 -45902
rect 33627 -46172 33653 -45928
rect 33653 -46172 33897 -45928
rect 33897 -46172 33923 -45928
rect 33627 -46198 33923 -46172
rect 33967 -46198 34263 -45902
rect -74473 -46538 -74177 -46242
rect -73473 -46538 -73177 -46242
rect -72473 -46538 -72177 -46242
rect -71473 -46538 -71177 -46242
rect -70473 -46538 -70177 -46242
rect -69473 -46538 -69177 -46242
rect -68473 -46538 -68177 -46242
rect -67473 -46538 -67177 -46242
rect -66473 -46538 -66177 -46242
rect -65473 -46538 -65177 -46242
rect -64473 -46538 -64177 -46242
rect -63473 -46538 -63177 -46242
rect -62473 -46538 -62177 -46242
rect -61473 -46538 -61177 -46242
rect -60473 -46538 -60177 -46242
rect -59473 -46538 -59177 -46242
rect -58473 -46538 -58177 -46242
rect -57473 -46538 -57177 -46242
rect -56473 -46538 -56177 -46242
rect -55473 -46538 -55177 -46242
rect -54473 -46538 -54177 -46242
rect -53473 -46538 -53177 -46242
rect -52473 -46538 -52177 -46242
rect -51473 -46538 -51177 -46242
rect -50473 -46538 -50177 -46242
rect -49473 -46538 -49177 -46242
rect 8627 -46538 8923 -46242
rect 9627 -46538 9923 -46242
rect 10627 -46538 10923 -46242
rect 11627 -46538 11923 -46242
rect 12627 -46538 12923 -46242
rect 13627 -46538 13923 -46242
rect 14627 -46538 14923 -46242
rect 15627 -46538 15923 -46242
rect 16627 -46538 16923 -46242
rect 17627 -46538 17923 -46242
rect 18627 -46538 18923 -46242
rect 19627 -46538 19923 -46242
rect 20627 -46538 20923 -46242
rect 21627 -46538 21923 -46242
rect 22627 -46538 22923 -46242
rect 23627 -46538 23923 -46242
rect 24627 -46538 24923 -46242
rect 25627 -46538 25923 -46242
rect 26627 -46538 26923 -46242
rect 27627 -46538 27923 -46242
rect 28627 -46538 28923 -46242
rect 29627 -46538 29923 -46242
rect 30627 -46538 30923 -46242
rect 31627 -46538 31923 -46242
rect 32627 -46538 32923 -46242
rect 33627 -46538 33923 -46242
<< metal3 >>
rect -74485 38542 -74165 38550
rect -74485 38238 -74477 38542
rect -74173 38238 -74165 38542
rect -74485 38210 -74165 38238
rect -73485 38542 -73165 38550
rect -73485 38238 -73477 38542
rect -73173 38238 -73165 38542
rect -73485 38210 -73165 38238
rect -72485 38542 -72165 38550
rect -72485 38238 -72477 38542
rect -72173 38238 -72165 38542
rect -72485 38210 -72165 38238
rect -71485 38542 -71165 38550
rect -71485 38238 -71477 38542
rect -71173 38238 -71165 38542
rect -71485 38210 -71165 38238
rect -70485 38542 -70165 38550
rect -70485 38238 -70477 38542
rect -70173 38238 -70165 38542
rect -70485 38210 -70165 38238
rect -69485 38542 -69165 38550
rect -69485 38238 -69477 38542
rect -69173 38238 -69165 38542
rect -69485 38210 -69165 38238
rect -68485 38542 -68165 38550
rect -68485 38238 -68477 38542
rect -68173 38238 -68165 38542
rect -68485 38210 -68165 38238
rect -67485 38542 -67165 38550
rect -67485 38238 -67477 38542
rect -67173 38238 -67165 38542
rect -67485 38210 -67165 38238
rect -66485 38542 -66165 38550
rect -66485 38238 -66477 38542
rect -66173 38238 -66165 38542
rect -66485 38210 -66165 38238
rect -65485 38542 -65165 38550
rect -65485 38238 -65477 38542
rect -65173 38238 -65165 38542
rect -65485 38210 -65165 38238
rect -64485 38542 -64165 38550
rect -64485 38238 -64477 38542
rect -64173 38238 -64165 38542
rect -64485 38210 -64165 38238
rect -63485 38542 -63165 38550
rect -63485 38238 -63477 38542
rect -63173 38238 -63165 38542
rect -63485 38210 -63165 38238
rect -62485 38542 -62165 38550
rect -62485 38238 -62477 38542
rect -62173 38238 -62165 38542
rect -62485 38210 -62165 38238
rect -61485 38542 -61165 38550
rect -61485 38238 -61477 38542
rect -61173 38238 -61165 38542
rect -61485 38210 -61165 38238
rect -60485 38542 -60165 38550
rect -60485 38238 -60477 38542
rect -60173 38238 -60165 38542
rect -60485 38210 -60165 38238
rect -59485 38542 -59165 38550
rect -59485 38238 -59477 38542
rect -59173 38238 -59165 38542
rect -59485 38210 -59165 38238
rect -74825 38202 -58825 38210
rect -74825 37898 -74817 38202
rect -74513 37898 -74477 38202
rect -74173 37898 -74137 38202
rect -73513 37898 -73477 38202
rect -73173 37898 -73137 38202
rect -72513 37898 -72477 38202
rect -72173 37898 -72137 38202
rect -71513 37898 -71477 38202
rect -71173 37898 -71137 38202
rect -70513 37898 -70477 38202
rect -70173 37898 -70137 38202
rect -69513 37898 -69477 38202
rect -69173 37898 -69137 38202
rect -68513 37898 -68477 38202
rect -68173 37898 -68137 38202
rect -67513 37898 -67477 38202
rect -67173 37898 -67137 38202
rect -66513 37898 -66477 38202
rect -66173 37898 -66137 38202
rect -65513 37898 -65477 38202
rect -65173 37898 -65137 38202
rect -64513 37898 -64477 38202
rect -64173 37898 -64137 38202
rect -63513 37898 -63477 38202
rect -63173 37898 -63137 38202
rect -62513 37898 -62477 38202
rect -62173 37898 -62137 38202
rect -61513 37898 -61477 38202
rect -61173 37898 -61137 38202
rect -60513 37898 -60477 38202
rect -60173 37898 -60137 38202
rect -59513 37898 -59477 38202
rect -59173 37898 -59137 38202
rect -58833 37898 -58825 38202
rect -74825 37890 -58825 37898
rect -74485 37862 -74165 37890
rect -74485 37238 -74477 37862
rect -74173 37238 -74165 37862
rect -74485 37210 -74165 37238
rect -73485 37862 -73165 37890
rect -73485 37238 -73477 37862
rect -73173 37238 -73165 37862
rect -73485 37210 -73165 37238
rect -72485 37862 -72165 37890
rect -72485 37238 -72477 37862
rect -72173 37238 -72165 37862
rect -72485 37210 -72165 37238
rect -71485 37862 -71165 37890
rect -71485 37238 -71477 37862
rect -71173 37238 -71165 37862
rect -71485 37210 -71165 37238
rect -70485 37862 -70165 37890
rect -70485 37238 -70477 37862
rect -70173 37238 -70165 37862
rect -70485 37210 -70165 37238
rect -69485 37862 -69165 37890
rect -69485 37238 -69477 37862
rect -69173 37238 -69165 37862
rect -69485 37210 -69165 37238
rect -68485 37862 -68165 37890
rect -68485 37238 -68477 37862
rect -68173 37238 -68165 37862
rect -68485 37210 -68165 37238
rect -67485 37862 -67165 37890
rect -67485 37238 -67477 37862
rect -67173 37238 -67165 37862
rect -67485 37210 -67165 37238
rect -66485 37862 -66165 37890
rect -66485 37238 -66477 37862
rect -66173 37238 -66165 37862
rect -66485 37210 -66165 37238
rect -65485 37862 -65165 37890
rect -65485 37238 -65477 37862
rect -65173 37238 -65165 37862
rect -65485 37210 -65165 37238
rect -64485 37862 -64165 37890
rect -64485 37238 -64477 37862
rect -64173 37238 -64165 37862
rect -64485 37210 -64165 37238
rect -63485 37862 -63165 37890
rect -63485 37238 -63477 37862
rect -63173 37238 -63165 37862
rect -63485 37210 -63165 37238
rect -62485 37862 -62165 37890
rect -62485 37238 -62477 37862
rect -62173 37238 -62165 37862
rect -62485 37210 -62165 37238
rect -61485 37862 -61165 37890
rect -61485 37238 -61477 37862
rect -61173 37238 -61165 37862
rect -61485 37210 -61165 37238
rect -60485 37862 -60165 37890
rect -60485 37238 -60477 37862
rect -60173 37238 -60165 37862
rect -60485 37210 -60165 37238
rect -59485 37862 -59165 37890
rect -59485 37238 -59477 37862
rect -59173 37238 -59165 37862
rect -59485 37210 -59165 37238
rect -74825 37202 -58825 37210
rect -74825 36898 -74817 37202
rect -74513 36898 -74477 37202
rect -74173 36898 -74137 37202
rect -73513 36898 -73477 37202
rect -73173 36898 -73137 37202
rect -72513 36898 -72477 37202
rect -72173 36898 -72137 37202
rect -71513 36898 -71477 37202
rect -71173 36898 -71137 37202
rect -70513 36898 -70477 37202
rect -70173 36898 -70137 37202
rect -69513 36898 -69477 37202
rect -69173 36898 -69137 37202
rect -68513 36898 -68477 37202
rect -68173 36898 -68137 37202
rect -67513 36898 -67477 37202
rect -67173 36898 -67137 37202
rect -66513 36898 -66477 37202
rect -66173 36898 -66137 37202
rect -65513 36898 -65477 37202
rect -65173 36898 -65137 37202
rect -64513 36898 -64477 37202
rect -64173 36898 -64137 37202
rect -63513 36898 -63477 37202
rect -63173 36898 -63137 37202
rect -62513 36898 -62477 37202
rect -62173 36898 -62137 37202
rect -61513 36898 -61477 37202
rect -61173 36898 -61137 37202
rect -60513 36898 -60477 37202
rect -60173 36898 -60137 37202
rect -59513 36898 -59477 37202
rect -59173 36898 -59137 37202
rect -58833 36898 -58825 37202
rect -74825 36890 -58825 36898
rect -74485 36862 -74165 36890
rect -74485 36238 -74477 36862
rect -74173 36238 -74165 36862
rect -74485 36210 -74165 36238
rect -73485 36862 -73165 36890
rect -73485 36238 -73477 36862
rect -73173 36238 -73165 36862
rect -73485 36210 -73165 36238
rect -72485 36862 -72165 36890
rect -72485 36238 -72477 36862
rect -72173 36238 -72165 36862
rect -72485 36210 -72165 36238
rect -71485 36862 -71165 36890
rect -71485 36238 -71477 36862
rect -71173 36238 -71165 36862
rect -71485 36210 -71165 36238
rect -70485 36862 -70165 36890
rect -70485 36238 -70477 36862
rect -70173 36238 -70165 36862
rect -70485 36210 -70165 36238
rect -69485 36862 -69165 36890
rect -69485 36238 -69477 36862
rect -69173 36238 -69165 36862
rect -69485 36210 -69165 36238
rect -68485 36862 -68165 36890
rect -68485 36238 -68477 36862
rect -68173 36238 -68165 36862
rect -68485 36210 -68165 36238
rect -67485 36862 -67165 36890
rect -67485 36238 -67477 36862
rect -67173 36238 -67165 36862
rect -67485 36210 -67165 36238
rect -66485 36862 -66165 36890
rect -66485 36238 -66477 36862
rect -66173 36238 -66165 36862
rect -66485 36210 -66165 36238
rect -65485 36862 -65165 36890
rect -65485 36238 -65477 36862
rect -65173 36238 -65165 36862
rect -65485 36210 -65165 36238
rect -64485 36862 -64165 36890
rect -64485 36238 -64477 36862
rect -64173 36238 -64165 36862
rect -64485 36210 -64165 36238
rect -63485 36862 -63165 36890
rect -63485 36238 -63477 36862
rect -63173 36238 -63165 36862
rect -63485 36210 -63165 36238
rect -62485 36862 -62165 36890
rect -62485 36238 -62477 36862
rect -62173 36238 -62165 36862
rect -62485 36210 -62165 36238
rect -61485 36862 -61165 36890
rect -61485 36238 -61477 36862
rect -61173 36238 -61165 36862
rect -61485 36210 -61165 36238
rect -60485 36862 -60165 36890
rect -60485 36238 -60477 36862
rect -60173 36238 -60165 36862
rect -60485 36210 -60165 36238
rect -59485 36862 -59165 36890
rect -59485 36238 -59477 36862
rect -59173 36238 -59165 36862
rect -59485 36210 -59165 36238
rect -74825 36202 -58825 36210
rect -74825 35898 -74817 36202
rect -74513 35898 -74477 36202
rect -74173 35898 -74137 36202
rect -73513 35898 -73477 36202
rect -73173 35898 -73137 36202
rect -72513 35898 -72477 36202
rect -72173 35898 -72137 36202
rect -71513 35898 -71477 36202
rect -71173 35898 -71137 36202
rect -70513 35898 -70477 36202
rect -70173 35898 -70137 36202
rect -69513 35898 -69477 36202
rect -69173 35898 -69137 36202
rect -68513 35898 -68477 36202
rect -68173 35898 -68137 36202
rect -67513 35898 -67477 36202
rect -67173 35898 -67137 36202
rect -66513 35898 -66477 36202
rect -66173 35898 -66137 36202
rect -65513 35898 -65477 36202
rect -65173 35898 -65137 36202
rect -64513 35898 -64477 36202
rect -64173 35898 -64137 36202
rect -63513 35898 -63477 36202
rect -63173 35898 -63137 36202
rect -62513 35898 -62477 36202
rect -62173 35898 -62137 36202
rect -61513 35898 -61477 36202
rect -61173 35898 -61137 36202
rect -60513 35898 -60477 36202
rect -60173 35898 -60137 36202
rect -59513 35898 -59477 36202
rect -59173 35898 -59137 36202
rect -58833 35898 -58825 36202
rect -74825 35890 -58825 35898
rect -74485 35862 -74165 35890
rect -74485 35238 -74477 35862
rect -74173 35238 -74165 35862
rect -74485 35210 -74165 35238
rect -73485 35862 -73165 35890
rect -73485 35238 -73477 35862
rect -73173 35238 -73165 35862
rect -73485 35210 -73165 35238
rect -72485 35862 -72165 35890
rect -72485 35238 -72477 35862
rect -72173 35238 -72165 35862
rect -72485 35210 -72165 35238
rect -71485 35862 -71165 35890
rect -71485 35238 -71477 35862
rect -71173 35238 -71165 35862
rect -71485 35210 -71165 35238
rect -70485 35862 -70165 35890
rect -70485 35238 -70477 35862
rect -70173 35238 -70165 35862
rect -70485 35210 -70165 35238
rect -69485 35862 -69165 35890
rect -69485 35238 -69477 35862
rect -69173 35238 -69165 35862
rect -69485 35210 -69165 35238
rect -68485 35862 -68165 35890
rect -68485 35238 -68477 35862
rect -68173 35238 -68165 35862
rect -68485 35210 -68165 35238
rect -67485 35862 -67165 35890
rect -67485 35238 -67477 35862
rect -67173 35238 -67165 35862
rect -67485 35210 -67165 35238
rect -66485 35862 -66165 35890
rect -66485 35238 -66477 35862
rect -66173 35238 -66165 35862
rect -66485 35210 -66165 35238
rect -65485 35862 -65165 35890
rect -65485 35238 -65477 35862
rect -65173 35238 -65165 35862
rect -65485 35210 -65165 35238
rect -64485 35862 -64165 35890
rect -64485 35238 -64477 35862
rect -64173 35238 -64165 35862
rect -64485 35210 -64165 35238
rect -63485 35862 -63165 35890
rect -63485 35238 -63477 35862
rect -63173 35238 -63165 35862
rect -63485 35210 -63165 35238
rect -62485 35862 -62165 35890
rect -62485 35238 -62477 35862
rect -62173 35238 -62165 35862
rect -62485 35210 -62165 35238
rect -61485 35862 -61165 35890
rect -61485 35238 -61477 35862
rect -61173 35238 -61165 35862
rect -61485 35210 -61165 35238
rect -60485 35862 -60165 35890
rect -60485 35238 -60477 35862
rect -60173 35238 -60165 35862
rect -60485 35210 -60165 35238
rect -59485 35862 -59165 35890
rect -59485 35238 -59477 35862
rect -59173 35238 -59165 35862
rect -59485 35210 -59165 35238
rect -74825 35202 -58825 35210
rect -74825 34898 -74817 35202
rect -74513 34898 -74477 35202
rect -74173 34898 -74137 35202
rect -73513 34898 -73477 35202
rect -73173 34898 -73137 35202
rect -72513 34898 -72477 35202
rect -72173 34898 -72137 35202
rect -71513 34898 -71477 35202
rect -71173 34898 -71137 35202
rect -70513 34898 -70477 35202
rect -70173 34898 -70137 35202
rect -69513 34898 -69477 35202
rect -69173 34898 -69137 35202
rect -68513 34898 -68477 35202
rect -68173 34898 -68137 35202
rect -67513 34898 -67477 35202
rect -67173 34898 -67137 35202
rect -66513 34898 -66477 35202
rect -66173 34898 -66137 35202
rect -65513 34898 -65477 35202
rect -65173 34898 -65137 35202
rect -64513 34898 -64477 35202
rect -64173 34898 -64137 35202
rect -63513 34898 -63477 35202
rect -63173 34898 -63137 35202
rect -62513 34898 -62477 35202
rect -62173 34898 -62137 35202
rect -61513 34898 -61477 35202
rect -61173 34898 -61137 35202
rect -60513 34898 -60477 35202
rect -60173 34898 -60137 35202
rect -59513 34898 -59477 35202
rect -59173 34898 -59137 35202
rect -58833 34898 -58825 35202
rect -74825 34890 -58825 34898
rect -74485 34862 -74165 34890
rect -74485 34238 -74477 34862
rect -74173 34238 -74165 34862
rect -74485 34210 -74165 34238
rect -73485 34862 -73165 34890
rect -73485 34238 -73477 34862
rect -73173 34238 -73165 34862
rect -73485 34210 -73165 34238
rect -72485 34862 -72165 34890
rect -72485 34238 -72477 34862
rect -72173 34238 -72165 34862
rect -72485 34210 -72165 34238
rect -71485 34862 -71165 34890
rect -71485 34238 -71477 34862
rect -71173 34238 -71165 34862
rect -71485 34210 -71165 34238
rect -70485 34862 -70165 34890
rect -70485 34238 -70477 34862
rect -70173 34238 -70165 34862
rect -70485 34210 -70165 34238
rect -69485 34862 -69165 34890
rect -69485 34238 -69477 34862
rect -69173 34238 -69165 34862
rect -69485 34210 -69165 34238
rect -68485 34862 -68165 34890
rect -68485 34238 -68477 34862
rect -68173 34238 -68165 34862
rect -68485 34210 -68165 34238
rect -67485 34862 -67165 34890
rect -67485 34238 -67477 34862
rect -67173 34238 -67165 34862
rect -67485 34210 -67165 34238
rect -66485 34862 -66165 34890
rect -66485 34238 -66477 34862
rect -66173 34238 -66165 34862
rect -66485 34210 -66165 34238
rect -65485 34862 -65165 34890
rect -65485 34238 -65477 34862
rect -65173 34238 -65165 34862
rect -65485 34210 -65165 34238
rect -64485 34862 -64165 34890
rect -64485 34238 -64477 34862
rect -64173 34238 -64165 34862
rect -64485 34210 -64165 34238
rect -63485 34862 -63165 34890
rect -63485 34238 -63477 34862
rect -63173 34238 -63165 34862
rect -63485 34210 -63165 34238
rect -62485 34862 -62165 34890
rect -62485 34238 -62477 34862
rect -62173 34238 -62165 34862
rect -62485 34210 -62165 34238
rect -61485 34862 -61165 34890
rect -61485 34238 -61477 34862
rect -61173 34238 -61165 34862
rect -61485 34210 -61165 34238
rect -60485 34862 -60165 34890
rect -60485 34238 -60477 34862
rect -60173 34238 -60165 34862
rect -60485 34210 -60165 34238
rect -59485 34862 -59165 34890
rect -59485 34238 -59477 34862
rect -59173 34238 -59165 34862
rect -59485 34210 -59165 34238
rect -74825 34202 -58825 34210
rect -74825 33898 -74817 34202
rect -74513 33898 -74477 34202
rect -74173 33898 -74137 34202
rect -73513 33898 -73477 34202
rect -73173 33898 -73137 34202
rect -72513 33898 -72477 34202
rect -72173 33898 -72137 34202
rect -71513 33898 -71477 34202
rect -71173 33898 -71137 34202
rect -70513 33898 -70477 34202
rect -70173 33898 -70137 34202
rect -69513 33898 -69477 34202
rect -69173 33898 -69137 34202
rect -68513 33898 -68477 34202
rect -68173 33898 -68137 34202
rect -67513 33898 -67477 34202
rect -67173 33898 -67137 34202
rect -66513 33898 -66477 34202
rect -66173 33898 -66137 34202
rect -65513 33898 -65477 34202
rect -65173 33898 -65137 34202
rect -64513 33898 -64477 34202
rect -64173 33898 -64137 34202
rect -63513 33898 -63477 34202
rect -63173 33898 -63137 34202
rect -62513 33898 -62477 34202
rect -62173 33898 -62137 34202
rect -61513 33898 -61477 34202
rect -61173 33898 -61137 34202
rect -60513 33898 -60477 34202
rect -60173 33898 -60137 34202
rect -59513 33898 -59477 34202
rect -59173 33898 -59137 34202
rect -58833 33898 -58825 34202
rect -74825 33890 -58825 33898
rect -74485 33862 -74165 33890
rect -74485 33238 -74477 33862
rect -74173 33238 -74165 33862
rect -74485 33210 -74165 33238
rect -73485 33862 -73165 33890
rect -73485 33238 -73477 33862
rect -73173 33238 -73165 33862
rect -73485 33210 -73165 33238
rect -72485 33862 -72165 33890
rect -72485 33238 -72477 33862
rect -72173 33238 -72165 33862
rect -72485 33210 -72165 33238
rect -71485 33862 -71165 33890
rect -71485 33238 -71477 33862
rect -71173 33238 -71165 33862
rect -71485 33210 -71165 33238
rect -70485 33862 -70165 33890
rect -70485 33238 -70477 33862
rect -70173 33238 -70165 33862
rect -70485 33210 -70165 33238
rect -69485 33862 -69165 33890
rect -69485 33238 -69477 33862
rect -69173 33238 -69165 33862
rect -69485 33210 -69165 33238
rect -68485 33862 -68165 33890
rect -68485 33238 -68477 33862
rect -68173 33238 -68165 33862
rect -68485 33210 -68165 33238
rect -67485 33862 -67165 33890
rect -67485 33238 -67477 33862
rect -67173 33238 -67165 33862
rect -67485 33210 -67165 33238
rect -66485 33862 -66165 33890
rect -66485 33238 -66477 33862
rect -66173 33238 -66165 33862
rect -66485 33210 -66165 33238
rect -65485 33862 -65165 33890
rect -65485 33238 -65477 33862
rect -65173 33238 -65165 33862
rect -65485 33210 -65165 33238
rect -64485 33862 -64165 33890
rect -64485 33238 -64477 33862
rect -64173 33238 -64165 33862
rect -64485 33210 -64165 33238
rect -63485 33862 -63165 33890
rect -63485 33238 -63477 33862
rect -63173 33238 -63165 33862
rect -63485 33210 -63165 33238
rect -62485 33862 -62165 33890
rect -62485 33238 -62477 33862
rect -62173 33238 -62165 33862
rect -62485 33210 -62165 33238
rect -61485 33862 -61165 33890
rect -61485 33238 -61477 33862
rect -61173 33238 -61165 33862
rect -61485 33210 -61165 33238
rect -60485 33862 -60165 33890
rect -60485 33238 -60477 33862
rect -60173 33238 -60165 33862
rect -60485 33210 -60165 33238
rect -59485 33862 -59165 33890
rect -59485 33238 -59477 33862
rect -59173 33238 -59165 33862
rect -59485 33210 -59165 33238
rect -74825 33202 -58825 33210
rect -74825 32898 -74817 33202
rect -74513 32898 -74477 33202
rect -74173 32898 -74137 33202
rect -73513 32898 -73477 33202
rect -73173 32898 -73137 33202
rect -72513 32898 -72477 33202
rect -72173 32898 -72137 33202
rect -71513 32898 -71477 33202
rect -71173 32898 -71137 33202
rect -70513 32898 -70477 33202
rect -70173 32898 -70137 33202
rect -69513 32898 -69477 33202
rect -69173 32898 -69137 33202
rect -68513 32898 -68477 33202
rect -68173 32898 -68137 33202
rect -67513 32898 -67477 33202
rect -67173 32898 -67137 33202
rect -66513 32898 -66477 33202
rect -66173 32898 -66137 33202
rect -65513 32898 -65477 33202
rect -65173 32898 -65137 33202
rect -64513 32898 -64477 33202
rect -64173 32898 -64137 33202
rect -63513 32898 -63477 33202
rect -63173 32898 -63137 33202
rect -62513 32898 -62477 33202
rect -62173 32898 -62137 33202
rect -61513 32898 -61477 33202
rect -61173 32898 -61137 33202
rect -60513 32898 -60477 33202
rect -60173 32898 -60137 33202
rect -59513 32898 -59477 33202
rect -59173 32898 -59137 33202
rect -58833 32898 -58825 33202
rect -74825 32890 -58825 32898
rect -57352 33076 -56752 48242
rect -27789 40573 -12989 47031
rect -50437 36573 4504 40573
rect 16011 38550 30811 47031
rect 9994 38542 10314 38550
rect 9994 38238 10002 38542
rect 10306 38238 10314 38542
rect 9994 38210 10314 38238
rect 10994 38542 11314 38550
rect 10994 38238 11002 38542
rect 11306 38238 11314 38542
rect 10994 38210 11314 38238
rect 11994 38542 12314 38550
rect 11994 38238 12002 38542
rect 12306 38238 12314 38542
rect 11994 38210 12314 38238
rect 12994 38542 13314 38550
rect 12994 38238 13002 38542
rect 13306 38238 13314 38542
rect 12994 38210 13314 38238
rect 13994 38542 14314 38550
rect 13994 38238 14002 38542
rect 14306 38238 14314 38542
rect 13994 38210 14314 38238
rect 14994 38542 32314 38550
rect 14994 38238 15002 38542
rect 15306 38238 16002 38542
rect 16306 38238 17002 38542
rect 17306 38238 18002 38542
rect 18306 38238 19002 38542
rect 19306 38238 20002 38542
rect 20306 38238 21002 38542
rect 21306 38238 22002 38542
rect 22306 38238 23002 38542
rect 23306 38238 24002 38542
rect 24306 38238 25002 38542
rect 25306 38238 26002 38542
rect 26306 38238 27002 38542
rect 27306 38238 28002 38542
rect 28306 38238 29002 38542
rect 29306 38238 30002 38542
rect 30306 38238 31002 38542
rect 31306 38238 32002 38542
rect 32306 38238 32314 38542
rect 14994 38210 32314 38238
rect 32994 38542 33314 38550
rect 32994 38238 33002 38542
rect 33306 38238 33314 38542
rect 32994 38210 33314 38238
rect 33994 38542 34314 38550
rect 33994 38238 34002 38542
rect 34306 38238 34314 38542
rect 33994 38210 34314 38238
rect 9654 38202 34654 38210
rect 9654 37898 9662 38202
rect 9966 37898 10002 38202
rect 10306 37898 10342 38202
rect 10966 37898 11002 38202
rect 11306 37898 11342 38202
rect 11966 37898 12002 38202
rect 12306 37898 12342 38202
rect 12966 37898 13002 38202
rect 13306 37898 13342 38202
rect 13966 37898 14002 38202
rect 14306 37898 14342 38202
rect 14966 37898 15002 38202
rect 15306 37898 15342 38202
rect 15966 37898 16002 38202
rect 16306 37898 16342 38202
rect 16966 37898 17002 38202
rect 17306 37898 17342 38202
rect 17966 37898 18002 38202
rect 18306 37898 18342 38202
rect 18966 37898 19002 38202
rect 19306 37898 19342 38202
rect 19966 37898 20002 38202
rect 20306 37898 20342 38202
rect 20966 37898 21002 38202
rect 21306 37898 21342 38202
rect 21966 37898 22002 38202
rect 22306 37898 22342 38202
rect 22966 37898 23002 38202
rect 23306 37898 23342 38202
rect 23966 37898 24002 38202
rect 24306 37898 24342 38202
rect 24966 37898 25002 38202
rect 25306 37898 25342 38202
rect 25966 37898 26002 38202
rect 26306 37898 26342 38202
rect 26966 37898 27002 38202
rect 27306 37898 27342 38202
rect 27966 37898 28002 38202
rect 28306 37898 28342 38202
rect 28966 37898 29002 38202
rect 29306 37898 29342 38202
rect 29966 37898 30002 38202
rect 30306 37898 30342 38202
rect 30966 37898 31002 38202
rect 31306 37898 31342 38202
rect 31966 37898 32002 38202
rect 32306 37898 32342 38202
rect 32966 37898 33002 38202
rect 33306 37898 33342 38202
rect 33966 37898 34002 38202
rect 34306 37898 34342 38202
rect 34646 37898 34654 38202
rect 9654 37890 34654 37898
rect 9994 37862 10314 37890
rect 9994 37238 10002 37862
rect 10306 37238 10314 37862
rect 9994 37210 10314 37238
rect 10994 37862 11314 37890
rect 10994 37238 11002 37862
rect 11306 37238 11314 37862
rect 10994 37210 11314 37238
rect 11994 37862 12314 37890
rect 11994 37238 12002 37862
rect 12306 37238 12314 37862
rect 11994 37210 12314 37238
rect 12994 37862 13314 37890
rect 12994 37238 13002 37862
rect 13306 37238 13314 37862
rect 12994 37210 13314 37238
rect 13994 37862 14314 37890
rect 13994 37238 14002 37862
rect 14306 37238 14314 37862
rect 13994 37210 14314 37238
rect 14994 37862 15314 37890
rect 14994 37238 15002 37862
rect 15306 37238 15314 37862
rect 14994 37210 15314 37238
rect 15994 37862 16314 37890
rect 15994 37238 16002 37862
rect 16306 37238 16314 37862
rect 15994 37210 16314 37238
rect 16994 37862 17314 37890
rect 16994 37238 17002 37862
rect 17306 37238 17314 37862
rect 16994 37210 17314 37238
rect 17994 37862 18314 37890
rect 17994 37238 18002 37862
rect 18306 37238 18314 37862
rect 17994 37210 18314 37238
rect 18994 37862 19314 37890
rect 18994 37238 19002 37862
rect 19306 37238 19314 37862
rect 18994 37210 19314 37238
rect 19994 37862 20314 37890
rect 19994 37238 20002 37862
rect 20306 37238 20314 37862
rect 19994 37210 20314 37238
rect 20994 37862 21314 37890
rect 20994 37238 21002 37862
rect 21306 37238 21314 37862
rect 20994 37210 21314 37238
rect 21994 37862 22314 37890
rect 21994 37238 22002 37862
rect 22306 37238 22314 37862
rect 21994 37210 22314 37238
rect 22994 37862 23314 37890
rect 22994 37238 23002 37862
rect 23306 37238 23314 37862
rect 22994 37210 23314 37238
rect 23994 37862 24314 37890
rect 23994 37238 24002 37862
rect 24306 37238 24314 37862
rect 23994 37210 24314 37238
rect 24994 37862 25314 37890
rect 24994 37238 25002 37862
rect 25306 37238 25314 37862
rect 24994 37210 25314 37238
rect 25994 37862 26314 37890
rect 25994 37238 26002 37862
rect 26306 37238 26314 37862
rect 25994 37210 26314 37238
rect 26994 37862 27314 37890
rect 26994 37238 27002 37862
rect 27306 37238 27314 37862
rect 26994 37210 27314 37238
rect 27994 37862 28314 37890
rect 27994 37238 28002 37862
rect 28306 37238 28314 37862
rect 27994 37210 28314 37238
rect 28994 37862 29314 37890
rect 28994 37238 29002 37862
rect 29306 37238 29314 37862
rect 28994 37210 29314 37238
rect 29994 37862 30314 37890
rect 29994 37238 30002 37862
rect 30306 37238 30314 37862
rect 29994 37210 30314 37238
rect 30994 37862 31314 37890
rect 30994 37238 31002 37862
rect 31306 37238 31314 37862
rect 30994 37210 31314 37238
rect 31994 37862 32314 37890
rect 31994 37238 32002 37862
rect 32306 37238 32314 37862
rect 31994 37210 32314 37238
rect 32994 37862 33314 37890
rect 32994 37238 33002 37862
rect 33306 37238 33314 37862
rect 32994 37210 33314 37238
rect 33994 37862 34314 37890
rect 33994 37238 34002 37862
rect 34306 37238 34314 37862
rect 33994 37210 34314 37238
rect 9654 37202 34654 37210
rect 9654 36898 9662 37202
rect 9966 36898 10002 37202
rect 10306 36898 10342 37202
rect 10966 36898 11002 37202
rect 11306 36898 11342 37202
rect 11966 36898 12002 37202
rect 12306 36898 12342 37202
rect 12966 36898 13002 37202
rect 13306 36898 13342 37202
rect 13966 36898 14002 37202
rect 14306 36898 14342 37202
rect 14966 36898 15002 37202
rect 15306 36898 15342 37202
rect 15966 36898 16002 37202
rect 16306 36898 16342 37202
rect 16966 36898 17002 37202
rect 17306 36898 17342 37202
rect 17966 36898 18002 37202
rect 18306 36898 18342 37202
rect 18966 36898 19002 37202
rect 19306 36898 19342 37202
rect 19966 36898 20002 37202
rect 20306 36898 20342 37202
rect 20966 36898 21002 37202
rect 21306 36898 21342 37202
rect 21966 36898 22002 37202
rect 22306 36898 22342 37202
rect 22966 36898 23002 37202
rect 23306 36898 23342 37202
rect 23966 36898 24002 37202
rect 24306 36898 24342 37202
rect 24966 36898 25002 37202
rect 25306 36898 25342 37202
rect 25966 36898 26002 37202
rect 26306 36898 26342 37202
rect 26966 36898 27002 37202
rect 27306 36898 27342 37202
rect 27966 36898 28002 37202
rect 28306 36898 28342 37202
rect 28966 36898 29002 37202
rect 29306 36898 29342 37202
rect 29966 36898 30002 37202
rect 30306 36898 30342 37202
rect 30966 36898 31002 37202
rect 31306 36898 31342 37202
rect 31966 36898 32002 37202
rect 32306 36898 32342 37202
rect 32966 36898 33002 37202
rect 33306 36898 33342 37202
rect 33966 36898 34002 37202
rect 34306 36898 34342 37202
rect 34646 36898 34654 37202
rect 9654 36890 34654 36898
rect -50437 34164 -48843 36573
rect -50437 33548 -50428 34164
rect -48852 33548 -48843 34164
rect -50437 33539 -48843 33548
rect 2910 34164 4504 36573
rect 9994 36862 10314 36890
rect 9994 36238 10002 36862
rect 10306 36238 10314 36862
rect 9994 36210 10314 36238
rect 10994 36862 11314 36890
rect 10994 36238 11002 36862
rect 11306 36238 11314 36862
rect 10994 36210 11314 36238
rect 11994 36862 12314 36890
rect 11994 36238 12002 36862
rect 12306 36238 12314 36862
rect 11994 36210 12314 36238
rect 12994 36862 13314 36890
rect 12994 36238 13002 36862
rect 13306 36238 13314 36862
rect 12994 36210 13314 36238
rect 13994 36862 14314 36890
rect 13994 36238 14002 36862
rect 14306 36238 14314 36862
rect 13994 36210 14314 36238
rect 14994 36862 15314 36890
rect 14994 36238 15002 36862
rect 15306 36238 15314 36862
rect 14994 36210 15314 36238
rect 15994 36862 16314 36890
rect 15994 36238 16002 36862
rect 16306 36238 16314 36862
rect 15994 36210 16314 36238
rect 16994 36862 17314 36890
rect 16994 36238 17002 36862
rect 17306 36238 17314 36862
rect 16994 36210 17314 36238
rect 17994 36862 18314 36890
rect 17994 36238 18002 36862
rect 18306 36238 18314 36862
rect 17994 36210 18314 36238
rect 18994 36862 19314 36890
rect 18994 36238 19002 36862
rect 19306 36238 19314 36862
rect 18994 36210 19314 36238
rect 19994 36862 20314 36890
rect 19994 36238 20002 36862
rect 20306 36238 20314 36862
rect 19994 36210 20314 36238
rect 20994 36862 21314 36890
rect 20994 36238 21002 36862
rect 21306 36238 21314 36862
rect 20994 36210 21314 36238
rect 21994 36862 22314 36890
rect 21994 36238 22002 36862
rect 22306 36238 22314 36862
rect 21994 36210 22314 36238
rect 22994 36862 23314 36890
rect 22994 36238 23002 36862
rect 23306 36238 23314 36862
rect 22994 36210 23314 36238
rect 23994 36862 24314 36890
rect 23994 36238 24002 36862
rect 24306 36238 24314 36862
rect 23994 36210 24314 36238
rect 24994 36862 25314 36890
rect 24994 36238 25002 36862
rect 25306 36238 25314 36862
rect 24994 36210 25314 36238
rect 25994 36862 26314 36890
rect 25994 36238 26002 36862
rect 26306 36238 26314 36862
rect 25994 36210 26314 36238
rect 26994 36862 27314 36890
rect 26994 36238 27002 36862
rect 27306 36238 27314 36862
rect 26994 36210 27314 36238
rect 27994 36862 28314 36890
rect 27994 36238 28002 36862
rect 28306 36238 28314 36862
rect 27994 36210 28314 36238
rect 28994 36862 29314 36890
rect 28994 36238 29002 36862
rect 29306 36238 29314 36862
rect 28994 36210 29314 36238
rect 29994 36862 30314 36890
rect 29994 36238 30002 36862
rect 30306 36238 30314 36862
rect 29994 36210 30314 36238
rect 30994 36862 31314 36890
rect 30994 36238 31002 36862
rect 31306 36238 31314 36862
rect 30994 36210 31314 36238
rect 31994 36862 32314 36890
rect 31994 36238 32002 36862
rect 32306 36238 32314 36862
rect 31994 36210 32314 36238
rect 32994 36862 33314 36890
rect 32994 36238 33002 36862
rect 33306 36238 33314 36862
rect 32994 36210 33314 36238
rect 33994 36862 34314 36890
rect 33994 36238 34002 36862
rect 34306 36238 34314 36862
rect 33994 36210 34314 36238
rect 9654 36202 34654 36210
rect 9654 35898 9662 36202
rect 9966 35898 10002 36202
rect 10306 35898 10342 36202
rect 10966 35898 11002 36202
rect 11306 35898 11342 36202
rect 11966 35898 12002 36202
rect 12306 35898 12342 36202
rect 12966 35898 13002 36202
rect 13306 35898 13342 36202
rect 13966 35898 14002 36202
rect 14306 35898 14342 36202
rect 14966 35898 15002 36202
rect 15306 35898 15342 36202
rect 15966 35898 16002 36202
rect 16306 35898 16342 36202
rect 16966 35898 17002 36202
rect 17306 35898 17342 36202
rect 17966 35898 18002 36202
rect 18306 35898 18342 36202
rect 18966 35898 19002 36202
rect 19306 35898 19342 36202
rect 19966 35898 20002 36202
rect 20306 35898 20342 36202
rect 20966 35898 21002 36202
rect 21306 35898 21342 36202
rect 21966 35898 22002 36202
rect 22306 35898 22342 36202
rect 22966 35898 23002 36202
rect 23306 35898 23342 36202
rect 23966 35898 24002 36202
rect 24306 35898 24342 36202
rect 24966 35898 25002 36202
rect 25306 35898 25342 36202
rect 25966 35898 26002 36202
rect 26306 35898 26342 36202
rect 26966 35898 27002 36202
rect 27306 35898 27342 36202
rect 27966 35898 28002 36202
rect 28306 35898 28342 36202
rect 28966 35898 29002 36202
rect 29306 35898 29342 36202
rect 29966 35898 30002 36202
rect 30306 35898 30342 36202
rect 30966 35898 31002 36202
rect 31306 35898 31342 36202
rect 31966 35898 32002 36202
rect 32306 35898 32342 36202
rect 32966 35898 33002 36202
rect 33306 35898 33342 36202
rect 33966 35898 34002 36202
rect 34306 35898 34342 36202
rect 34646 35898 34654 36202
rect 9654 35890 34654 35898
rect 9994 35862 10314 35890
rect 9994 35238 10002 35862
rect 10306 35238 10314 35862
rect 9994 35210 10314 35238
rect 10994 35862 11314 35890
rect 10994 35238 11002 35862
rect 11306 35238 11314 35862
rect 10994 35210 11314 35238
rect 11994 35862 12314 35890
rect 11994 35238 12002 35862
rect 12306 35238 12314 35862
rect 11994 35210 12314 35238
rect 12994 35862 13314 35890
rect 12994 35238 13002 35862
rect 13306 35238 13314 35862
rect 12994 35210 13314 35238
rect 13994 35862 14314 35890
rect 13994 35238 14002 35862
rect 14306 35238 14314 35862
rect 13994 35210 14314 35238
rect 14994 35862 15314 35890
rect 14994 35238 15002 35862
rect 15306 35238 15314 35862
rect 14994 35210 15314 35238
rect 15994 35862 16314 35890
rect 15994 35238 16002 35862
rect 16306 35238 16314 35862
rect 15994 35210 16314 35238
rect 16994 35862 17314 35890
rect 16994 35238 17002 35862
rect 17306 35238 17314 35862
rect 16994 35210 17314 35238
rect 17994 35862 18314 35890
rect 17994 35238 18002 35862
rect 18306 35238 18314 35862
rect 17994 35210 18314 35238
rect 18994 35862 19314 35890
rect 18994 35238 19002 35862
rect 19306 35238 19314 35862
rect 18994 35210 19314 35238
rect 19994 35862 20314 35890
rect 19994 35238 20002 35862
rect 20306 35238 20314 35862
rect 19994 35210 20314 35238
rect 20994 35862 21314 35890
rect 20994 35238 21002 35862
rect 21306 35238 21314 35862
rect 20994 35210 21314 35238
rect 21994 35862 22314 35890
rect 21994 35238 22002 35862
rect 22306 35238 22314 35862
rect 21994 35210 22314 35238
rect 22994 35862 23314 35890
rect 22994 35238 23002 35862
rect 23306 35238 23314 35862
rect 22994 35210 23314 35238
rect 23994 35862 24314 35890
rect 23994 35238 24002 35862
rect 24306 35238 24314 35862
rect 23994 35210 24314 35238
rect 24994 35862 25314 35890
rect 24994 35238 25002 35862
rect 25306 35238 25314 35862
rect 24994 35210 25314 35238
rect 25994 35862 26314 35890
rect 25994 35238 26002 35862
rect 26306 35238 26314 35862
rect 25994 35210 26314 35238
rect 26994 35862 27314 35890
rect 26994 35238 27002 35862
rect 27306 35238 27314 35862
rect 26994 35210 27314 35238
rect 27994 35862 28314 35890
rect 27994 35238 28002 35862
rect 28306 35238 28314 35862
rect 27994 35210 28314 35238
rect 28994 35862 29314 35890
rect 28994 35238 29002 35862
rect 29306 35238 29314 35862
rect 28994 35210 29314 35238
rect 29994 35862 30314 35890
rect 29994 35238 30002 35862
rect 30306 35238 30314 35862
rect 29994 35210 30314 35238
rect 30994 35862 31314 35890
rect 30994 35238 31002 35862
rect 31306 35238 31314 35862
rect 30994 35210 31314 35238
rect 31994 35862 32314 35890
rect 31994 35238 32002 35862
rect 32306 35238 32314 35862
rect 31994 35210 32314 35238
rect 32994 35862 33314 35890
rect 32994 35238 33002 35862
rect 33306 35238 33314 35862
rect 32994 35210 33314 35238
rect 33994 35862 34314 35890
rect 33994 35238 34002 35862
rect 34306 35238 34314 35862
rect 33994 35210 34314 35238
rect 9654 35202 34654 35210
rect 9654 34898 9662 35202
rect 9966 34898 10002 35202
rect 10306 34898 10342 35202
rect 10966 34898 11002 35202
rect 11306 34898 11342 35202
rect 11966 34898 12002 35202
rect 12306 34898 12342 35202
rect 12966 34898 13002 35202
rect 13306 34898 13342 35202
rect 13966 34898 14002 35202
rect 14306 34898 14342 35202
rect 14966 34898 15002 35202
rect 15306 34898 15342 35202
rect 15966 34898 16002 35202
rect 16306 34898 16342 35202
rect 16966 34898 17002 35202
rect 17306 34898 17342 35202
rect 17966 34898 18002 35202
rect 18306 34898 18342 35202
rect 18966 34898 19002 35202
rect 19306 34898 19342 35202
rect 19966 34898 20002 35202
rect 20306 34898 20342 35202
rect 20966 34898 21002 35202
rect 21306 34898 21342 35202
rect 21966 34898 22002 35202
rect 22306 34898 22342 35202
rect 22966 34898 23002 35202
rect 23306 34898 23342 35202
rect 23966 34898 24002 35202
rect 24306 34898 24342 35202
rect 24966 34898 25002 35202
rect 25306 34898 25342 35202
rect 25966 34898 26002 35202
rect 26306 34898 26342 35202
rect 26966 34898 27002 35202
rect 27306 34898 27342 35202
rect 27966 34898 28002 35202
rect 28306 34898 28342 35202
rect 28966 34898 29002 35202
rect 29306 34898 29342 35202
rect 29966 34898 30002 35202
rect 30306 34898 30342 35202
rect 30966 34898 31002 35202
rect 31306 34898 31342 35202
rect 31966 34898 32002 35202
rect 32306 34898 32342 35202
rect 32966 34898 33002 35202
rect 33306 34898 33342 35202
rect 33966 34898 34002 35202
rect 34306 34898 34342 35202
rect 34646 34898 34654 35202
rect 9654 34890 34654 34898
rect 9994 34862 10314 34890
rect 9994 34238 10002 34862
rect 10306 34238 10314 34862
rect 9994 34210 10314 34238
rect 10994 34862 11314 34890
rect 10994 34238 11002 34862
rect 11306 34238 11314 34862
rect 10994 34210 11314 34238
rect 11994 34862 12314 34890
rect 11994 34238 12002 34862
rect 12306 34238 12314 34862
rect 11994 34210 12314 34238
rect 12994 34862 13314 34890
rect 12994 34238 13002 34862
rect 13306 34238 13314 34862
rect 12994 34210 13314 34238
rect 13994 34862 14314 34890
rect 13994 34238 14002 34862
rect 14306 34238 14314 34862
rect 13994 34210 14314 34238
rect 14994 34862 15314 34890
rect 14994 34238 15002 34862
rect 15306 34238 15314 34862
rect 14994 34210 15314 34238
rect 15994 34862 16314 34890
rect 15994 34238 16002 34862
rect 16306 34238 16314 34862
rect 15994 34210 16314 34238
rect 16994 34862 17314 34890
rect 16994 34238 17002 34862
rect 17306 34238 17314 34862
rect 16994 34210 17314 34238
rect 17994 34862 18314 34890
rect 17994 34238 18002 34862
rect 18306 34238 18314 34862
rect 17994 34210 18314 34238
rect 18994 34862 19314 34890
rect 18994 34238 19002 34862
rect 19306 34238 19314 34862
rect 18994 34210 19314 34238
rect 19994 34862 20314 34890
rect 19994 34238 20002 34862
rect 20306 34238 20314 34862
rect 19994 34210 20314 34238
rect 20994 34862 21314 34890
rect 20994 34238 21002 34862
rect 21306 34238 21314 34862
rect 20994 34210 21314 34238
rect 21994 34862 22314 34890
rect 21994 34238 22002 34862
rect 22306 34238 22314 34862
rect 21994 34210 22314 34238
rect 22994 34862 23314 34890
rect 22994 34238 23002 34862
rect 23306 34238 23314 34862
rect 22994 34210 23314 34238
rect 23994 34862 24314 34890
rect 23994 34238 24002 34862
rect 24306 34238 24314 34862
rect 23994 34210 24314 34238
rect 24994 34862 25314 34890
rect 24994 34238 25002 34862
rect 25306 34238 25314 34862
rect 24994 34210 25314 34238
rect 25994 34862 26314 34890
rect 25994 34238 26002 34862
rect 26306 34238 26314 34862
rect 25994 34210 26314 34238
rect 26994 34862 27314 34890
rect 26994 34238 27002 34862
rect 27306 34238 27314 34862
rect 26994 34210 27314 34238
rect 27994 34862 28314 34890
rect 27994 34238 28002 34862
rect 28306 34238 28314 34862
rect 27994 34210 28314 34238
rect 28994 34862 29314 34890
rect 28994 34238 29002 34862
rect 29306 34238 29314 34862
rect 28994 34210 29314 34238
rect 29994 34862 30314 34890
rect 29994 34238 30002 34862
rect 30306 34238 30314 34862
rect 29994 34210 30314 34238
rect 30994 34862 31314 34890
rect 30994 34238 31002 34862
rect 31306 34238 31314 34862
rect 30994 34210 31314 34238
rect 31994 34862 32314 34890
rect 31994 34238 32002 34862
rect 32306 34238 32314 34862
rect 31994 34210 32314 34238
rect 32994 34862 33314 34890
rect 32994 34238 33002 34862
rect 33306 34238 33314 34862
rect 32994 34210 33314 34238
rect 33994 34862 34314 34890
rect 33994 34238 34002 34862
rect 34306 34238 34314 34862
rect 33994 34210 34314 34238
rect 2910 33548 2919 34164
rect 4495 33548 4504 34164
rect 9654 34202 34654 34210
rect 9654 33898 9662 34202
rect 9966 33898 10002 34202
rect 10306 33898 10342 34202
rect 10966 33898 11002 34202
rect 11306 33898 11342 34202
rect 11966 33898 12002 34202
rect 12306 33898 12342 34202
rect 12966 33898 13002 34202
rect 13306 33898 13342 34202
rect 13966 33898 14002 34202
rect 14306 33898 14342 34202
rect 14966 33898 15002 34202
rect 15306 33898 15342 34202
rect 15966 33898 16002 34202
rect 16306 33898 16342 34202
rect 16966 33898 17002 34202
rect 17306 33898 17342 34202
rect 17966 33898 18002 34202
rect 18306 33898 18342 34202
rect 18966 33898 19002 34202
rect 19306 33898 19342 34202
rect 19966 33898 20002 34202
rect 20306 33898 20342 34202
rect 20966 33898 21002 34202
rect 21306 33898 21342 34202
rect 21966 33898 22002 34202
rect 22306 33898 22342 34202
rect 22966 33898 23002 34202
rect 23306 33898 23342 34202
rect 23966 33898 24002 34202
rect 24306 33898 24342 34202
rect 24966 33898 25002 34202
rect 25306 33898 25342 34202
rect 25966 33898 26002 34202
rect 26306 33898 26342 34202
rect 26966 33898 27002 34202
rect 27306 33898 27342 34202
rect 27966 33898 28002 34202
rect 28306 33898 28342 34202
rect 28966 33898 29002 34202
rect 29306 33898 29342 34202
rect 29966 33898 30002 34202
rect 30306 33898 30342 34202
rect 30966 33898 31002 34202
rect 31306 33898 31342 34202
rect 31966 33898 32002 34202
rect 32306 33898 32342 34202
rect 32966 33898 33002 34202
rect 33306 33898 33342 34202
rect 33966 33898 34002 34202
rect 34306 33898 34342 34202
rect 34646 33898 34654 34202
rect 9654 33890 34654 33898
rect 2910 33539 4504 33548
rect 9994 33862 10314 33890
rect 9994 33238 10002 33862
rect 10306 33238 10314 33862
rect 9994 33210 10314 33238
rect 10994 33862 11314 33890
rect 10994 33238 11002 33862
rect 11306 33238 11314 33862
rect 10994 33210 11314 33238
rect 11994 33862 12314 33890
rect 11994 33238 12002 33862
rect 12306 33238 12314 33862
rect 11994 33210 12314 33238
rect 12994 33862 13314 33890
rect 12994 33238 13002 33862
rect 13306 33238 13314 33862
rect 12994 33210 13314 33238
rect 13994 33862 14314 33890
rect 13994 33238 14002 33862
rect 14306 33238 14314 33862
rect 13994 33210 14314 33238
rect 14994 33862 15314 33890
rect 14994 33238 15002 33862
rect 15306 33238 15314 33862
rect 14994 33210 15314 33238
rect 15994 33862 16314 33890
rect 15994 33238 16002 33862
rect 16306 33238 16314 33862
rect 15994 33210 16314 33238
rect 16994 33862 17314 33890
rect 16994 33238 17002 33862
rect 17306 33238 17314 33862
rect 16994 33210 17314 33238
rect 17994 33862 18314 33890
rect 17994 33238 18002 33862
rect 18306 33238 18314 33862
rect 17994 33210 18314 33238
rect 18994 33862 19314 33890
rect 18994 33238 19002 33862
rect 19306 33238 19314 33862
rect 18994 33210 19314 33238
rect 19994 33862 20314 33890
rect 19994 33238 20002 33862
rect 20306 33238 20314 33862
rect 19994 33210 20314 33238
rect 20994 33862 21314 33890
rect 20994 33238 21002 33862
rect 21306 33238 21314 33862
rect 20994 33210 21314 33238
rect 21994 33862 22314 33890
rect 21994 33238 22002 33862
rect 22306 33238 22314 33862
rect 21994 33210 22314 33238
rect 22994 33862 23314 33890
rect 22994 33238 23002 33862
rect 23306 33238 23314 33862
rect 22994 33210 23314 33238
rect 23994 33862 24314 33890
rect 23994 33238 24002 33862
rect 24306 33238 24314 33862
rect 23994 33210 24314 33238
rect 24994 33862 25314 33890
rect 24994 33238 25002 33862
rect 25306 33238 25314 33862
rect 24994 33210 25314 33238
rect 25994 33862 26314 33890
rect 25994 33238 26002 33862
rect 26306 33238 26314 33862
rect 25994 33210 26314 33238
rect 26994 33862 27314 33890
rect 26994 33238 27002 33862
rect 27306 33238 27314 33862
rect 26994 33210 27314 33238
rect 27994 33862 28314 33890
rect 27994 33238 28002 33862
rect 28306 33238 28314 33862
rect 27994 33210 28314 33238
rect 28994 33862 29314 33890
rect 28994 33238 29002 33862
rect 29306 33238 29314 33862
rect 28994 33210 29314 33238
rect 29994 33862 30314 33890
rect 29994 33238 30002 33862
rect 30306 33238 30314 33862
rect 29994 33210 30314 33238
rect 30994 33862 31314 33890
rect 30994 33238 31002 33862
rect 31306 33238 31314 33862
rect 30994 33210 31314 33238
rect 31994 33862 32314 33890
rect 31994 33238 32002 33862
rect 32306 33238 32314 33862
rect 31994 33210 32314 33238
rect 32994 33862 33314 33890
rect 32994 33238 33002 33862
rect 33306 33238 33314 33862
rect 32994 33210 33314 33238
rect 33994 33862 34314 33890
rect 33994 33238 34002 33862
rect 34306 33238 34314 33862
rect 33994 33210 34314 33238
rect 9654 33202 34654 33210
rect -57352 32967 -50570 33076
rect -74485 32862 -74165 32890
rect -74485 32238 -74477 32862
rect -74173 32238 -74165 32862
rect -74485 32210 -74165 32238
rect -73485 32862 -73165 32890
rect -73485 32238 -73477 32862
rect -73173 32238 -73165 32862
rect -73485 32210 -73165 32238
rect -72485 32862 -72165 32890
rect -72485 32238 -72477 32862
rect -72173 32238 -72165 32862
rect -72485 32210 -72165 32238
rect -71485 32862 -71165 32890
rect -71485 32238 -71477 32862
rect -71173 32238 -71165 32862
rect -71485 32210 -71165 32238
rect -70485 32862 -70165 32890
rect -70485 32238 -70477 32862
rect -70173 32238 -70165 32862
rect -70485 32210 -70165 32238
rect -69485 32862 -69165 32890
rect -69485 32238 -69477 32862
rect -69173 32238 -69165 32862
rect -69485 32210 -69165 32238
rect -68485 32862 -68165 32890
rect -68485 32238 -68477 32862
rect -68173 32238 -68165 32862
rect -68485 32210 -68165 32238
rect -67485 32862 -67165 32890
rect -67485 32238 -67477 32862
rect -67173 32238 -67165 32862
rect -67485 32210 -67165 32238
rect -66485 32862 -66165 32890
rect -66485 32238 -66477 32862
rect -66173 32238 -66165 32862
rect -66485 32210 -66165 32238
rect -65485 32862 -65165 32890
rect -65485 32238 -65477 32862
rect -65173 32238 -65165 32862
rect -65485 32210 -65165 32238
rect -64485 32862 -64165 32890
rect -64485 32238 -64477 32862
rect -64173 32238 -64165 32862
rect -64485 32210 -64165 32238
rect -63485 32862 -63165 32890
rect -63485 32238 -63477 32862
rect -63173 32238 -63165 32862
rect -63485 32210 -63165 32238
rect -62485 32862 -62165 32890
rect -62485 32238 -62477 32862
rect -62173 32238 -62165 32862
rect -62485 32210 -62165 32238
rect -61485 32862 -61165 32890
rect -61485 32238 -61477 32862
rect -61173 32238 -61165 32862
rect -61485 32210 -61165 32238
rect -60485 32862 -60165 32890
rect -60485 32238 -60477 32862
rect -60173 32238 -60165 32862
rect -60485 32210 -60165 32238
rect -59485 32862 -59165 32890
rect -59485 32238 -59477 32862
rect -59173 32238 -59165 32862
rect -57352 32591 -50955 32967
rect -50579 32591 -50570 32967
rect 9654 32898 9662 33202
rect 9966 32898 10002 33202
rect 10306 32898 10342 33202
rect 10966 32898 11002 33202
rect 11306 32898 11342 33202
rect 11966 32898 12002 33202
rect 12306 32898 12342 33202
rect 12966 32898 13002 33202
rect 13306 32898 13342 33202
rect 13966 32898 14002 33202
rect 14306 32898 14342 33202
rect 14966 32898 15002 33202
rect 15306 32898 15342 33202
rect 15966 32898 16002 33202
rect 16306 32898 16342 33202
rect 16966 32898 17002 33202
rect 17306 32898 17342 33202
rect 17966 32898 18002 33202
rect 18306 32898 18342 33202
rect 18966 32898 19002 33202
rect 19306 32898 19342 33202
rect 19966 32898 20002 33202
rect 20306 32898 20342 33202
rect 20966 32898 21002 33202
rect 21306 32898 21342 33202
rect 21966 32898 22002 33202
rect 22306 32898 22342 33202
rect 22966 32898 23002 33202
rect 23306 32898 23342 33202
rect 23966 32898 24002 33202
rect 24306 32898 24342 33202
rect 24966 32898 25002 33202
rect 25306 32898 25342 33202
rect 25966 32898 26002 33202
rect 26306 32898 26342 33202
rect 26966 32898 27002 33202
rect 27306 32898 27342 33202
rect 27966 32898 28002 33202
rect 28306 32898 28342 33202
rect 28966 32898 29002 33202
rect 29306 32898 29342 33202
rect 29966 32898 30002 33202
rect 30306 32898 30342 33202
rect 30966 32898 31002 33202
rect 31306 32898 31342 33202
rect 31966 32898 32002 33202
rect 32306 32898 32342 33202
rect 32966 32898 33002 33202
rect 33306 32898 33342 33202
rect 33966 32898 34002 33202
rect 34306 32898 34342 33202
rect 34646 32898 34654 33202
rect 9654 32890 34654 32898
rect -57352 32476 -50570 32591
rect 9994 32862 10314 32890
rect -59485 32210 -59165 32238
rect 9994 32238 10002 32862
rect 10306 32238 10314 32862
rect 9994 32210 10314 32238
rect 10994 32862 11314 32890
rect 10994 32238 11002 32862
rect 11306 32238 11314 32862
rect 10994 32210 11314 32238
rect 11994 32862 12314 32890
rect 11994 32238 12002 32862
rect 12306 32238 12314 32862
rect 11994 32210 12314 32238
rect 12994 32862 13314 32890
rect 12994 32238 13002 32862
rect 13306 32238 13314 32862
rect 12994 32210 13314 32238
rect 13994 32862 14314 32890
rect 13994 32238 14002 32862
rect 14306 32238 14314 32862
rect 13994 32210 14314 32238
rect 14994 32862 15314 32890
rect 14994 32238 15002 32862
rect 15306 32238 15314 32862
rect 14994 32210 15314 32238
rect 15994 32862 16314 32890
rect 15994 32238 16002 32862
rect 16306 32238 16314 32862
rect 15994 32210 16314 32238
rect 16994 32862 17314 32890
rect 16994 32238 17002 32862
rect 17306 32238 17314 32862
rect 16994 32210 17314 32238
rect 17994 32862 18314 32890
rect 17994 32238 18002 32862
rect 18306 32238 18314 32862
rect 17994 32210 18314 32238
rect 18994 32862 19314 32890
rect 18994 32238 19002 32862
rect 19306 32238 19314 32862
rect 18994 32210 19314 32238
rect 19994 32862 20314 32890
rect 19994 32238 20002 32862
rect 20306 32238 20314 32862
rect 19994 32210 20314 32238
rect 20994 32862 21314 32890
rect 20994 32238 21002 32862
rect 21306 32238 21314 32862
rect 20994 32210 21314 32238
rect 21994 32862 22314 32890
rect 21994 32238 22002 32862
rect 22306 32238 22314 32862
rect 21994 32210 22314 32238
rect 22994 32862 23314 32890
rect 22994 32238 23002 32862
rect 23306 32238 23314 32862
rect 22994 32210 23314 32238
rect 23994 32862 24314 32890
rect 23994 32238 24002 32862
rect 24306 32238 24314 32862
rect 23994 32210 24314 32238
rect 24994 32862 25314 32890
rect 24994 32238 25002 32862
rect 25306 32238 25314 32862
rect 24994 32210 25314 32238
rect 25994 32862 26314 32890
rect 25994 32238 26002 32862
rect 26306 32238 26314 32862
rect 25994 32210 26314 32238
rect 26994 32862 27314 32890
rect 26994 32238 27002 32862
rect 27306 32238 27314 32862
rect 26994 32210 27314 32238
rect 27994 32862 28314 32890
rect 27994 32238 28002 32862
rect 28306 32238 28314 32862
rect 27994 32210 28314 32238
rect 28994 32862 29314 32890
rect 28994 32238 29002 32862
rect 29306 32238 29314 32862
rect 28994 32210 29314 32238
rect 29994 32862 30314 32890
rect 29994 32238 30002 32862
rect 30306 32238 30314 32862
rect 29994 32210 30314 32238
rect 30994 32862 31314 32890
rect 30994 32238 31002 32862
rect 31306 32238 31314 32862
rect 30994 32210 31314 32238
rect 31994 32862 32314 32890
rect 31994 32238 32002 32862
rect 32306 32238 32314 32862
rect 31994 32210 32314 32238
rect 32994 32862 33314 32890
rect 32994 32238 33002 32862
rect 33306 32238 33314 32862
rect 32994 32210 33314 32238
rect 33994 32862 34314 32890
rect 33994 32238 34002 32862
rect 34306 32238 34314 32862
rect 33994 32210 34314 32238
rect -74825 32202 -58825 32210
rect -74825 31898 -74817 32202
rect -74513 31898 -74477 32202
rect -74173 31898 -74137 32202
rect -73513 31898 -73477 32202
rect -73173 31898 -73137 32202
rect -72513 31898 -72477 32202
rect -72173 31898 -72137 32202
rect -71513 31898 -71477 32202
rect -71173 31898 -71137 32202
rect -70513 31898 -70477 32202
rect -70173 31898 -70137 32202
rect -69513 31898 -69477 32202
rect -69173 31898 -69137 32202
rect -68513 31898 -68477 32202
rect -68173 31898 -68137 32202
rect -67513 31898 -67477 32202
rect -67173 31898 -67137 32202
rect -66513 31898 -66477 32202
rect -66173 31898 -66137 32202
rect -65513 31898 -65477 32202
rect -65173 31898 -65137 32202
rect -64513 31898 -64477 32202
rect -64173 31898 -64137 32202
rect -63513 31898 -63477 32202
rect -63173 31898 -63137 32202
rect -62513 31898 -62477 32202
rect -62173 31898 -62137 32202
rect -61513 31898 -61477 32202
rect -61173 31898 -61137 32202
rect -60513 31898 -60477 32202
rect -60173 31898 -60137 32202
rect -59513 31898 -59477 32202
rect -59173 31898 -59137 32202
rect -58833 31898 -58825 32202
rect -74825 31890 -58825 31898
rect 9654 32202 34654 32210
rect 9654 31898 9662 32202
rect 9966 31898 10002 32202
rect 10306 31898 10342 32202
rect 10966 31898 11002 32202
rect 11306 31898 11342 32202
rect 11966 31898 12002 32202
rect 12306 31898 12342 32202
rect 12966 31898 13002 32202
rect 13306 31898 13342 32202
rect 13966 31898 14002 32202
rect 14306 31898 14342 32202
rect 14966 31898 15002 32202
rect 15306 31898 15342 32202
rect 15966 31898 16002 32202
rect 16306 31898 16342 32202
rect 16966 31898 17002 32202
rect 17306 31898 17342 32202
rect 17966 31898 18002 32202
rect 18306 31898 18342 32202
rect 18966 31898 19002 32202
rect 19306 31898 19342 32202
rect 19966 31898 20002 32202
rect 20306 31898 20342 32202
rect 20966 31898 21002 32202
rect 21306 31898 21342 32202
rect 21966 31898 22002 32202
rect 22306 31898 22342 32202
rect 22966 31898 23002 32202
rect 23306 31898 23342 32202
rect 23966 31898 24002 32202
rect 24306 31898 24342 32202
rect 24966 31898 25002 32202
rect 25306 31898 25342 32202
rect 25966 31898 26002 32202
rect 26306 31898 26342 32202
rect 26966 31898 27002 32202
rect 27306 31898 27342 32202
rect 27966 31898 28002 32202
rect 28306 31898 28342 32202
rect 28966 31898 29002 32202
rect 29306 31898 29342 32202
rect 29966 31898 30002 32202
rect 30306 31898 30342 32202
rect 30966 31898 31002 32202
rect 31306 31898 31342 32202
rect 31966 31898 32002 32202
rect 32306 31898 32342 32202
rect 32966 31898 33002 32202
rect 33306 31898 33342 32202
rect 33966 31898 34002 32202
rect 34306 31898 34342 32202
rect 34646 31898 34654 32202
rect 9654 31890 34654 31898
rect -74485 31862 -74165 31890
rect -74485 31238 -74477 31862
rect -74173 31238 -74165 31862
rect -74485 31210 -74165 31238
rect -73485 31862 -73165 31890
rect -73485 31238 -73477 31862
rect -73173 31238 -73165 31862
rect -73485 31210 -73165 31238
rect -72485 31862 -72165 31890
rect -72485 31238 -72477 31862
rect -72173 31238 -72165 31862
rect -72485 31210 -72165 31238
rect -71485 31862 -71165 31890
rect -71485 31238 -71477 31862
rect -71173 31238 -71165 31862
rect -71485 31210 -71165 31238
rect -70485 31862 -70165 31890
rect -70485 31238 -70477 31862
rect -70173 31238 -70165 31862
rect -70485 31210 -70165 31238
rect -69485 31862 -69165 31890
rect -69485 31238 -69477 31862
rect -69173 31238 -69165 31862
rect -69485 31210 -69165 31238
rect -68485 31862 -68165 31890
rect -68485 31238 -68477 31862
rect -68173 31238 -68165 31862
rect -68485 31210 -68165 31238
rect -67485 31862 -67165 31890
rect -67485 31238 -67477 31862
rect -67173 31238 -67165 31862
rect -67485 31210 -67165 31238
rect -66485 31862 -66165 31890
rect -66485 31238 -66477 31862
rect -66173 31238 -66165 31862
rect -66485 31210 -66165 31238
rect -65485 31862 -65165 31890
rect -65485 31238 -65477 31862
rect -65173 31238 -65165 31862
rect -65485 31210 -65165 31238
rect -64485 31862 -64165 31890
rect -64485 31238 -64477 31862
rect -64173 31238 -64165 31862
rect -64485 31210 -64165 31238
rect -63485 31862 -63165 31890
rect -63485 31238 -63477 31862
rect -63173 31238 -63165 31862
rect -63485 31210 -63165 31238
rect -62485 31862 -62165 31890
rect -62485 31238 -62477 31862
rect -62173 31238 -62165 31862
rect -62485 31210 -62165 31238
rect -61485 31862 -61165 31890
rect -61485 31238 -61477 31862
rect -61173 31238 -61165 31862
rect -61485 31210 -61165 31238
rect -60485 31862 -60165 31890
rect -60485 31238 -60477 31862
rect -60173 31238 -60165 31862
rect -60485 31210 -60165 31238
rect -59485 31862 -59165 31890
rect -59485 31238 -59477 31862
rect -59173 31238 -59165 31862
rect -59485 31210 -59165 31238
rect 9994 31862 10314 31890
rect 9994 31238 10002 31862
rect 10306 31238 10314 31862
rect 9994 31210 10314 31238
rect 10994 31862 11314 31890
rect 10994 31238 11002 31862
rect 11306 31238 11314 31862
rect 10994 31210 11314 31238
rect 11994 31862 12314 31890
rect 11994 31238 12002 31862
rect 12306 31238 12314 31862
rect 11994 31210 12314 31238
rect 12994 31862 13314 31890
rect 12994 31238 13002 31862
rect 13306 31238 13314 31862
rect 12994 31210 13314 31238
rect 13994 31862 14314 31890
rect 13994 31238 14002 31862
rect 14306 31238 14314 31862
rect 13994 31210 14314 31238
rect 14994 31862 15314 31890
rect 14994 31238 15002 31862
rect 15306 31238 15314 31862
rect 14994 31210 15314 31238
rect 15994 31862 16314 31890
rect 15994 31238 16002 31862
rect 16306 31238 16314 31862
rect 15994 31210 16314 31238
rect 16994 31862 17314 31890
rect 16994 31238 17002 31862
rect 17306 31238 17314 31862
rect 16994 31210 17314 31238
rect 17994 31862 18314 31890
rect 17994 31238 18002 31862
rect 18306 31238 18314 31862
rect 17994 31210 18314 31238
rect 18994 31862 19314 31890
rect 18994 31238 19002 31862
rect 19306 31238 19314 31862
rect 18994 31210 19314 31238
rect 19994 31862 20314 31890
rect 19994 31238 20002 31862
rect 20306 31238 20314 31862
rect 19994 31210 20314 31238
rect 20994 31862 21314 31890
rect 20994 31238 21002 31862
rect 21306 31238 21314 31862
rect 20994 31210 21314 31238
rect 21994 31862 22314 31890
rect 21994 31238 22002 31862
rect 22306 31238 22314 31862
rect 21994 31210 22314 31238
rect 22994 31862 23314 31890
rect 22994 31238 23002 31862
rect 23306 31238 23314 31862
rect 22994 31210 23314 31238
rect 23994 31862 24314 31890
rect 23994 31238 24002 31862
rect 24306 31238 24314 31862
rect 23994 31210 24314 31238
rect 24994 31862 25314 31890
rect 24994 31238 25002 31862
rect 25306 31238 25314 31862
rect 24994 31210 25314 31238
rect 25994 31862 26314 31890
rect 25994 31238 26002 31862
rect 26306 31238 26314 31862
rect 25994 31210 26314 31238
rect 26994 31862 27314 31890
rect 26994 31238 27002 31862
rect 27306 31238 27314 31862
rect 26994 31210 27314 31238
rect 27994 31862 28314 31890
rect 27994 31238 28002 31862
rect 28306 31238 28314 31862
rect 27994 31210 28314 31238
rect 28994 31862 29314 31890
rect 28994 31238 29002 31862
rect 29306 31238 29314 31862
rect 28994 31210 29314 31238
rect 29994 31862 30314 31890
rect 29994 31238 30002 31862
rect 30306 31238 30314 31862
rect 29994 31210 30314 31238
rect 30994 31862 31314 31890
rect 30994 31238 31002 31862
rect 31306 31238 31314 31862
rect 30994 31210 31314 31238
rect 31994 31862 32314 31890
rect 31994 31238 32002 31862
rect 32306 31238 32314 31862
rect 31994 31210 32314 31238
rect 32994 31862 33314 31890
rect 32994 31238 33002 31862
rect 33306 31238 33314 31862
rect 32994 31210 33314 31238
rect 33994 31862 34314 31890
rect 33994 31238 34002 31862
rect 34306 31238 34314 31862
rect 33994 31210 34314 31238
rect -74825 31202 -58825 31210
rect -74825 30898 -74817 31202
rect -74513 30898 -74477 31202
rect -74173 30898 -74137 31202
rect -73513 30898 -73477 31202
rect -73173 30898 -73137 31202
rect -72513 30898 -72477 31202
rect -72173 30898 -72137 31202
rect -71513 30898 -71477 31202
rect -71173 30898 -71137 31202
rect -70513 30898 -70477 31202
rect -70173 30898 -70137 31202
rect -69513 30898 -69477 31202
rect -69173 30898 -69137 31202
rect -68513 30898 -68477 31202
rect -68173 30898 -68137 31202
rect -67513 30898 -67477 31202
rect -67173 30898 -67137 31202
rect -66513 30898 -66477 31202
rect -66173 30898 -66137 31202
rect -65513 30898 -65477 31202
rect -65173 30898 -65137 31202
rect -64513 30898 -64477 31202
rect -64173 30898 -64137 31202
rect -63513 30898 -63477 31202
rect -63173 30898 -63137 31202
rect -62513 30898 -62477 31202
rect -62173 30898 -62137 31202
rect -61513 30898 -61477 31202
rect -61173 30898 -61137 31202
rect -60513 30898 -60477 31202
rect -60173 30898 -60137 31202
rect -59513 30898 -59477 31202
rect -59173 30898 -59137 31202
rect -58833 30898 -58825 31202
rect -74825 30890 -58825 30898
rect 9654 31202 34654 31210
rect 9654 30898 9662 31202
rect 9966 30898 10002 31202
rect 10306 30898 10342 31202
rect 10966 30898 11002 31202
rect 11306 30898 11342 31202
rect 11966 30898 12002 31202
rect 12306 30898 12342 31202
rect 12966 30898 13002 31202
rect 13306 30898 13342 31202
rect 13966 30898 14002 31202
rect 14306 30898 14342 31202
rect 14966 30898 15002 31202
rect 15306 30898 15342 31202
rect 15966 30898 16002 31202
rect 16306 30898 16342 31202
rect 16966 30898 17002 31202
rect 17306 30898 17342 31202
rect 17966 30898 18002 31202
rect 18306 30898 18342 31202
rect 18966 30898 19002 31202
rect 19306 30898 19342 31202
rect 19966 30898 20002 31202
rect 20306 30898 20342 31202
rect 20966 30898 21002 31202
rect 21306 30898 21342 31202
rect 21966 30898 22002 31202
rect 22306 30898 22342 31202
rect 22966 30898 23002 31202
rect 23306 30898 23342 31202
rect 23966 30898 24002 31202
rect 24306 30898 24342 31202
rect 24966 30898 25002 31202
rect 25306 30898 25342 31202
rect 25966 30898 26002 31202
rect 26306 30898 26342 31202
rect 26966 30898 27002 31202
rect 27306 30898 27342 31202
rect 27966 30898 28002 31202
rect 28306 30898 28342 31202
rect 28966 30898 29002 31202
rect 29306 30898 29342 31202
rect 29966 30898 30002 31202
rect 30306 30898 30342 31202
rect 30966 30898 31002 31202
rect 31306 30898 31342 31202
rect 31966 30898 32002 31202
rect 32306 30898 32342 31202
rect 32966 30898 33002 31202
rect 33306 30898 33342 31202
rect 33966 30898 34002 31202
rect 34306 30898 34342 31202
rect 34646 30898 34654 31202
rect 9654 30890 34654 30898
rect -74485 30862 -74165 30890
rect -74485 30238 -74477 30862
rect -74173 30238 -74165 30862
rect -74485 30210 -74165 30238
rect -73485 30862 -73165 30890
rect -73485 30238 -73477 30862
rect -73173 30238 -73165 30862
rect -73485 30210 -73165 30238
rect -72485 30862 -72165 30890
rect -72485 30238 -72477 30862
rect -72173 30238 -72165 30862
rect -72485 30210 -72165 30238
rect -71485 30862 -71165 30890
rect -71485 30238 -71477 30862
rect -71173 30238 -71165 30862
rect -71485 30210 -71165 30238
rect -70485 30862 -70165 30890
rect -70485 30238 -70477 30862
rect -70173 30238 -70165 30862
rect -70485 30210 -70165 30238
rect -69485 30862 -69165 30890
rect -69485 30238 -69477 30862
rect -69173 30238 -69165 30862
rect -69485 30210 -69165 30238
rect -68485 30862 -68165 30890
rect -68485 30238 -68477 30862
rect -68173 30238 -68165 30862
rect -68485 30210 -68165 30238
rect -67485 30862 -67165 30890
rect -67485 30238 -67477 30862
rect -67173 30238 -67165 30862
rect -67485 30210 -67165 30238
rect -66485 30862 -66165 30890
rect -66485 30238 -66477 30862
rect -66173 30238 -66165 30862
rect -66485 30210 -66165 30238
rect -65485 30862 -65165 30890
rect -65485 30238 -65477 30862
rect -65173 30238 -65165 30862
rect -65485 30210 -65165 30238
rect -64485 30862 -64165 30890
rect -64485 30238 -64477 30862
rect -64173 30238 -64165 30862
rect -64485 30210 -64165 30238
rect -63485 30862 -63165 30890
rect -63485 30238 -63477 30862
rect -63173 30238 -63165 30862
rect -63485 30210 -63165 30238
rect -62485 30862 -62165 30890
rect -62485 30238 -62477 30862
rect -62173 30238 -62165 30862
rect -62485 30210 -62165 30238
rect -61485 30862 -61165 30890
rect -61485 30238 -61477 30862
rect -61173 30238 -61165 30862
rect -61485 30210 -61165 30238
rect -60485 30862 -60165 30890
rect -60485 30238 -60477 30862
rect -60173 30238 -60165 30862
rect -60485 30210 -60165 30238
rect -59485 30862 -59165 30890
rect -59485 30238 -59477 30862
rect -59173 30238 -59165 30862
rect -59485 30210 -59165 30238
rect 9994 30862 10314 30890
rect 9994 30238 10002 30862
rect 10306 30238 10314 30862
rect 9994 30210 10314 30238
rect 10994 30862 11314 30890
rect 10994 30238 11002 30862
rect 11306 30238 11314 30862
rect 10994 30210 11314 30238
rect 11994 30862 12314 30890
rect 11994 30238 12002 30862
rect 12306 30238 12314 30862
rect 11994 30210 12314 30238
rect 12994 30862 13314 30890
rect 12994 30238 13002 30862
rect 13306 30238 13314 30862
rect 12994 30210 13314 30238
rect 13994 30862 14314 30890
rect 13994 30238 14002 30862
rect 14306 30238 14314 30862
rect 13994 30210 14314 30238
rect 14994 30862 15314 30890
rect 14994 30238 15002 30862
rect 15306 30238 15314 30862
rect 14994 30210 15314 30238
rect 15994 30862 16314 30890
rect 15994 30238 16002 30862
rect 16306 30238 16314 30862
rect 15994 30210 16314 30238
rect 16994 30862 17314 30890
rect 16994 30238 17002 30862
rect 17306 30238 17314 30862
rect 16994 30210 17314 30238
rect 17994 30862 18314 30890
rect 17994 30238 18002 30862
rect 18306 30238 18314 30862
rect 17994 30210 18314 30238
rect 18994 30862 19314 30890
rect 18994 30238 19002 30862
rect 19306 30238 19314 30862
rect 18994 30210 19314 30238
rect 19994 30862 20314 30890
rect 19994 30238 20002 30862
rect 20306 30238 20314 30862
rect 19994 30210 20314 30238
rect 20994 30862 21314 30890
rect 20994 30238 21002 30862
rect 21306 30238 21314 30862
rect 20994 30210 21314 30238
rect 21994 30862 22314 30890
rect 21994 30238 22002 30862
rect 22306 30238 22314 30862
rect 21994 30210 22314 30238
rect 22994 30862 23314 30890
rect 22994 30238 23002 30862
rect 23306 30238 23314 30862
rect 22994 30210 23314 30238
rect 23994 30862 24314 30890
rect 23994 30238 24002 30862
rect 24306 30238 24314 30862
rect 23994 30210 24314 30238
rect 24994 30862 25314 30890
rect 24994 30238 25002 30862
rect 25306 30238 25314 30862
rect 24994 30210 25314 30238
rect 25994 30862 26314 30890
rect 25994 30238 26002 30862
rect 26306 30238 26314 30862
rect 25994 30210 26314 30238
rect 26994 30862 27314 30890
rect 26994 30238 27002 30862
rect 27306 30238 27314 30862
rect 26994 30210 27314 30238
rect 27994 30862 28314 30890
rect 27994 30238 28002 30862
rect 28306 30238 28314 30862
rect 27994 30210 28314 30238
rect 28994 30862 29314 30890
rect 28994 30238 29002 30862
rect 29306 30238 29314 30862
rect 28994 30210 29314 30238
rect 29994 30862 30314 30890
rect 29994 30238 30002 30862
rect 30306 30238 30314 30862
rect 29994 30210 30314 30238
rect 30994 30862 31314 30890
rect 30994 30238 31002 30862
rect 31306 30238 31314 30862
rect 30994 30210 31314 30238
rect 31994 30862 32314 30890
rect 31994 30238 32002 30862
rect 32306 30238 32314 30862
rect 31994 30210 32314 30238
rect 32994 30862 33314 30890
rect 32994 30238 33002 30862
rect 33306 30238 33314 30862
rect 32994 30210 33314 30238
rect 33994 30862 34314 30890
rect 33994 30238 34002 30862
rect 34306 30238 34314 30862
rect 33994 30210 34314 30238
rect -74825 30202 -58825 30210
rect -74825 29898 -74817 30202
rect -74513 29898 -74477 30202
rect -74173 29898 -74137 30202
rect -73513 29898 -73477 30202
rect -73173 29898 -73137 30202
rect -72513 29898 -72477 30202
rect -72173 29898 -72137 30202
rect -71513 29898 -71477 30202
rect -71173 29898 -71137 30202
rect -70513 29898 -70477 30202
rect -70173 29898 -70137 30202
rect -69513 29898 -69477 30202
rect -69173 29898 -69137 30202
rect -68513 29898 -68477 30202
rect -68173 29898 -68137 30202
rect -67513 29898 -67477 30202
rect -67173 29898 -67137 30202
rect -66513 29898 -66477 30202
rect -66173 29898 -66137 30202
rect -65513 29898 -65477 30202
rect -65173 29898 -65137 30202
rect -64513 29898 -64477 30202
rect -64173 29898 -64137 30202
rect -63513 29898 -63477 30202
rect -63173 29898 -63137 30202
rect -62513 29898 -62477 30202
rect -62173 29898 -62137 30202
rect -61513 29898 -61477 30202
rect -61173 29898 -61137 30202
rect -60513 29898 -60477 30202
rect -60173 29898 -60137 30202
rect -59513 29898 -59477 30202
rect -59173 29898 -59137 30202
rect -58833 29898 -58825 30202
rect -74825 29890 -58825 29898
rect 9654 30202 34654 30210
rect 9654 29898 9662 30202
rect 9966 29898 10002 30202
rect 10306 29898 10342 30202
rect 10966 29898 11002 30202
rect 11306 29898 11342 30202
rect 11966 29898 12002 30202
rect 12306 29898 12342 30202
rect 12966 29898 13002 30202
rect 13306 29898 13342 30202
rect 13966 29898 14002 30202
rect 14306 29898 14342 30202
rect 14966 29898 15002 30202
rect 15306 29898 15342 30202
rect 15966 29898 16002 30202
rect 16306 29898 16342 30202
rect 16966 29898 17002 30202
rect 17306 29898 17342 30202
rect 17966 29898 18002 30202
rect 18306 29898 18342 30202
rect 18966 29898 19002 30202
rect 19306 29898 19342 30202
rect 19966 29898 20002 30202
rect 20306 29898 20342 30202
rect 20966 29898 21002 30202
rect 21306 29898 21342 30202
rect 21966 29898 22002 30202
rect 22306 29898 22342 30202
rect 22966 29898 23002 30202
rect 23306 29898 23342 30202
rect 23966 29898 24002 30202
rect 24306 29898 24342 30202
rect 24966 29898 25002 30202
rect 25306 29898 25342 30202
rect 25966 29898 26002 30202
rect 26306 29898 26342 30202
rect 26966 29898 27002 30202
rect 27306 29898 27342 30202
rect 27966 29898 28002 30202
rect 28306 29898 28342 30202
rect 28966 29898 29002 30202
rect 29306 29898 29342 30202
rect 29966 29898 30002 30202
rect 30306 29898 30342 30202
rect 30966 29898 31002 30202
rect 31306 29898 31342 30202
rect 31966 29898 32002 30202
rect 32306 29898 32342 30202
rect 32966 29898 33002 30202
rect 33306 29898 33342 30202
rect 33966 29898 34002 30202
rect 34306 29898 34342 30202
rect 34646 29898 34654 30202
rect 9654 29890 34654 29898
rect -74485 29862 -74165 29890
rect -74485 29238 -74477 29862
rect -74173 29238 -74165 29862
rect -74485 29210 -74165 29238
rect -73485 29862 -73165 29890
rect -73485 29238 -73477 29862
rect -73173 29238 -73165 29862
rect -73485 29210 -73165 29238
rect -72485 29862 -72165 29890
rect -72485 29238 -72477 29862
rect -72173 29238 -72165 29862
rect -72485 29210 -72165 29238
rect -71485 29862 -71165 29890
rect -71485 29238 -71477 29862
rect -71173 29238 -71165 29862
rect -71485 29210 -71165 29238
rect -70485 29862 -70165 29890
rect -70485 29238 -70477 29862
rect -70173 29238 -70165 29862
rect -70485 29210 -70165 29238
rect -69485 29862 -69165 29890
rect -69485 29238 -69477 29862
rect -69173 29238 -69165 29862
rect -69485 29210 -69165 29238
rect -68485 29862 -68165 29890
rect -68485 29238 -68477 29862
rect -68173 29238 -68165 29862
rect -68485 29210 -68165 29238
rect -67485 29862 -67165 29890
rect -67485 29238 -67477 29862
rect -67173 29238 -67165 29862
rect -67485 29210 -67165 29238
rect -66485 29862 -66165 29890
rect -66485 29238 -66477 29862
rect -66173 29238 -66165 29862
rect -66485 29210 -66165 29238
rect -65485 29862 -65165 29890
rect -65485 29238 -65477 29862
rect -65173 29238 -65165 29862
rect -65485 29210 -65165 29238
rect -64485 29862 -64165 29890
rect -64485 29238 -64477 29862
rect -64173 29238 -64165 29862
rect -64485 29210 -64165 29238
rect -63485 29862 -63165 29890
rect -63485 29238 -63477 29862
rect -63173 29238 -63165 29862
rect -63485 29210 -63165 29238
rect -62485 29862 -62165 29890
rect -62485 29238 -62477 29862
rect -62173 29238 -62165 29862
rect -62485 29210 -62165 29238
rect -61485 29862 -61165 29890
rect -61485 29238 -61477 29862
rect -61173 29238 -61165 29862
rect -61485 29210 -61165 29238
rect -60485 29862 -60165 29890
rect -60485 29238 -60477 29862
rect -60173 29238 -60165 29862
rect -60485 29210 -60165 29238
rect -59485 29862 -59165 29890
rect -59485 29238 -59477 29862
rect -59173 29238 -59165 29862
rect -59485 29210 -59165 29238
rect 9994 29862 10314 29890
rect 9994 29238 10002 29862
rect 10306 29238 10314 29862
rect 9994 29210 10314 29238
rect 10994 29862 11314 29890
rect 10994 29238 11002 29862
rect 11306 29238 11314 29862
rect 10994 29210 11314 29238
rect 11994 29862 12314 29890
rect 11994 29238 12002 29862
rect 12306 29238 12314 29862
rect 11994 29210 12314 29238
rect 12994 29862 13314 29890
rect 12994 29238 13002 29862
rect 13306 29238 13314 29862
rect 12994 29210 13314 29238
rect 13994 29862 14314 29890
rect 13994 29238 14002 29862
rect 14306 29238 14314 29862
rect 13994 29210 14314 29238
rect 14994 29862 15314 29890
rect 14994 29238 15002 29862
rect 15306 29238 15314 29862
rect 14994 29210 15314 29238
rect 15994 29862 16314 29890
rect 15994 29238 16002 29862
rect 16306 29238 16314 29862
rect 15994 29210 16314 29238
rect 16994 29862 17314 29890
rect 16994 29238 17002 29862
rect 17306 29238 17314 29862
rect 16994 29210 17314 29238
rect 17994 29862 18314 29890
rect 17994 29238 18002 29862
rect 18306 29238 18314 29862
rect 17994 29210 18314 29238
rect 18994 29862 19314 29890
rect 18994 29238 19002 29862
rect 19306 29238 19314 29862
rect 18994 29210 19314 29238
rect 19994 29862 20314 29890
rect 19994 29238 20002 29862
rect 20306 29238 20314 29862
rect 19994 29210 20314 29238
rect 20994 29862 21314 29890
rect 20994 29238 21002 29862
rect 21306 29238 21314 29862
rect 20994 29210 21314 29238
rect 21994 29862 22314 29890
rect 21994 29238 22002 29862
rect 22306 29238 22314 29862
rect 21994 29210 22314 29238
rect 22994 29862 23314 29890
rect 22994 29238 23002 29862
rect 23306 29238 23314 29862
rect 22994 29210 23314 29238
rect 23994 29862 24314 29890
rect 23994 29238 24002 29862
rect 24306 29238 24314 29862
rect 23994 29210 24314 29238
rect 24994 29862 25314 29890
rect 24994 29238 25002 29862
rect 25306 29238 25314 29862
rect 24994 29210 25314 29238
rect 25994 29862 26314 29890
rect 25994 29238 26002 29862
rect 26306 29238 26314 29862
rect 25994 29210 26314 29238
rect 26994 29862 27314 29890
rect 26994 29238 27002 29862
rect 27306 29238 27314 29862
rect 26994 29210 27314 29238
rect 27994 29862 28314 29890
rect 27994 29238 28002 29862
rect 28306 29238 28314 29862
rect 27994 29210 28314 29238
rect 28994 29862 29314 29890
rect 28994 29238 29002 29862
rect 29306 29238 29314 29862
rect 28994 29210 29314 29238
rect 29994 29862 30314 29890
rect 29994 29238 30002 29862
rect 30306 29238 30314 29862
rect 29994 29210 30314 29238
rect 30994 29862 31314 29890
rect 30994 29238 31002 29862
rect 31306 29238 31314 29862
rect 30994 29210 31314 29238
rect 31994 29862 32314 29890
rect 31994 29238 32002 29862
rect 32306 29238 32314 29862
rect 31994 29210 32314 29238
rect 32994 29862 33314 29890
rect 32994 29238 33002 29862
rect 33306 29238 33314 29862
rect 32994 29210 33314 29238
rect 33994 29862 34314 29890
rect 33994 29238 34002 29862
rect 34306 29238 34314 29862
rect 33994 29210 34314 29238
rect -74825 29202 -58825 29210
rect -74825 28898 -74817 29202
rect -74513 28898 -74477 29202
rect -74173 28898 -74137 29202
rect -73513 28898 -73477 29202
rect -73173 28898 -73137 29202
rect -72513 28898 -72477 29202
rect -72173 28898 -72137 29202
rect -71513 28898 -71477 29202
rect -71173 28898 -71137 29202
rect -70513 28898 -70477 29202
rect -70173 28898 -70137 29202
rect -69513 28898 -69477 29202
rect -69173 28898 -69137 29202
rect -68513 28898 -68477 29202
rect -68173 28898 -68137 29202
rect -67513 28898 -67477 29202
rect -67173 28898 -67137 29202
rect -66513 28898 -66477 29202
rect -66173 28898 -66137 29202
rect -65513 28898 -65477 29202
rect -65173 28898 -65137 29202
rect -64513 28898 -64477 29202
rect -64173 28898 -64137 29202
rect -63513 28898 -63477 29202
rect -63173 28898 -63137 29202
rect -62513 28898 -62477 29202
rect -62173 28898 -62137 29202
rect -61513 28898 -61477 29202
rect -61173 28898 -61137 29202
rect -60513 28898 -60477 29202
rect -60173 28898 -60137 29202
rect -59513 28898 -59477 29202
rect -59173 28898 -59137 29202
rect -58833 28898 -58825 29202
rect -74825 28890 -58825 28898
rect 9654 29202 34654 29210
rect 9654 28898 9662 29202
rect 9966 28898 10002 29202
rect 10306 28898 10342 29202
rect 10966 28898 11002 29202
rect 11306 28898 11342 29202
rect 11966 28898 12002 29202
rect 12306 28898 12342 29202
rect 12966 28898 13002 29202
rect 13306 28898 13342 29202
rect 13966 28898 14002 29202
rect 14306 28898 14342 29202
rect 14966 28898 15002 29202
rect 15306 28898 15342 29202
rect 15966 28898 16002 29202
rect 16306 28898 16342 29202
rect 16966 28898 17002 29202
rect 17306 28898 17342 29202
rect 17966 28898 18002 29202
rect 18306 28898 18342 29202
rect 18966 28898 19002 29202
rect 19306 28898 19342 29202
rect 19966 28898 20002 29202
rect 20306 28898 20342 29202
rect 20966 28898 21002 29202
rect 21306 28898 21342 29202
rect 21966 28898 22002 29202
rect 22306 28898 22342 29202
rect 22966 28898 23002 29202
rect 23306 28898 23342 29202
rect 23966 28898 24002 29202
rect 24306 28898 24342 29202
rect 24966 28898 25002 29202
rect 25306 28898 25342 29202
rect 25966 28898 26002 29202
rect 26306 28898 26342 29202
rect 26966 28898 27002 29202
rect 27306 28898 27342 29202
rect 27966 28898 28002 29202
rect 28306 28898 28342 29202
rect 28966 28898 29002 29202
rect 29306 28898 29342 29202
rect 29966 28898 30002 29202
rect 30306 28898 30342 29202
rect 30966 28898 31002 29202
rect 31306 28898 31342 29202
rect 31966 28898 32002 29202
rect 32306 28898 32342 29202
rect 32966 28898 33002 29202
rect 33306 28898 33342 29202
rect 33966 28898 34002 29202
rect 34306 28898 34342 29202
rect 34646 28898 34654 29202
rect 9654 28890 34654 28898
rect -74485 28862 -74165 28890
rect -74485 28558 -74477 28862
rect -74173 28558 -74165 28862
rect -74485 28550 -74165 28558
rect -73485 28862 -73165 28890
rect -73485 28558 -73477 28862
rect -73173 28558 -73165 28862
rect -73485 28550 -73165 28558
rect -72485 28862 -72165 28890
rect -72485 28558 -72477 28862
rect -72173 28558 -72165 28862
rect -72485 28550 -72165 28558
rect -71485 28862 -71165 28890
rect -71485 28558 -71477 28862
rect -71173 28558 -71165 28862
rect -71485 28550 -71165 28558
rect -70485 28862 -70165 28890
rect -70485 28558 -70477 28862
rect -70173 28558 -70165 28862
rect -70485 28550 -70165 28558
rect -69485 28862 -69165 28890
rect -69485 28558 -69477 28862
rect -69173 28558 -69165 28862
rect -69485 28550 -69165 28558
rect -68485 28862 -68165 28890
rect -68485 28558 -68477 28862
rect -68173 28558 -68165 28862
rect -68485 28550 -68165 28558
rect -67485 28862 -67165 28890
rect -67485 28558 -67477 28862
rect -67173 28558 -67165 28862
rect -67485 28550 -67165 28558
rect -66485 28862 -66165 28890
rect -66485 28558 -66477 28862
rect -66173 28558 -66165 28862
rect -66485 28550 -66165 28558
rect -65485 28862 -65165 28890
rect -65485 28558 -65477 28862
rect -65173 28558 -65165 28862
rect -65485 28550 -65165 28558
rect -64485 28862 -64165 28890
rect -64485 28558 -64477 28862
rect -64173 28558 -64165 28862
rect -64485 28550 -64165 28558
rect -63485 28862 -63165 28890
rect -63485 28558 -63477 28862
rect -63173 28558 -63165 28862
rect -63485 28550 -63165 28558
rect -62485 28862 -62165 28890
rect -62485 28558 -62477 28862
rect -62173 28558 -62165 28862
rect -62485 28550 -62165 28558
rect -61485 28862 -61165 28890
rect -61485 28558 -61477 28862
rect -61173 28558 -61165 28862
rect -61485 28550 -61165 28558
rect -60485 28862 -60165 28890
rect -60485 28558 -60477 28862
rect -60173 28558 -60165 28862
rect -60485 28550 -60165 28558
rect -59485 28862 -59165 28890
rect -59485 28558 -59477 28862
rect -59173 28558 -59165 28862
rect -59485 28550 -59165 28558
rect 9994 28862 10314 28890
rect 9994 28558 10002 28862
rect 10306 28558 10314 28862
rect 9994 28550 10314 28558
rect 10994 28862 11314 28890
rect 10994 28558 11002 28862
rect 11306 28558 11314 28862
rect 10994 28550 11314 28558
rect 11994 28862 12314 28890
rect 11994 28558 12002 28862
rect 12306 28558 12314 28862
rect 11994 28550 12314 28558
rect 12994 28862 13314 28890
rect 12994 28558 13002 28862
rect 13306 28558 13314 28862
rect 12994 28550 13314 28558
rect 13994 28862 14314 28890
rect 13994 28558 14002 28862
rect 14306 28558 14314 28862
rect 13994 28550 14314 28558
rect 14994 28862 15314 28890
rect 14994 28558 15002 28862
rect 15306 28558 15314 28862
rect 14994 28550 15314 28558
rect 15994 28862 16314 28890
rect 15994 28558 16002 28862
rect 16306 28558 16314 28862
rect 15994 28550 16314 28558
rect 16994 28862 17314 28890
rect 16994 28558 17002 28862
rect 17306 28558 17314 28862
rect 16994 28550 17314 28558
rect 17994 28862 18314 28890
rect 17994 28558 18002 28862
rect 18306 28558 18314 28862
rect 17994 28550 18314 28558
rect 18994 28862 19314 28890
rect 18994 28558 19002 28862
rect 19306 28558 19314 28862
rect 18994 28550 19314 28558
rect 19994 28862 20314 28890
rect 19994 28558 20002 28862
rect 20306 28558 20314 28862
rect 19994 28550 20314 28558
rect 20994 28862 21314 28890
rect 20994 28558 21002 28862
rect 21306 28558 21314 28862
rect 20994 28550 21314 28558
rect 21994 28862 22314 28890
rect 21994 28558 22002 28862
rect 22306 28558 22314 28862
rect 21994 28550 22314 28558
rect 22994 28862 23314 28890
rect 22994 28558 23002 28862
rect 23306 28558 23314 28862
rect 22994 28550 23314 28558
rect 23994 28862 24314 28890
rect 23994 28558 24002 28862
rect 24306 28558 24314 28862
rect 23994 28550 24314 28558
rect 24994 28862 25314 28890
rect 24994 28558 25002 28862
rect 25306 28558 25314 28862
rect 24994 28550 25314 28558
rect 25994 28862 26314 28890
rect 25994 28558 26002 28862
rect 26306 28558 26314 28862
rect 25994 28550 26314 28558
rect 26994 28862 27314 28890
rect 26994 28558 27002 28862
rect 27306 28558 27314 28862
rect 26994 28550 27314 28558
rect 27994 28862 28314 28890
rect 27994 28558 28002 28862
rect 28306 28558 28314 28862
rect 27994 28550 28314 28558
rect 28994 28862 29314 28890
rect 28994 28558 29002 28862
rect 29306 28558 29314 28862
rect 28994 28550 29314 28558
rect 29994 28862 30314 28890
rect 29994 28558 30002 28862
rect 30306 28558 30314 28862
rect 29994 28550 30314 28558
rect 30994 28862 31314 28890
rect 30994 28558 31002 28862
rect 31306 28558 31314 28862
rect 30994 28550 31314 28558
rect 31994 28862 32314 28890
rect 31994 28558 32002 28862
rect 32306 28558 32314 28862
rect 31994 28550 32314 28558
rect 32994 28862 33314 28890
rect 32994 28558 33002 28862
rect 33306 28558 33314 28862
rect 32994 28550 33314 28558
rect 33994 28862 34314 28890
rect 33994 28558 34002 28862
rect 34306 28558 34314 28862
rect 33994 28550 34314 28558
rect -72825 25947 -60825 26000
rect -72825 16043 -72782 25947
rect -60878 16043 -60825 25947
rect -72825 16000 -60825 16043
rect 20275 25952 32275 26000
rect 20275 16048 20318 25952
rect 32222 16048 32275 25952
rect 20275 16000 32275 16048
rect -21216 15122 -19300 15128
rect -21216 13858 -21210 15122
rect -19306 13858 -19300 15122
rect -21216 13852 -19300 13858
rect -42440 13802 -40660 13850
rect -42440 7898 -42382 13802
rect -40718 7898 -40660 13802
rect -42440 7850 -40660 7898
rect 110 13802 1890 13850
rect 110 7898 168 13802
rect 1832 7898 1890 13802
rect 110 7850 1890 7898
rect -42440 2312 -40660 2350
rect -42440 -2312 -42382 2312
rect -40718 -2312 -40660 2312
rect -42440 -2350 -40660 -2312
rect 110 2312 1890 2350
rect 110 -2312 168 2312
rect 1832 -2312 1890 2312
rect 110 -2350 1890 -2312
rect -42440 -7898 -40660 -7850
rect -42440 -13802 -42382 -7898
rect -40718 -13802 -40660 -7898
rect -42440 -13850 -40660 -13802
rect 110 -7898 1890 -7850
rect 110 -13802 168 -7898
rect 1832 -13802 1890 -7898
rect 110 -13850 1890 -13802
rect -72825 -16048 -60825 -16000
rect -72825 -25952 -72782 -16048
rect -60878 -25952 -60825 -16048
rect -72825 -26000 -60825 -25952
rect 20275 -16048 32275 -16000
rect 20275 -25952 20318 -16048
rect 32222 -25952 32275 -16048
rect 20275 -26000 32275 -25952
rect -74485 -28558 -74165 -28550
rect -74485 -28862 -74477 -28558
rect -74173 -28862 -74165 -28558
rect -74485 -28890 -74165 -28862
rect -73485 -28558 -73165 -28550
rect -73485 -28862 -73477 -28558
rect -73173 -28862 -73165 -28558
rect -73485 -28890 -73165 -28862
rect -72485 -28558 -72165 -28550
rect -72485 -28862 -72477 -28558
rect -72173 -28862 -72165 -28558
rect -72485 -28890 -72165 -28862
rect -71485 -28558 -71165 -28550
rect -71485 -28862 -71477 -28558
rect -71173 -28862 -71165 -28558
rect -71485 -28890 -71165 -28862
rect -70485 -28558 -70165 -28550
rect -70485 -28862 -70477 -28558
rect -70173 -28862 -70165 -28558
rect -70485 -28890 -70165 -28862
rect -69485 -28558 -69165 -28550
rect -69485 -28862 -69477 -28558
rect -69173 -28862 -69165 -28558
rect -69485 -28890 -69165 -28862
rect -68485 -28558 -68165 -28550
rect -68485 -28862 -68477 -28558
rect -68173 -28862 -68165 -28558
rect -68485 -28890 -68165 -28862
rect -67485 -28558 -67165 -28550
rect -67485 -28862 -67477 -28558
rect -67173 -28862 -67165 -28558
rect -67485 -28890 -67165 -28862
rect -66485 -28558 -66165 -28550
rect -66485 -28862 -66477 -28558
rect -66173 -28862 -66165 -28558
rect -66485 -28890 -66165 -28862
rect -65485 -28558 -65165 -28550
rect -65485 -28862 -65477 -28558
rect -65173 -28862 -65165 -28558
rect -65485 -28890 -65165 -28862
rect -64485 -28558 -64165 -28550
rect -64485 -28862 -64477 -28558
rect -64173 -28862 -64165 -28558
rect -64485 -28890 -64165 -28862
rect -63485 -28558 -63165 -28550
rect -63485 -28862 -63477 -28558
rect -63173 -28862 -63165 -28558
rect -63485 -28890 -63165 -28862
rect -62485 -28558 -62165 -28550
rect -62485 -28862 -62477 -28558
rect -62173 -28862 -62165 -28558
rect -62485 -28890 -62165 -28862
rect -61485 -28558 -61165 -28550
rect -61485 -28862 -61477 -28558
rect -61173 -28862 -61165 -28558
rect -61485 -28890 -61165 -28862
rect -60485 -28558 -60165 -28550
rect -60485 -28862 -60477 -28558
rect -60173 -28862 -60165 -28558
rect -60485 -28890 -60165 -28862
rect -59485 -28558 -59165 -28550
rect -59485 -28862 -59477 -28558
rect -59173 -28862 -59165 -28558
rect -59485 -28890 -59165 -28862
rect -58485 -28558 -58165 -28550
rect -58485 -28862 -58477 -28558
rect -58173 -28862 -58165 -28558
rect -58485 -28890 -58165 -28862
rect -57485 -28558 -57165 -28550
rect -57485 -28862 -57477 -28558
rect -57173 -28862 -57165 -28558
rect -57485 -28890 -57165 -28862
rect -56485 -28558 -56165 -28550
rect -56485 -28862 -56477 -28558
rect -56173 -28862 -56165 -28558
rect -56485 -28890 -56165 -28862
rect -55485 -28558 -55165 -28550
rect -55485 -28862 -55477 -28558
rect -55173 -28862 -55165 -28558
rect -55485 -28890 -55165 -28862
rect -54485 -28558 -54165 -28550
rect -54485 -28862 -54477 -28558
rect -54173 -28862 -54165 -28558
rect -54485 -28890 -54165 -28862
rect -53485 -28558 -53165 -28550
rect -53485 -28862 -53477 -28558
rect -53173 -28862 -53165 -28558
rect -53485 -28890 -53165 -28862
rect -52485 -28558 -52165 -28550
rect -52485 -28862 -52477 -28558
rect -52173 -28862 -52165 -28558
rect -52485 -28890 -52165 -28862
rect -51485 -28558 -51165 -28550
rect -51485 -28862 -51477 -28558
rect -51173 -28862 -51165 -28558
rect -51485 -28890 -51165 -28862
rect -50485 -28558 -50165 -28550
rect -50485 -28862 -50477 -28558
rect -50173 -28862 -50165 -28558
rect -50485 -28890 -50165 -28862
rect -49485 -28558 -49165 -28550
rect -49485 -28862 -49477 -28558
rect -49173 -28862 -49165 -28558
rect -49485 -28890 -49165 -28862
rect 8615 -28558 8935 -28550
rect 8615 -28862 8623 -28558
rect 8927 -28862 8935 -28558
rect 8615 -28890 8935 -28862
rect 9615 -28558 9935 -28550
rect 9615 -28862 9623 -28558
rect 9927 -28862 9935 -28558
rect 9615 -28890 9935 -28862
rect 10615 -28558 10935 -28550
rect 10615 -28862 10623 -28558
rect 10927 -28862 10935 -28558
rect 10615 -28890 10935 -28862
rect 11615 -28558 11935 -28550
rect 11615 -28862 11623 -28558
rect 11927 -28862 11935 -28558
rect 11615 -28890 11935 -28862
rect 12615 -28558 12935 -28550
rect 12615 -28862 12623 -28558
rect 12927 -28862 12935 -28558
rect 12615 -28890 12935 -28862
rect 13615 -28558 13935 -28550
rect 13615 -28862 13623 -28558
rect 13927 -28862 13935 -28558
rect 13615 -28890 13935 -28862
rect 14615 -28558 14935 -28550
rect 14615 -28862 14623 -28558
rect 14927 -28862 14935 -28558
rect 14615 -28890 14935 -28862
rect 15615 -28558 15935 -28550
rect 15615 -28862 15623 -28558
rect 15927 -28862 15935 -28558
rect 15615 -28890 15935 -28862
rect 16615 -28558 16935 -28550
rect 16615 -28862 16623 -28558
rect 16927 -28862 16935 -28558
rect 16615 -28890 16935 -28862
rect 17615 -28558 17935 -28550
rect 17615 -28862 17623 -28558
rect 17927 -28862 17935 -28558
rect 17615 -28890 17935 -28862
rect 18615 -28558 18935 -28550
rect 18615 -28862 18623 -28558
rect 18927 -28862 18935 -28558
rect 18615 -28890 18935 -28862
rect 19615 -28558 19935 -28550
rect 19615 -28862 19623 -28558
rect 19927 -28862 19935 -28558
rect 19615 -28890 19935 -28862
rect 20615 -28558 20935 -28550
rect 20615 -28862 20623 -28558
rect 20927 -28862 20935 -28558
rect 20615 -28890 20935 -28862
rect 21615 -28558 21935 -28550
rect 21615 -28862 21623 -28558
rect 21927 -28862 21935 -28558
rect 21615 -28890 21935 -28862
rect 22615 -28558 22935 -28550
rect 22615 -28862 22623 -28558
rect 22927 -28862 22935 -28558
rect 22615 -28890 22935 -28862
rect 23615 -28558 23935 -28550
rect 23615 -28862 23623 -28558
rect 23927 -28862 23935 -28558
rect 23615 -28890 23935 -28862
rect 24615 -28558 24935 -28550
rect 24615 -28862 24623 -28558
rect 24927 -28862 24935 -28558
rect 24615 -28890 24935 -28862
rect 25615 -28558 25935 -28550
rect 25615 -28862 25623 -28558
rect 25927 -28862 25935 -28558
rect 25615 -28890 25935 -28862
rect 26615 -28558 26935 -28550
rect 26615 -28862 26623 -28558
rect 26927 -28862 26935 -28558
rect 26615 -28890 26935 -28862
rect 27615 -28558 27935 -28550
rect 27615 -28862 27623 -28558
rect 27927 -28862 27935 -28558
rect 27615 -28890 27935 -28862
rect 28615 -28558 28935 -28550
rect 28615 -28862 28623 -28558
rect 28927 -28862 28935 -28558
rect 28615 -28890 28935 -28862
rect 29615 -28558 29935 -28550
rect 29615 -28862 29623 -28558
rect 29927 -28862 29935 -28558
rect 29615 -28890 29935 -28862
rect 30615 -28558 30935 -28550
rect 30615 -28862 30623 -28558
rect 30927 -28862 30935 -28558
rect 30615 -28890 30935 -28862
rect 31615 -28558 31935 -28550
rect 31615 -28862 31623 -28558
rect 31927 -28862 31935 -28558
rect 31615 -28890 31935 -28862
rect 32615 -28558 32935 -28550
rect 32615 -28862 32623 -28558
rect 32927 -28862 32935 -28558
rect 32615 -28890 32935 -28862
rect 33615 -28558 33935 -28550
rect 33615 -28862 33623 -28558
rect 33927 -28862 33935 -28558
rect 33615 -28890 33935 -28862
rect -74825 -28898 -48825 -28890
rect -74825 -29202 -74817 -28898
rect -74513 -29202 -74477 -28898
rect -74173 -29202 -74137 -28898
rect -73513 -29202 -73477 -28898
rect -73173 -29202 -73137 -28898
rect -72513 -29202 -72477 -28898
rect -72173 -29202 -72137 -28898
rect -71513 -29202 -71477 -28898
rect -71173 -29202 -71137 -28898
rect -70513 -29202 -70477 -28898
rect -70173 -29202 -70137 -28898
rect -69513 -29202 -69477 -28898
rect -69173 -29202 -69137 -28898
rect -68513 -29202 -68477 -28898
rect -68173 -29202 -68137 -28898
rect -67513 -29202 -67477 -28898
rect -67173 -29202 -67137 -28898
rect -66513 -29202 -66477 -28898
rect -66173 -29202 -66137 -28898
rect -65513 -29202 -65477 -28898
rect -65173 -29202 -65137 -28898
rect -64513 -29202 -64477 -28898
rect -64173 -29202 -64137 -28898
rect -63513 -29202 -63477 -28898
rect -63173 -29202 -63137 -28898
rect -62513 -29202 -62477 -28898
rect -62173 -29202 -62137 -28898
rect -61513 -29202 -61477 -28898
rect -61173 -29202 -61137 -28898
rect -60513 -29202 -60477 -28898
rect -60173 -29202 -60137 -28898
rect -59513 -29202 -59477 -28898
rect -59173 -29202 -59137 -28898
rect -58513 -29202 -58477 -28898
rect -58173 -29202 -58137 -28898
rect -57513 -29202 -57477 -28898
rect -57173 -29202 -57137 -28898
rect -56513 -29202 -56477 -28898
rect -56173 -29202 -56137 -28898
rect -55513 -29202 -55477 -28898
rect -55173 -29202 -55137 -28898
rect -54513 -29202 -54477 -28898
rect -54173 -29202 -54137 -28898
rect -53513 -29202 -53477 -28898
rect -53173 -29202 -53137 -28898
rect -52513 -29202 -52477 -28898
rect -52173 -29202 -52137 -28898
rect -51513 -29202 -51477 -28898
rect -51173 -29202 -51137 -28898
rect -50513 -29202 -50477 -28898
rect -50173 -29202 -50137 -28898
rect -49513 -29202 -49477 -28898
rect -49173 -29202 -49137 -28898
rect -48833 -29202 -48825 -28898
rect -74825 -29210 -48825 -29202
rect 8275 -28898 34275 -28890
rect 8275 -29202 8283 -28898
rect 8587 -29202 8623 -28898
rect 8927 -29202 8963 -28898
rect 9587 -29202 9623 -28898
rect 9927 -29202 9963 -28898
rect 10587 -29202 10623 -28898
rect 10927 -29202 10963 -28898
rect 11587 -29202 11623 -28898
rect 11927 -29202 11963 -28898
rect 12587 -29202 12623 -28898
rect 12927 -29202 12963 -28898
rect 13587 -29202 13623 -28898
rect 13927 -29202 13963 -28898
rect 14587 -29202 14623 -28898
rect 14927 -29202 14963 -28898
rect 15587 -29202 15623 -28898
rect 15927 -29202 15963 -28898
rect 16587 -29202 16623 -28898
rect 16927 -29202 16963 -28898
rect 17587 -29202 17623 -28898
rect 17927 -29202 17963 -28898
rect 18587 -29202 18623 -28898
rect 18927 -29202 18963 -28898
rect 19587 -29202 19623 -28898
rect 19927 -29202 19963 -28898
rect 20587 -29202 20623 -28898
rect 20927 -29202 20963 -28898
rect 21587 -29202 21623 -28898
rect 21927 -29202 21963 -28898
rect 22587 -29202 22623 -28898
rect 22927 -29202 22963 -28898
rect 23587 -29202 23623 -28898
rect 23927 -29202 23963 -28898
rect 24587 -29202 24623 -28898
rect 24927 -29202 24963 -28898
rect 25587 -29202 25623 -28898
rect 25927 -29202 25963 -28898
rect 26587 -29202 26623 -28898
rect 26927 -29202 26963 -28898
rect 27587 -29202 27623 -28898
rect 27927 -29202 27963 -28898
rect 28587 -29202 28623 -28898
rect 28927 -29202 28963 -28898
rect 29587 -29202 29623 -28898
rect 29927 -29202 29963 -28898
rect 30587 -29202 30623 -28898
rect 30927 -29202 30963 -28898
rect 31587 -29202 31623 -28898
rect 31927 -29202 31963 -28898
rect 32587 -29202 32623 -28898
rect 32927 -29202 32963 -28898
rect 33587 -29202 33623 -28898
rect 33927 -29202 33963 -28898
rect 34267 -29202 34275 -28898
rect 8275 -29210 34275 -29202
rect -74485 -29238 -74165 -29210
rect -74485 -29862 -74477 -29238
rect -74173 -29862 -74165 -29238
rect -74485 -29890 -74165 -29862
rect -73485 -29238 -73165 -29210
rect -73485 -29862 -73477 -29238
rect -73173 -29862 -73165 -29238
rect -73485 -29890 -73165 -29862
rect -72485 -29238 -72165 -29210
rect -72485 -29862 -72477 -29238
rect -72173 -29862 -72165 -29238
rect -72485 -29890 -72165 -29862
rect -71485 -29238 -71165 -29210
rect -71485 -29862 -71477 -29238
rect -71173 -29862 -71165 -29238
rect -71485 -29890 -71165 -29862
rect -70485 -29238 -70165 -29210
rect -70485 -29862 -70477 -29238
rect -70173 -29862 -70165 -29238
rect -70485 -29890 -70165 -29862
rect -69485 -29238 -69165 -29210
rect -69485 -29862 -69477 -29238
rect -69173 -29862 -69165 -29238
rect -69485 -29890 -69165 -29862
rect -68485 -29238 -68165 -29210
rect -68485 -29862 -68477 -29238
rect -68173 -29862 -68165 -29238
rect -68485 -29890 -68165 -29862
rect -67485 -29238 -67165 -29210
rect -67485 -29862 -67477 -29238
rect -67173 -29862 -67165 -29238
rect -67485 -29890 -67165 -29862
rect -66485 -29238 -66165 -29210
rect -66485 -29862 -66477 -29238
rect -66173 -29862 -66165 -29238
rect -66485 -29890 -66165 -29862
rect -65485 -29238 -65165 -29210
rect -65485 -29862 -65477 -29238
rect -65173 -29862 -65165 -29238
rect -65485 -29890 -65165 -29862
rect -64485 -29238 -64165 -29210
rect -64485 -29862 -64477 -29238
rect -64173 -29862 -64165 -29238
rect -64485 -29890 -64165 -29862
rect -63485 -29238 -63165 -29210
rect -63485 -29862 -63477 -29238
rect -63173 -29862 -63165 -29238
rect -63485 -29890 -63165 -29862
rect -62485 -29238 -62165 -29210
rect -62485 -29862 -62477 -29238
rect -62173 -29862 -62165 -29238
rect -62485 -29890 -62165 -29862
rect -61485 -29238 -61165 -29210
rect -61485 -29862 -61477 -29238
rect -61173 -29862 -61165 -29238
rect -61485 -29890 -61165 -29862
rect -60485 -29238 -60165 -29210
rect -60485 -29862 -60477 -29238
rect -60173 -29862 -60165 -29238
rect -60485 -29890 -60165 -29862
rect -59485 -29238 -59165 -29210
rect -59485 -29862 -59477 -29238
rect -59173 -29862 -59165 -29238
rect -59485 -29890 -59165 -29862
rect -58485 -29238 -58165 -29210
rect -58485 -29862 -58477 -29238
rect -58173 -29862 -58165 -29238
rect -58485 -29890 -58165 -29862
rect -57485 -29238 -57165 -29210
rect -57485 -29862 -57477 -29238
rect -57173 -29862 -57165 -29238
rect -57485 -29890 -57165 -29862
rect -56485 -29238 -56165 -29210
rect -56485 -29862 -56477 -29238
rect -56173 -29862 -56165 -29238
rect -56485 -29890 -56165 -29862
rect -55485 -29238 -55165 -29210
rect -55485 -29862 -55477 -29238
rect -55173 -29862 -55165 -29238
rect -55485 -29890 -55165 -29862
rect -54485 -29238 -54165 -29210
rect -54485 -29862 -54477 -29238
rect -54173 -29862 -54165 -29238
rect -54485 -29890 -54165 -29862
rect -53485 -29238 -53165 -29210
rect -53485 -29862 -53477 -29238
rect -53173 -29862 -53165 -29238
rect -53485 -29890 -53165 -29862
rect -52485 -29238 -52165 -29210
rect -52485 -29862 -52477 -29238
rect -52173 -29862 -52165 -29238
rect -52485 -29890 -52165 -29862
rect -51485 -29238 -51165 -29210
rect -51485 -29862 -51477 -29238
rect -51173 -29862 -51165 -29238
rect -51485 -29890 -51165 -29862
rect -50485 -29238 -50165 -29210
rect -50485 -29862 -50477 -29238
rect -50173 -29862 -50165 -29238
rect -50485 -29890 -50165 -29862
rect -49485 -29238 -49165 -29210
rect -49485 -29862 -49477 -29238
rect -49173 -29862 -49165 -29238
rect -49485 -29890 -49165 -29862
rect 8615 -29238 8935 -29210
rect 8615 -29862 8623 -29238
rect 8927 -29862 8935 -29238
rect 8615 -29890 8935 -29862
rect 9615 -29238 9935 -29210
rect 9615 -29862 9623 -29238
rect 9927 -29862 9935 -29238
rect 9615 -29890 9935 -29862
rect 10615 -29238 10935 -29210
rect 10615 -29862 10623 -29238
rect 10927 -29862 10935 -29238
rect 10615 -29890 10935 -29862
rect 11615 -29238 11935 -29210
rect 11615 -29862 11623 -29238
rect 11927 -29862 11935 -29238
rect 11615 -29890 11935 -29862
rect 12615 -29238 12935 -29210
rect 12615 -29862 12623 -29238
rect 12927 -29862 12935 -29238
rect 12615 -29890 12935 -29862
rect 13615 -29238 13935 -29210
rect 13615 -29862 13623 -29238
rect 13927 -29862 13935 -29238
rect 13615 -29890 13935 -29862
rect 14615 -29238 14935 -29210
rect 14615 -29862 14623 -29238
rect 14927 -29862 14935 -29238
rect 14615 -29890 14935 -29862
rect 15615 -29238 15935 -29210
rect 15615 -29862 15623 -29238
rect 15927 -29862 15935 -29238
rect 15615 -29890 15935 -29862
rect 16615 -29238 16935 -29210
rect 16615 -29862 16623 -29238
rect 16927 -29862 16935 -29238
rect 16615 -29890 16935 -29862
rect 17615 -29238 17935 -29210
rect 17615 -29862 17623 -29238
rect 17927 -29862 17935 -29238
rect 17615 -29890 17935 -29862
rect 18615 -29238 18935 -29210
rect 18615 -29862 18623 -29238
rect 18927 -29862 18935 -29238
rect 18615 -29890 18935 -29862
rect 19615 -29238 19935 -29210
rect 19615 -29862 19623 -29238
rect 19927 -29862 19935 -29238
rect 19615 -29890 19935 -29862
rect 20615 -29238 20935 -29210
rect 20615 -29862 20623 -29238
rect 20927 -29862 20935 -29238
rect 20615 -29890 20935 -29862
rect 21615 -29238 21935 -29210
rect 21615 -29862 21623 -29238
rect 21927 -29862 21935 -29238
rect 21615 -29890 21935 -29862
rect 22615 -29238 22935 -29210
rect 22615 -29862 22623 -29238
rect 22927 -29862 22935 -29238
rect 22615 -29890 22935 -29862
rect 23615 -29238 23935 -29210
rect 23615 -29862 23623 -29238
rect 23927 -29862 23935 -29238
rect 23615 -29890 23935 -29862
rect 24615 -29238 24935 -29210
rect 24615 -29862 24623 -29238
rect 24927 -29862 24935 -29238
rect 24615 -29890 24935 -29862
rect 25615 -29238 25935 -29210
rect 25615 -29862 25623 -29238
rect 25927 -29862 25935 -29238
rect 25615 -29890 25935 -29862
rect 26615 -29238 26935 -29210
rect 26615 -29862 26623 -29238
rect 26927 -29862 26935 -29238
rect 26615 -29890 26935 -29862
rect 27615 -29238 27935 -29210
rect 27615 -29862 27623 -29238
rect 27927 -29862 27935 -29238
rect 27615 -29890 27935 -29862
rect 28615 -29238 28935 -29210
rect 28615 -29862 28623 -29238
rect 28927 -29862 28935 -29238
rect 28615 -29890 28935 -29862
rect 29615 -29238 29935 -29210
rect 29615 -29862 29623 -29238
rect 29927 -29862 29935 -29238
rect 29615 -29890 29935 -29862
rect 30615 -29238 30935 -29210
rect 30615 -29862 30623 -29238
rect 30927 -29862 30935 -29238
rect 30615 -29890 30935 -29862
rect 31615 -29238 31935 -29210
rect 31615 -29862 31623 -29238
rect 31927 -29862 31935 -29238
rect 31615 -29890 31935 -29862
rect 32615 -29238 32935 -29210
rect 32615 -29862 32623 -29238
rect 32927 -29862 32935 -29238
rect 32615 -29890 32935 -29862
rect 33615 -29238 33935 -29210
rect 33615 -29862 33623 -29238
rect 33927 -29862 33935 -29238
rect 33615 -29890 33935 -29862
rect -74825 -29898 -48825 -29890
rect -74825 -30202 -74817 -29898
rect -74513 -30202 -74477 -29898
rect -74173 -30202 -74137 -29898
rect -73513 -30202 -73477 -29898
rect -73173 -30202 -73137 -29898
rect -72513 -30202 -72477 -29898
rect -72173 -30202 -72137 -29898
rect -71513 -30202 -71477 -29898
rect -71173 -30202 -71137 -29898
rect -70513 -30202 -70477 -29898
rect -70173 -30202 -70137 -29898
rect -69513 -30202 -69477 -29898
rect -69173 -30202 -69137 -29898
rect -68513 -30202 -68477 -29898
rect -68173 -30202 -68137 -29898
rect -67513 -30202 -67477 -29898
rect -67173 -30202 -67137 -29898
rect -66513 -30202 -66477 -29898
rect -66173 -30202 -66137 -29898
rect -65513 -30202 -65477 -29898
rect -65173 -30202 -65137 -29898
rect -64513 -30202 -64477 -29898
rect -64173 -30202 -64137 -29898
rect -63513 -30202 -63477 -29898
rect -63173 -30202 -63137 -29898
rect -62513 -30202 -62477 -29898
rect -62173 -30202 -62137 -29898
rect -61513 -30202 -61477 -29898
rect -61173 -30202 -61137 -29898
rect -60513 -30202 -60477 -29898
rect -60173 -30202 -60137 -29898
rect -59513 -30202 -59477 -29898
rect -59173 -30202 -59137 -29898
rect -58513 -30202 -58477 -29898
rect -58173 -30202 -58137 -29898
rect -57513 -30202 -57477 -29898
rect -57173 -30202 -57137 -29898
rect -56513 -30202 -56477 -29898
rect -56173 -30202 -56137 -29898
rect -55513 -30202 -55477 -29898
rect -55173 -30202 -55137 -29898
rect -54513 -30202 -54477 -29898
rect -54173 -30202 -54137 -29898
rect -53513 -30202 -53477 -29898
rect -53173 -30202 -53137 -29898
rect -52513 -30202 -52477 -29898
rect -52173 -30202 -52137 -29898
rect -51513 -30202 -51477 -29898
rect -51173 -30202 -51137 -29898
rect -50513 -30202 -50477 -29898
rect -50173 -30202 -50137 -29898
rect -49513 -30202 -49477 -29898
rect -49173 -30202 -49137 -29898
rect -48833 -30202 -48825 -29898
rect -74825 -30210 -48825 -30202
rect 8275 -29898 34275 -29890
rect 8275 -30202 8283 -29898
rect 8587 -30202 8623 -29898
rect 8927 -30202 8963 -29898
rect 9587 -30202 9623 -29898
rect 9927 -30202 9963 -29898
rect 10587 -30202 10623 -29898
rect 10927 -30202 10963 -29898
rect 11587 -30202 11623 -29898
rect 11927 -30202 11963 -29898
rect 12587 -30202 12623 -29898
rect 12927 -30202 12963 -29898
rect 13587 -30202 13623 -29898
rect 13927 -30202 13963 -29898
rect 14587 -30202 14623 -29898
rect 14927 -30202 14963 -29898
rect 15587 -30202 15623 -29898
rect 15927 -30202 15963 -29898
rect 16587 -30202 16623 -29898
rect 16927 -30202 16963 -29898
rect 17587 -30202 17623 -29898
rect 17927 -30202 17963 -29898
rect 18587 -30202 18623 -29898
rect 18927 -30202 18963 -29898
rect 19587 -30202 19623 -29898
rect 19927 -30202 19963 -29898
rect 20587 -30202 20623 -29898
rect 20927 -30202 20963 -29898
rect 21587 -30202 21623 -29898
rect 21927 -30202 21963 -29898
rect 22587 -30202 22623 -29898
rect 22927 -30202 22963 -29898
rect 23587 -30202 23623 -29898
rect 23927 -30202 23963 -29898
rect 24587 -30202 24623 -29898
rect 24927 -30202 24963 -29898
rect 25587 -30202 25623 -29898
rect 25927 -30202 25963 -29898
rect 26587 -30202 26623 -29898
rect 26927 -30202 26963 -29898
rect 27587 -30202 27623 -29898
rect 27927 -30202 27963 -29898
rect 28587 -30202 28623 -29898
rect 28927 -30202 28963 -29898
rect 29587 -30202 29623 -29898
rect 29927 -30202 29963 -29898
rect 30587 -30202 30623 -29898
rect 30927 -30202 30963 -29898
rect 31587 -30202 31623 -29898
rect 31927 -30202 31963 -29898
rect 32587 -30202 32623 -29898
rect 32927 -30202 32963 -29898
rect 33587 -30202 33623 -29898
rect 33927 -30202 33963 -29898
rect 34267 -30202 34275 -29898
rect 8275 -30210 34275 -30202
rect -74485 -30238 -74165 -30210
rect -74485 -30862 -74477 -30238
rect -74173 -30862 -74165 -30238
rect -74485 -30890 -74165 -30862
rect -73485 -30238 -73165 -30210
rect -73485 -30862 -73477 -30238
rect -73173 -30862 -73165 -30238
rect -73485 -30890 -73165 -30862
rect -72485 -30238 -72165 -30210
rect -72485 -30862 -72477 -30238
rect -72173 -30862 -72165 -30238
rect -72485 -30890 -72165 -30862
rect -71485 -30238 -71165 -30210
rect -71485 -30862 -71477 -30238
rect -71173 -30862 -71165 -30238
rect -71485 -30890 -71165 -30862
rect -70485 -30238 -70165 -30210
rect -70485 -30862 -70477 -30238
rect -70173 -30862 -70165 -30238
rect -70485 -30890 -70165 -30862
rect -69485 -30238 -69165 -30210
rect -69485 -30862 -69477 -30238
rect -69173 -30862 -69165 -30238
rect -69485 -30890 -69165 -30862
rect -68485 -30238 -68165 -30210
rect -68485 -30862 -68477 -30238
rect -68173 -30862 -68165 -30238
rect -68485 -30890 -68165 -30862
rect -67485 -30238 -67165 -30210
rect -67485 -30862 -67477 -30238
rect -67173 -30862 -67165 -30238
rect -67485 -30890 -67165 -30862
rect -66485 -30238 -66165 -30210
rect -66485 -30862 -66477 -30238
rect -66173 -30862 -66165 -30238
rect -66485 -30890 -66165 -30862
rect -65485 -30238 -65165 -30210
rect -65485 -30862 -65477 -30238
rect -65173 -30862 -65165 -30238
rect -65485 -30890 -65165 -30862
rect -64485 -30238 -64165 -30210
rect -64485 -30862 -64477 -30238
rect -64173 -30862 -64165 -30238
rect -64485 -30890 -64165 -30862
rect -63485 -30238 -63165 -30210
rect -63485 -30862 -63477 -30238
rect -63173 -30862 -63165 -30238
rect -63485 -30890 -63165 -30862
rect -62485 -30238 -62165 -30210
rect -62485 -30862 -62477 -30238
rect -62173 -30862 -62165 -30238
rect -62485 -30890 -62165 -30862
rect -61485 -30238 -61165 -30210
rect -61485 -30862 -61477 -30238
rect -61173 -30862 -61165 -30238
rect -61485 -30890 -61165 -30862
rect -60485 -30238 -60165 -30210
rect -60485 -30862 -60477 -30238
rect -60173 -30862 -60165 -30238
rect -60485 -30890 -60165 -30862
rect -59485 -30238 -59165 -30210
rect -59485 -30862 -59477 -30238
rect -59173 -30862 -59165 -30238
rect -59485 -30890 -59165 -30862
rect -58485 -30238 -58165 -30210
rect -58485 -30862 -58477 -30238
rect -58173 -30862 -58165 -30238
rect -58485 -30890 -58165 -30862
rect -57485 -30238 -57165 -30210
rect -57485 -30862 -57477 -30238
rect -57173 -30862 -57165 -30238
rect -57485 -30890 -57165 -30862
rect -56485 -30238 -56165 -30210
rect -56485 -30862 -56477 -30238
rect -56173 -30862 -56165 -30238
rect -56485 -30890 -56165 -30862
rect -55485 -30238 -55165 -30210
rect -55485 -30862 -55477 -30238
rect -55173 -30862 -55165 -30238
rect -55485 -30890 -55165 -30862
rect -54485 -30238 -54165 -30210
rect -54485 -30862 -54477 -30238
rect -54173 -30862 -54165 -30238
rect -54485 -30890 -54165 -30862
rect -53485 -30238 -53165 -30210
rect -53485 -30862 -53477 -30238
rect -53173 -30862 -53165 -30238
rect -53485 -30890 -53165 -30862
rect -52485 -30238 -52165 -30210
rect -52485 -30862 -52477 -30238
rect -52173 -30862 -52165 -30238
rect -52485 -30890 -52165 -30862
rect -51485 -30238 -51165 -30210
rect -51485 -30862 -51477 -30238
rect -51173 -30862 -51165 -30238
rect -51485 -30890 -51165 -30862
rect -50485 -30238 -50165 -30210
rect -50485 -30862 -50477 -30238
rect -50173 -30862 -50165 -30238
rect -50485 -30890 -50165 -30862
rect -49485 -30238 -49165 -30210
rect -49485 -30862 -49477 -30238
rect -49173 -30862 -49165 -30238
rect -49485 -30890 -49165 -30862
rect 8615 -30238 8935 -30210
rect 8615 -30862 8623 -30238
rect 8927 -30862 8935 -30238
rect 8615 -30890 8935 -30862
rect 9615 -30238 9935 -30210
rect 9615 -30862 9623 -30238
rect 9927 -30862 9935 -30238
rect 9615 -30890 9935 -30862
rect 10615 -30238 10935 -30210
rect 10615 -30862 10623 -30238
rect 10927 -30862 10935 -30238
rect 10615 -30890 10935 -30862
rect 11615 -30238 11935 -30210
rect 11615 -30862 11623 -30238
rect 11927 -30862 11935 -30238
rect 11615 -30890 11935 -30862
rect 12615 -30238 12935 -30210
rect 12615 -30862 12623 -30238
rect 12927 -30862 12935 -30238
rect 12615 -30890 12935 -30862
rect 13615 -30238 13935 -30210
rect 13615 -30862 13623 -30238
rect 13927 -30862 13935 -30238
rect 13615 -30890 13935 -30862
rect 14615 -30238 14935 -30210
rect 14615 -30862 14623 -30238
rect 14927 -30862 14935 -30238
rect 14615 -30890 14935 -30862
rect 15615 -30238 15935 -30210
rect 15615 -30862 15623 -30238
rect 15927 -30862 15935 -30238
rect 15615 -30890 15935 -30862
rect 16615 -30238 16935 -30210
rect 16615 -30862 16623 -30238
rect 16927 -30862 16935 -30238
rect 16615 -30890 16935 -30862
rect 17615 -30238 17935 -30210
rect 17615 -30862 17623 -30238
rect 17927 -30862 17935 -30238
rect 17615 -30890 17935 -30862
rect 18615 -30238 18935 -30210
rect 18615 -30862 18623 -30238
rect 18927 -30862 18935 -30238
rect 18615 -30890 18935 -30862
rect 19615 -30238 19935 -30210
rect 19615 -30862 19623 -30238
rect 19927 -30862 19935 -30238
rect 19615 -30890 19935 -30862
rect 20615 -30238 20935 -30210
rect 20615 -30862 20623 -30238
rect 20927 -30862 20935 -30238
rect 20615 -30890 20935 -30862
rect 21615 -30238 21935 -30210
rect 21615 -30862 21623 -30238
rect 21927 -30862 21935 -30238
rect 21615 -30890 21935 -30862
rect 22615 -30238 22935 -30210
rect 22615 -30862 22623 -30238
rect 22927 -30862 22935 -30238
rect 22615 -30890 22935 -30862
rect 23615 -30238 23935 -30210
rect 23615 -30862 23623 -30238
rect 23927 -30862 23935 -30238
rect 23615 -30890 23935 -30862
rect 24615 -30238 24935 -30210
rect 24615 -30862 24623 -30238
rect 24927 -30862 24935 -30238
rect 24615 -30890 24935 -30862
rect 25615 -30238 25935 -30210
rect 25615 -30862 25623 -30238
rect 25927 -30862 25935 -30238
rect 25615 -30890 25935 -30862
rect 26615 -30238 26935 -30210
rect 26615 -30862 26623 -30238
rect 26927 -30862 26935 -30238
rect 26615 -30890 26935 -30862
rect 27615 -30238 27935 -30210
rect 27615 -30862 27623 -30238
rect 27927 -30862 27935 -30238
rect 27615 -30890 27935 -30862
rect 28615 -30238 28935 -30210
rect 28615 -30862 28623 -30238
rect 28927 -30862 28935 -30238
rect 28615 -30890 28935 -30862
rect 29615 -30238 29935 -30210
rect 29615 -30862 29623 -30238
rect 29927 -30862 29935 -30238
rect 29615 -30890 29935 -30862
rect 30615 -30238 30935 -30210
rect 30615 -30862 30623 -30238
rect 30927 -30862 30935 -30238
rect 30615 -30890 30935 -30862
rect 31615 -30238 31935 -30210
rect 31615 -30862 31623 -30238
rect 31927 -30862 31935 -30238
rect 31615 -30890 31935 -30862
rect 32615 -30238 32935 -30210
rect 32615 -30862 32623 -30238
rect 32927 -30862 32935 -30238
rect 32615 -30890 32935 -30862
rect 33615 -30238 33935 -30210
rect 33615 -30862 33623 -30238
rect 33927 -30862 33935 -30238
rect 33615 -30890 33935 -30862
rect -74825 -30898 -48825 -30890
rect -74825 -31202 -74817 -30898
rect -74513 -31202 -74477 -30898
rect -74173 -31202 -74137 -30898
rect -73513 -31202 -73477 -30898
rect -73173 -31202 -73137 -30898
rect -72513 -31202 -72477 -30898
rect -72173 -31202 -72137 -30898
rect -71513 -31202 -71477 -30898
rect -71173 -31202 -71137 -30898
rect -70513 -31202 -70477 -30898
rect -70173 -31202 -70137 -30898
rect -69513 -31202 -69477 -30898
rect -69173 -31202 -69137 -30898
rect -68513 -31202 -68477 -30898
rect -68173 -31202 -68137 -30898
rect -67513 -31202 -67477 -30898
rect -67173 -31202 -67137 -30898
rect -66513 -31202 -66477 -30898
rect -66173 -31202 -66137 -30898
rect -65513 -31202 -65477 -30898
rect -65173 -31202 -65137 -30898
rect -64513 -31202 -64477 -30898
rect -64173 -31202 -64137 -30898
rect -63513 -31202 -63477 -30898
rect -63173 -31202 -63137 -30898
rect -62513 -31202 -62477 -30898
rect -62173 -31202 -62137 -30898
rect -61513 -31202 -61477 -30898
rect -61173 -31202 -61137 -30898
rect -60513 -31202 -60477 -30898
rect -60173 -31202 -60137 -30898
rect -59513 -31202 -59477 -30898
rect -59173 -31202 -59137 -30898
rect -58513 -31202 -58477 -30898
rect -58173 -31202 -58137 -30898
rect -57513 -31202 -57477 -30898
rect -57173 -31202 -57137 -30898
rect -56513 -31202 -56477 -30898
rect -56173 -31202 -56137 -30898
rect -55513 -31202 -55477 -30898
rect -55173 -31202 -55137 -30898
rect -54513 -31202 -54477 -30898
rect -54173 -31202 -54137 -30898
rect -53513 -31202 -53477 -30898
rect -53173 -31202 -53137 -30898
rect -52513 -31202 -52477 -30898
rect -52173 -31202 -52137 -30898
rect -51513 -31202 -51477 -30898
rect -51173 -31202 -51137 -30898
rect -50513 -31202 -50477 -30898
rect -50173 -31202 -50137 -30898
rect -49513 -31202 -49477 -30898
rect -49173 -31202 -49137 -30898
rect -48833 -31202 -48825 -30898
rect -74825 -31210 -48825 -31202
rect 8275 -30898 34275 -30890
rect 8275 -31202 8283 -30898
rect 8587 -31202 8623 -30898
rect 8927 -31202 8963 -30898
rect 9587 -31202 9623 -30898
rect 9927 -31202 9963 -30898
rect 10587 -31202 10623 -30898
rect 10927 -31202 10963 -30898
rect 11587 -31202 11623 -30898
rect 11927 -31202 11963 -30898
rect 12587 -31202 12623 -30898
rect 12927 -31202 12963 -30898
rect 13587 -31202 13623 -30898
rect 13927 -31202 13963 -30898
rect 14587 -31202 14623 -30898
rect 14927 -31202 14963 -30898
rect 15587 -31202 15623 -30898
rect 15927 -31202 15963 -30898
rect 16587 -31202 16623 -30898
rect 16927 -31202 16963 -30898
rect 17587 -31202 17623 -30898
rect 17927 -31202 17963 -30898
rect 18587 -31202 18623 -30898
rect 18927 -31202 18963 -30898
rect 19587 -31202 19623 -30898
rect 19927 -31202 19963 -30898
rect 20587 -31202 20623 -30898
rect 20927 -31202 20963 -30898
rect 21587 -31202 21623 -30898
rect 21927 -31202 21963 -30898
rect 22587 -31202 22623 -30898
rect 22927 -31202 22963 -30898
rect 23587 -31202 23623 -30898
rect 23927 -31202 23963 -30898
rect 24587 -31202 24623 -30898
rect 24927 -31202 24963 -30898
rect 25587 -31202 25623 -30898
rect 25927 -31202 25963 -30898
rect 26587 -31202 26623 -30898
rect 26927 -31202 26963 -30898
rect 27587 -31202 27623 -30898
rect 27927 -31202 27963 -30898
rect 28587 -31202 28623 -30898
rect 28927 -31202 28963 -30898
rect 29587 -31202 29623 -30898
rect 29927 -31202 29963 -30898
rect 30587 -31202 30623 -30898
rect 30927 -31202 30963 -30898
rect 31587 -31202 31623 -30898
rect 31927 -31202 31963 -30898
rect 32587 -31202 32623 -30898
rect 32927 -31202 32963 -30898
rect 33587 -31202 33623 -30898
rect 33927 -31202 33963 -30898
rect 34267 -31202 34275 -30898
rect 8275 -31210 34275 -31202
rect -74485 -31238 -74165 -31210
rect -74485 -31862 -74477 -31238
rect -74173 -31862 -74165 -31238
rect -74485 -31890 -74165 -31862
rect -73485 -31238 -73165 -31210
rect -73485 -31862 -73477 -31238
rect -73173 -31862 -73165 -31238
rect -73485 -31890 -73165 -31862
rect -72485 -31238 -72165 -31210
rect -72485 -31862 -72477 -31238
rect -72173 -31862 -72165 -31238
rect -72485 -31890 -72165 -31862
rect -71485 -31238 -71165 -31210
rect -71485 -31862 -71477 -31238
rect -71173 -31862 -71165 -31238
rect -71485 -31890 -71165 -31862
rect -70485 -31238 -70165 -31210
rect -70485 -31862 -70477 -31238
rect -70173 -31862 -70165 -31238
rect -70485 -31890 -70165 -31862
rect -69485 -31238 -69165 -31210
rect -69485 -31862 -69477 -31238
rect -69173 -31862 -69165 -31238
rect -69485 -31890 -69165 -31862
rect -68485 -31238 -68165 -31210
rect -68485 -31862 -68477 -31238
rect -68173 -31862 -68165 -31238
rect -68485 -31890 -68165 -31862
rect -67485 -31238 -67165 -31210
rect -67485 -31862 -67477 -31238
rect -67173 -31862 -67165 -31238
rect -67485 -31890 -67165 -31862
rect -66485 -31238 -66165 -31210
rect -66485 -31862 -66477 -31238
rect -66173 -31862 -66165 -31238
rect -66485 -31890 -66165 -31862
rect -65485 -31238 -65165 -31210
rect -65485 -31862 -65477 -31238
rect -65173 -31862 -65165 -31238
rect -65485 -31890 -65165 -31862
rect -64485 -31238 -64165 -31210
rect -64485 -31862 -64477 -31238
rect -64173 -31862 -64165 -31238
rect -64485 -31890 -64165 -31862
rect -63485 -31238 -63165 -31210
rect -63485 -31862 -63477 -31238
rect -63173 -31862 -63165 -31238
rect -63485 -31890 -63165 -31862
rect -62485 -31238 -62165 -31210
rect -62485 -31862 -62477 -31238
rect -62173 -31862 -62165 -31238
rect -62485 -31890 -62165 -31862
rect -61485 -31238 -61165 -31210
rect -61485 -31862 -61477 -31238
rect -61173 -31862 -61165 -31238
rect -61485 -31890 -61165 -31862
rect -60485 -31238 -60165 -31210
rect -60485 -31862 -60477 -31238
rect -60173 -31862 -60165 -31238
rect -60485 -31890 -60165 -31862
rect -59485 -31238 -59165 -31210
rect -59485 -31862 -59477 -31238
rect -59173 -31862 -59165 -31238
rect -59485 -31890 -59165 -31862
rect -58485 -31238 -58165 -31210
rect -58485 -31862 -58477 -31238
rect -58173 -31862 -58165 -31238
rect -58485 -31890 -58165 -31862
rect -57485 -31238 -57165 -31210
rect -57485 -31862 -57477 -31238
rect -57173 -31862 -57165 -31238
rect -57485 -31890 -57165 -31862
rect -56485 -31238 -56165 -31210
rect -56485 -31862 -56477 -31238
rect -56173 -31862 -56165 -31238
rect -56485 -31890 -56165 -31862
rect -55485 -31238 -55165 -31210
rect -55485 -31862 -55477 -31238
rect -55173 -31862 -55165 -31238
rect -55485 -31890 -55165 -31862
rect -54485 -31238 -54165 -31210
rect -54485 -31862 -54477 -31238
rect -54173 -31862 -54165 -31238
rect -54485 -31890 -54165 -31862
rect -53485 -31238 -53165 -31210
rect -53485 -31862 -53477 -31238
rect -53173 -31862 -53165 -31238
rect -53485 -31890 -53165 -31862
rect -52485 -31238 -52165 -31210
rect -52485 -31862 -52477 -31238
rect -52173 -31862 -52165 -31238
rect -52485 -31890 -52165 -31862
rect -51485 -31238 -51165 -31210
rect -51485 -31862 -51477 -31238
rect -51173 -31862 -51165 -31238
rect -51485 -31890 -51165 -31862
rect -50485 -31238 -50165 -31210
rect -50485 -31862 -50477 -31238
rect -50173 -31862 -50165 -31238
rect -50485 -31890 -50165 -31862
rect -49485 -31238 -49165 -31210
rect -49485 -31862 -49477 -31238
rect -49173 -31862 -49165 -31238
rect -49485 -31890 -49165 -31862
rect 8615 -31238 8935 -31210
rect 8615 -31862 8623 -31238
rect 8927 -31862 8935 -31238
rect 8615 -31890 8935 -31862
rect 9615 -31238 9935 -31210
rect 9615 -31862 9623 -31238
rect 9927 -31862 9935 -31238
rect 9615 -31890 9935 -31862
rect 10615 -31238 10935 -31210
rect 10615 -31862 10623 -31238
rect 10927 -31862 10935 -31238
rect 10615 -31890 10935 -31862
rect 11615 -31238 11935 -31210
rect 11615 -31862 11623 -31238
rect 11927 -31862 11935 -31238
rect 11615 -31890 11935 -31862
rect 12615 -31238 12935 -31210
rect 12615 -31862 12623 -31238
rect 12927 -31862 12935 -31238
rect 12615 -31890 12935 -31862
rect 13615 -31238 13935 -31210
rect 13615 -31862 13623 -31238
rect 13927 -31862 13935 -31238
rect 13615 -31890 13935 -31862
rect 14615 -31238 14935 -31210
rect 14615 -31862 14623 -31238
rect 14927 -31862 14935 -31238
rect 14615 -31890 14935 -31862
rect 15615 -31238 15935 -31210
rect 15615 -31862 15623 -31238
rect 15927 -31862 15935 -31238
rect 15615 -31890 15935 -31862
rect 16615 -31238 16935 -31210
rect 16615 -31862 16623 -31238
rect 16927 -31862 16935 -31238
rect 16615 -31890 16935 -31862
rect 17615 -31238 17935 -31210
rect 17615 -31862 17623 -31238
rect 17927 -31862 17935 -31238
rect 17615 -31890 17935 -31862
rect 18615 -31238 18935 -31210
rect 18615 -31862 18623 -31238
rect 18927 -31862 18935 -31238
rect 18615 -31890 18935 -31862
rect 19615 -31238 19935 -31210
rect 19615 -31862 19623 -31238
rect 19927 -31862 19935 -31238
rect 19615 -31890 19935 -31862
rect 20615 -31238 20935 -31210
rect 20615 -31862 20623 -31238
rect 20927 -31862 20935 -31238
rect 20615 -31890 20935 -31862
rect 21615 -31238 21935 -31210
rect 21615 -31862 21623 -31238
rect 21927 -31862 21935 -31238
rect 21615 -31890 21935 -31862
rect 22615 -31238 22935 -31210
rect 22615 -31862 22623 -31238
rect 22927 -31862 22935 -31238
rect 22615 -31890 22935 -31862
rect 23615 -31238 23935 -31210
rect 23615 -31862 23623 -31238
rect 23927 -31862 23935 -31238
rect 23615 -31890 23935 -31862
rect 24615 -31238 24935 -31210
rect 24615 -31862 24623 -31238
rect 24927 -31862 24935 -31238
rect 24615 -31890 24935 -31862
rect 25615 -31238 25935 -31210
rect 25615 -31862 25623 -31238
rect 25927 -31862 25935 -31238
rect 25615 -31890 25935 -31862
rect 26615 -31238 26935 -31210
rect 26615 -31862 26623 -31238
rect 26927 -31862 26935 -31238
rect 26615 -31890 26935 -31862
rect 27615 -31238 27935 -31210
rect 27615 -31862 27623 -31238
rect 27927 -31862 27935 -31238
rect 27615 -31890 27935 -31862
rect 28615 -31238 28935 -31210
rect 28615 -31862 28623 -31238
rect 28927 -31862 28935 -31238
rect 28615 -31890 28935 -31862
rect 29615 -31238 29935 -31210
rect 29615 -31862 29623 -31238
rect 29927 -31862 29935 -31238
rect 29615 -31890 29935 -31862
rect 30615 -31238 30935 -31210
rect 30615 -31862 30623 -31238
rect 30927 -31862 30935 -31238
rect 30615 -31890 30935 -31862
rect 31615 -31238 31935 -31210
rect 31615 -31862 31623 -31238
rect 31927 -31862 31935 -31238
rect 31615 -31890 31935 -31862
rect 32615 -31238 32935 -31210
rect 32615 -31862 32623 -31238
rect 32927 -31862 32935 -31238
rect 32615 -31890 32935 -31862
rect 33615 -31238 33935 -31210
rect 33615 -31862 33623 -31238
rect 33927 -31862 33935 -31238
rect 33615 -31890 33935 -31862
rect -74825 -31898 -48825 -31890
rect -74825 -32202 -74817 -31898
rect -74513 -32202 -74477 -31898
rect -74173 -32202 -74137 -31898
rect -73513 -32202 -73477 -31898
rect -73173 -32202 -73137 -31898
rect -72513 -32202 -72477 -31898
rect -72173 -32202 -72137 -31898
rect -71513 -32202 -71477 -31898
rect -71173 -32202 -71137 -31898
rect -70513 -32202 -70477 -31898
rect -70173 -32202 -70137 -31898
rect -69513 -32202 -69477 -31898
rect -69173 -32202 -69137 -31898
rect -68513 -32202 -68477 -31898
rect -68173 -32202 -68137 -31898
rect -67513 -32202 -67477 -31898
rect -67173 -32202 -67137 -31898
rect -66513 -32202 -66477 -31898
rect -66173 -32202 -66137 -31898
rect -65513 -32202 -65477 -31898
rect -65173 -32202 -65137 -31898
rect -64513 -32202 -64477 -31898
rect -64173 -32202 -64137 -31898
rect -63513 -32202 -63477 -31898
rect -63173 -32202 -63137 -31898
rect -62513 -32202 -62477 -31898
rect -62173 -32202 -62137 -31898
rect -61513 -32202 -61477 -31898
rect -61173 -32202 -61137 -31898
rect -60513 -32202 -60477 -31898
rect -60173 -32202 -60137 -31898
rect -59513 -32202 -59477 -31898
rect -59173 -32202 -59137 -31898
rect -58513 -32202 -58477 -31898
rect -58173 -32202 -58137 -31898
rect -57513 -32202 -57477 -31898
rect -57173 -32202 -57137 -31898
rect -56513 -32202 -56477 -31898
rect -56173 -32202 -56137 -31898
rect -55513 -32202 -55477 -31898
rect -55173 -32202 -55137 -31898
rect -54513 -32202 -54477 -31898
rect -54173 -32202 -54137 -31898
rect -53513 -32202 -53477 -31898
rect -53173 -32202 -53137 -31898
rect -52513 -32202 -52477 -31898
rect -52173 -32202 -52137 -31898
rect -51513 -32202 -51477 -31898
rect -51173 -32202 -51137 -31898
rect -50513 -32202 -50477 -31898
rect -50173 -32202 -50137 -31898
rect -49513 -32202 -49477 -31898
rect -49173 -32202 -49137 -31898
rect -48833 -32202 -48825 -31898
rect -74825 -32210 -48825 -32202
rect 8275 -31898 34275 -31890
rect 8275 -32202 8283 -31898
rect 8587 -32202 8623 -31898
rect 8927 -32202 8963 -31898
rect 9587 -32202 9623 -31898
rect 9927 -32202 9963 -31898
rect 10587 -32202 10623 -31898
rect 10927 -32202 10963 -31898
rect 11587 -32202 11623 -31898
rect 11927 -32202 11963 -31898
rect 12587 -32202 12623 -31898
rect 12927 -32202 12963 -31898
rect 13587 -32202 13623 -31898
rect 13927 -32202 13963 -31898
rect 14587 -32202 14623 -31898
rect 14927 -32202 14963 -31898
rect 15587 -32202 15623 -31898
rect 15927 -32202 15963 -31898
rect 16587 -32202 16623 -31898
rect 16927 -32202 16963 -31898
rect 17587 -32202 17623 -31898
rect 17927 -32202 17963 -31898
rect 18587 -32202 18623 -31898
rect 18927 -32202 18963 -31898
rect 19587 -32202 19623 -31898
rect 19927 -32202 19963 -31898
rect 20587 -32202 20623 -31898
rect 20927 -32202 20963 -31898
rect 21587 -32202 21623 -31898
rect 21927 -32202 21963 -31898
rect 22587 -32202 22623 -31898
rect 22927 -32202 22963 -31898
rect 23587 -32202 23623 -31898
rect 23927 -32202 23963 -31898
rect 24587 -32202 24623 -31898
rect 24927 -32202 24963 -31898
rect 25587 -32202 25623 -31898
rect 25927 -32202 25963 -31898
rect 26587 -32202 26623 -31898
rect 26927 -32202 26963 -31898
rect 27587 -32202 27623 -31898
rect 27927 -32202 27963 -31898
rect 28587 -32202 28623 -31898
rect 28927 -32202 28963 -31898
rect 29587 -32202 29623 -31898
rect 29927 -32202 29963 -31898
rect 30587 -32202 30623 -31898
rect 30927 -32202 30963 -31898
rect 31587 -32202 31623 -31898
rect 31927 -32202 31963 -31898
rect 32587 -32202 32623 -31898
rect 32927 -32202 32963 -31898
rect 33587 -32202 33623 -31898
rect 33927 -32202 33963 -31898
rect 34267 -32202 34275 -31898
rect 8275 -32210 34275 -32202
rect -74485 -32238 -74165 -32210
rect -74485 -32862 -74477 -32238
rect -74173 -32862 -74165 -32238
rect -74485 -32890 -74165 -32862
rect -73485 -32238 -73165 -32210
rect -73485 -32862 -73477 -32238
rect -73173 -32862 -73165 -32238
rect -73485 -32890 -73165 -32862
rect -72485 -32238 -72165 -32210
rect -72485 -32862 -72477 -32238
rect -72173 -32862 -72165 -32238
rect -72485 -32890 -72165 -32862
rect -71485 -32238 -71165 -32210
rect -71485 -32862 -71477 -32238
rect -71173 -32862 -71165 -32238
rect -71485 -32890 -71165 -32862
rect -70485 -32238 -70165 -32210
rect -70485 -32862 -70477 -32238
rect -70173 -32862 -70165 -32238
rect -70485 -32890 -70165 -32862
rect -69485 -32238 -69165 -32210
rect -69485 -32862 -69477 -32238
rect -69173 -32862 -69165 -32238
rect -69485 -32890 -69165 -32862
rect -68485 -32238 -68165 -32210
rect -68485 -32862 -68477 -32238
rect -68173 -32862 -68165 -32238
rect -68485 -32890 -68165 -32862
rect -67485 -32238 -67165 -32210
rect -67485 -32862 -67477 -32238
rect -67173 -32862 -67165 -32238
rect -67485 -32890 -67165 -32862
rect -66485 -32238 -66165 -32210
rect -66485 -32862 -66477 -32238
rect -66173 -32862 -66165 -32238
rect -66485 -32890 -66165 -32862
rect -65485 -32238 -65165 -32210
rect -65485 -32862 -65477 -32238
rect -65173 -32862 -65165 -32238
rect -65485 -32890 -65165 -32862
rect -64485 -32238 -64165 -32210
rect -64485 -32862 -64477 -32238
rect -64173 -32862 -64165 -32238
rect -64485 -32890 -64165 -32862
rect -63485 -32238 -63165 -32210
rect -63485 -32862 -63477 -32238
rect -63173 -32862 -63165 -32238
rect -63485 -32890 -63165 -32862
rect -62485 -32238 -62165 -32210
rect -62485 -32862 -62477 -32238
rect -62173 -32862 -62165 -32238
rect -62485 -32890 -62165 -32862
rect -61485 -32238 -61165 -32210
rect -61485 -32862 -61477 -32238
rect -61173 -32862 -61165 -32238
rect -61485 -32890 -61165 -32862
rect -60485 -32238 -60165 -32210
rect -60485 -32862 -60477 -32238
rect -60173 -32862 -60165 -32238
rect -60485 -32890 -60165 -32862
rect -59485 -32238 -59165 -32210
rect -59485 -32862 -59477 -32238
rect -59173 -32862 -59165 -32238
rect -59485 -32890 -59165 -32862
rect -58485 -32238 -58165 -32210
rect -58485 -32862 -58477 -32238
rect -58173 -32862 -58165 -32238
rect -58485 -32890 -58165 -32862
rect -57485 -32238 -57165 -32210
rect -57485 -32862 -57477 -32238
rect -57173 -32862 -57165 -32238
rect -57485 -32890 -57165 -32862
rect -56485 -32238 -56165 -32210
rect -56485 -32862 -56477 -32238
rect -56173 -32862 -56165 -32238
rect -56485 -32890 -56165 -32862
rect -55485 -32238 -55165 -32210
rect -55485 -32862 -55477 -32238
rect -55173 -32862 -55165 -32238
rect -55485 -32890 -55165 -32862
rect -54485 -32238 -54165 -32210
rect -54485 -32862 -54477 -32238
rect -54173 -32862 -54165 -32238
rect -54485 -32890 -54165 -32862
rect -53485 -32238 -53165 -32210
rect -53485 -32862 -53477 -32238
rect -53173 -32862 -53165 -32238
rect -53485 -32890 -53165 -32862
rect -52485 -32238 -52165 -32210
rect -52485 -32862 -52477 -32238
rect -52173 -32862 -52165 -32238
rect -52485 -32890 -52165 -32862
rect -51485 -32238 -51165 -32210
rect -51485 -32862 -51477 -32238
rect -51173 -32862 -51165 -32238
rect -51485 -32890 -51165 -32862
rect -50485 -32238 -50165 -32210
rect -50485 -32862 -50477 -32238
rect -50173 -32862 -50165 -32238
rect -50485 -32890 -50165 -32862
rect -49485 -32238 -49165 -32210
rect -49485 -32862 -49477 -32238
rect -49173 -32862 -49165 -32238
rect 8615 -32238 8935 -32210
rect -49485 -32890 -49165 -32862
rect -46275 -32598 -36275 -32550
rect -74825 -32898 -48825 -32890
rect -74825 -33202 -74817 -32898
rect -74513 -33202 -74477 -32898
rect -74173 -33202 -74137 -32898
rect -73513 -33202 -73477 -32898
rect -73173 -33202 -73137 -32898
rect -72513 -33202 -72477 -32898
rect -72173 -33202 -72137 -32898
rect -71513 -33202 -71477 -32898
rect -71173 -33202 -71137 -32898
rect -70513 -33202 -70477 -32898
rect -70173 -33202 -70137 -32898
rect -69513 -33202 -69477 -32898
rect -69173 -33202 -69137 -32898
rect -68513 -33202 -68477 -32898
rect -68173 -33202 -68137 -32898
rect -67513 -33202 -67477 -32898
rect -67173 -33202 -67137 -32898
rect -66513 -33202 -66477 -32898
rect -66173 -33202 -66137 -32898
rect -65513 -33202 -65477 -32898
rect -65173 -33202 -65137 -32898
rect -64513 -33202 -64477 -32898
rect -64173 -33202 -64137 -32898
rect -63513 -33202 -63477 -32898
rect -63173 -33202 -63137 -32898
rect -62513 -33202 -62477 -32898
rect -62173 -33202 -62137 -32898
rect -61513 -33202 -61477 -32898
rect -61173 -33202 -61137 -32898
rect -60513 -33202 -60477 -32898
rect -60173 -33202 -60137 -32898
rect -59513 -33202 -59477 -32898
rect -59173 -33202 -59137 -32898
rect -58513 -33202 -58477 -32898
rect -58173 -33202 -58137 -32898
rect -57513 -33202 -57477 -32898
rect -57173 -33202 -57137 -32898
rect -56513 -33202 -56477 -32898
rect -56173 -33202 -56137 -32898
rect -55513 -33202 -55477 -32898
rect -55173 -33202 -55137 -32898
rect -54513 -33202 -54477 -32898
rect -54173 -33202 -54137 -32898
rect -53513 -33202 -53477 -32898
rect -53173 -33202 -53137 -32898
rect -52513 -33202 -52477 -32898
rect -52173 -33202 -52137 -32898
rect -51513 -33202 -51477 -32898
rect -51173 -33202 -51137 -32898
rect -50513 -33202 -50477 -32898
rect -50173 -33202 -50137 -32898
rect -49513 -33202 -49477 -32898
rect -49173 -33202 -49137 -32898
rect -48833 -33202 -48825 -32898
rect -74825 -33210 -48825 -33202
rect -74485 -33238 -74165 -33210
rect -74485 -33862 -74477 -33238
rect -74173 -33862 -74165 -33238
rect -74485 -33890 -74165 -33862
rect -73485 -33238 -73165 -33210
rect -73485 -33862 -73477 -33238
rect -73173 -33862 -73165 -33238
rect -73485 -33890 -73165 -33862
rect -72485 -33238 -72165 -33210
rect -72485 -33862 -72477 -33238
rect -72173 -33862 -72165 -33238
rect -72485 -33890 -72165 -33862
rect -71485 -33238 -71165 -33210
rect -71485 -33862 -71477 -33238
rect -71173 -33862 -71165 -33238
rect -71485 -33890 -71165 -33862
rect -70485 -33238 -70165 -33210
rect -70485 -33862 -70477 -33238
rect -70173 -33862 -70165 -33238
rect -70485 -33890 -70165 -33862
rect -69485 -33238 -69165 -33210
rect -69485 -33862 -69477 -33238
rect -69173 -33862 -69165 -33238
rect -69485 -33890 -69165 -33862
rect -68485 -33238 -68165 -33210
rect -68485 -33862 -68477 -33238
rect -68173 -33862 -68165 -33238
rect -68485 -33890 -68165 -33862
rect -67485 -33238 -67165 -33210
rect -67485 -33862 -67477 -33238
rect -67173 -33862 -67165 -33238
rect -67485 -33890 -67165 -33862
rect -66485 -33238 -66165 -33210
rect -66485 -33862 -66477 -33238
rect -66173 -33862 -66165 -33238
rect -66485 -33890 -66165 -33862
rect -65485 -33238 -65165 -33210
rect -65485 -33862 -65477 -33238
rect -65173 -33862 -65165 -33238
rect -65485 -33890 -65165 -33862
rect -64485 -33238 -64165 -33210
rect -64485 -33862 -64477 -33238
rect -64173 -33862 -64165 -33238
rect -64485 -33890 -64165 -33862
rect -63485 -33238 -63165 -33210
rect -63485 -33862 -63477 -33238
rect -63173 -33862 -63165 -33238
rect -63485 -33890 -63165 -33862
rect -62485 -33238 -62165 -33210
rect -62485 -33862 -62477 -33238
rect -62173 -33862 -62165 -33238
rect -62485 -33890 -62165 -33862
rect -61485 -33238 -61165 -33210
rect -61485 -33862 -61477 -33238
rect -61173 -33862 -61165 -33238
rect -61485 -33890 -61165 -33862
rect -60485 -33238 -60165 -33210
rect -60485 -33862 -60477 -33238
rect -60173 -33862 -60165 -33238
rect -60485 -33890 -60165 -33862
rect -59485 -33238 -59165 -33210
rect -59485 -33862 -59477 -33238
rect -59173 -33862 -59165 -33238
rect -59485 -33890 -59165 -33862
rect -58485 -33238 -58165 -33210
rect -58485 -33862 -58477 -33238
rect -58173 -33862 -58165 -33238
rect -58485 -33890 -58165 -33862
rect -57485 -33238 -57165 -33210
rect -57485 -33862 -57477 -33238
rect -57173 -33862 -57165 -33238
rect -57485 -33890 -57165 -33862
rect -56485 -33238 -56165 -33210
rect -56485 -33862 -56477 -33238
rect -56173 -33862 -56165 -33238
rect -56485 -33890 -56165 -33862
rect -55485 -33238 -55165 -33210
rect -55485 -33862 -55477 -33238
rect -55173 -33862 -55165 -33238
rect -55485 -33890 -55165 -33862
rect -54485 -33238 -54165 -33210
rect -54485 -33862 -54477 -33238
rect -54173 -33862 -54165 -33238
rect -54485 -33890 -54165 -33862
rect -53485 -33238 -53165 -33210
rect -53485 -33862 -53477 -33238
rect -53173 -33862 -53165 -33238
rect -53485 -33890 -53165 -33862
rect -52485 -33238 -52165 -33210
rect -52485 -33862 -52477 -33238
rect -52173 -33862 -52165 -33238
rect -52485 -33890 -52165 -33862
rect -51485 -33238 -51165 -33210
rect -51485 -33862 -51477 -33238
rect -51173 -33862 -51165 -33238
rect -51485 -33890 -51165 -33862
rect -50485 -33238 -50165 -33210
rect -50485 -33862 -50477 -33238
rect -50173 -33862 -50165 -33238
rect -50485 -33890 -50165 -33862
rect -49485 -33238 -49165 -33210
rect -49485 -33862 -49477 -33238
rect -49173 -33862 -49165 -33238
rect -49485 -33890 -49165 -33862
rect -74825 -33898 -48825 -33890
rect -74825 -34202 -74817 -33898
rect -74513 -34202 -74477 -33898
rect -74173 -34202 -74137 -33898
rect -73513 -34202 -73477 -33898
rect -73173 -34202 -73137 -33898
rect -72513 -34202 -72477 -33898
rect -72173 -34202 -72137 -33898
rect -71513 -34202 -71477 -33898
rect -71173 -34202 -71137 -33898
rect -70513 -34202 -70477 -33898
rect -70173 -34202 -70137 -33898
rect -69513 -34202 -69477 -33898
rect -69173 -34202 -69137 -33898
rect -68513 -34202 -68477 -33898
rect -68173 -34202 -68137 -33898
rect -67513 -34202 -67477 -33898
rect -67173 -34202 -67137 -33898
rect -66513 -34202 -66477 -33898
rect -66173 -34202 -66137 -33898
rect -65513 -34202 -65477 -33898
rect -65173 -34202 -65137 -33898
rect -64513 -34202 -64477 -33898
rect -64173 -34202 -64137 -33898
rect -63513 -34202 -63477 -33898
rect -63173 -34202 -63137 -33898
rect -62513 -34202 -62477 -33898
rect -62173 -34202 -62137 -33898
rect -61513 -34202 -61477 -33898
rect -61173 -34202 -61137 -33898
rect -60513 -34202 -60477 -33898
rect -60173 -34202 -60137 -33898
rect -59513 -34202 -59477 -33898
rect -59173 -34202 -59137 -33898
rect -58513 -34202 -58477 -33898
rect -58173 -34202 -58137 -33898
rect -57513 -34202 -57477 -33898
rect -57173 -34202 -57137 -33898
rect -56513 -34202 -56477 -33898
rect -56173 -34202 -56137 -33898
rect -55513 -34202 -55477 -33898
rect -55173 -34202 -55137 -33898
rect -54513 -34202 -54477 -33898
rect -54173 -34202 -54137 -33898
rect -53513 -34202 -53477 -33898
rect -53173 -34202 -53137 -33898
rect -52513 -34202 -52477 -33898
rect -52173 -34202 -52137 -33898
rect -51513 -34202 -51477 -33898
rect -51173 -34202 -51137 -33898
rect -50513 -34202 -50477 -33898
rect -50173 -34202 -50137 -33898
rect -49513 -34202 -49477 -33898
rect -49173 -34202 -49137 -33898
rect -48833 -34202 -48825 -33898
rect -74825 -34210 -48825 -34202
rect -74485 -34238 -74165 -34210
rect -74485 -34862 -74477 -34238
rect -74173 -34862 -74165 -34238
rect -74485 -34890 -74165 -34862
rect -73485 -34238 -73165 -34210
rect -73485 -34862 -73477 -34238
rect -73173 -34862 -73165 -34238
rect -73485 -34890 -73165 -34862
rect -72485 -34238 -72165 -34210
rect -72485 -34862 -72477 -34238
rect -72173 -34862 -72165 -34238
rect -72485 -34890 -72165 -34862
rect -71485 -34238 -71165 -34210
rect -71485 -34862 -71477 -34238
rect -71173 -34862 -71165 -34238
rect -71485 -34890 -71165 -34862
rect -70485 -34238 -70165 -34210
rect -70485 -34862 -70477 -34238
rect -70173 -34862 -70165 -34238
rect -70485 -34890 -70165 -34862
rect -69485 -34238 -69165 -34210
rect -69485 -34862 -69477 -34238
rect -69173 -34862 -69165 -34238
rect -69485 -34890 -69165 -34862
rect -68485 -34238 -68165 -34210
rect -68485 -34862 -68477 -34238
rect -68173 -34862 -68165 -34238
rect -68485 -34890 -68165 -34862
rect -67485 -34238 -67165 -34210
rect -67485 -34862 -67477 -34238
rect -67173 -34862 -67165 -34238
rect -67485 -34890 -67165 -34862
rect -66485 -34238 -66165 -34210
rect -66485 -34862 -66477 -34238
rect -66173 -34862 -66165 -34238
rect -66485 -34890 -66165 -34862
rect -65485 -34238 -65165 -34210
rect -65485 -34862 -65477 -34238
rect -65173 -34862 -65165 -34238
rect -65485 -34890 -65165 -34862
rect -64485 -34238 -64165 -34210
rect -64485 -34862 -64477 -34238
rect -64173 -34862 -64165 -34238
rect -64485 -34890 -64165 -34862
rect -63485 -34238 -63165 -34210
rect -63485 -34862 -63477 -34238
rect -63173 -34862 -63165 -34238
rect -63485 -34890 -63165 -34862
rect -62485 -34238 -62165 -34210
rect -62485 -34862 -62477 -34238
rect -62173 -34862 -62165 -34238
rect -62485 -34890 -62165 -34862
rect -61485 -34238 -61165 -34210
rect -61485 -34862 -61477 -34238
rect -61173 -34862 -61165 -34238
rect -61485 -34890 -61165 -34862
rect -60485 -34238 -60165 -34210
rect -60485 -34862 -60477 -34238
rect -60173 -34862 -60165 -34238
rect -60485 -34890 -60165 -34862
rect -59485 -34238 -59165 -34210
rect -59485 -34862 -59477 -34238
rect -59173 -34862 -59165 -34238
rect -59485 -34890 -59165 -34862
rect -58485 -34238 -58165 -34210
rect -58485 -34862 -58477 -34238
rect -58173 -34862 -58165 -34238
rect -58485 -34890 -58165 -34862
rect -57485 -34238 -57165 -34210
rect -57485 -34862 -57477 -34238
rect -57173 -34862 -57165 -34238
rect -57485 -34890 -57165 -34862
rect -56485 -34238 -56165 -34210
rect -56485 -34862 -56477 -34238
rect -56173 -34862 -56165 -34238
rect -56485 -34890 -56165 -34862
rect -55485 -34238 -55165 -34210
rect -55485 -34862 -55477 -34238
rect -55173 -34862 -55165 -34238
rect -55485 -34890 -55165 -34862
rect -54485 -34238 -54165 -34210
rect -54485 -34862 -54477 -34238
rect -54173 -34862 -54165 -34238
rect -54485 -34890 -54165 -34862
rect -53485 -34238 -53165 -34210
rect -53485 -34862 -53477 -34238
rect -53173 -34862 -53165 -34238
rect -53485 -34890 -53165 -34862
rect -52485 -34238 -52165 -34210
rect -52485 -34862 -52477 -34238
rect -52173 -34862 -52165 -34238
rect -52485 -34890 -52165 -34862
rect -51485 -34238 -51165 -34210
rect -51485 -34862 -51477 -34238
rect -51173 -34862 -51165 -34238
rect -51485 -34890 -51165 -34862
rect -50485 -34238 -50165 -34210
rect -50485 -34862 -50477 -34238
rect -50173 -34862 -50165 -34238
rect -50485 -34890 -50165 -34862
rect -49485 -34238 -49165 -34210
rect -49485 -34862 -49477 -34238
rect -49173 -34862 -49165 -34238
rect -49485 -34890 -49165 -34862
rect -74825 -34898 -48825 -34890
rect -74825 -35202 -74817 -34898
rect -74513 -35202 -74477 -34898
rect -74173 -35202 -74137 -34898
rect -73513 -35202 -73477 -34898
rect -73173 -35202 -73137 -34898
rect -72513 -35202 -72477 -34898
rect -72173 -35202 -72137 -34898
rect -71513 -35202 -71477 -34898
rect -71173 -35202 -71137 -34898
rect -70513 -35202 -70477 -34898
rect -70173 -35202 -70137 -34898
rect -69513 -35202 -69477 -34898
rect -69173 -35202 -69137 -34898
rect -68513 -35202 -68477 -34898
rect -68173 -35202 -68137 -34898
rect -67513 -35202 -67477 -34898
rect -67173 -35202 -67137 -34898
rect -66513 -35202 -66477 -34898
rect -66173 -35202 -66137 -34898
rect -65513 -35202 -65477 -34898
rect -65173 -35202 -65137 -34898
rect -64513 -35202 -64477 -34898
rect -64173 -35202 -64137 -34898
rect -63513 -35202 -63477 -34898
rect -63173 -35202 -63137 -34898
rect -62513 -35202 -62477 -34898
rect -62173 -35202 -62137 -34898
rect -61513 -35202 -61477 -34898
rect -61173 -35202 -61137 -34898
rect -60513 -35202 -60477 -34898
rect -60173 -35202 -60137 -34898
rect -59513 -35202 -59477 -34898
rect -59173 -35202 -59137 -34898
rect -58513 -35202 -58477 -34898
rect -58173 -35202 -58137 -34898
rect -57513 -35202 -57477 -34898
rect -57173 -35202 -57137 -34898
rect -56513 -35202 -56477 -34898
rect -56173 -35202 -56137 -34898
rect -55513 -35202 -55477 -34898
rect -55173 -35202 -55137 -34898
rect -54513 -35202 -54477 -34898
rect -54173 -35202 -54137 -34898
rect -53513 -35202 -53477 -34898
rect -53173 -35202 -53137 -34898
rect -52513 -35202 -52477 -34898
rect -52173 -35202 -52137 -34898
rect -51513 -35202 -51477 -34898
rect -51173 -35202 -51137 -34898
rect -50513 -35202 -50477 -34898
rect -50173 -35202 -50137 -34898
rect -49513 -35202 -49477 -34898
rect -49173 -35202 -49137 -34898
rect -48833 -35202 -48825 -34898
rect -74825 -35210 -48825 -35202
rect -74485 -35238 -74165 -35210
rect -74485 -35862 -74477 -35238
rect -74173 -35862 -74165 -35238
rect -74485 -35890 -74165 -35862
rect -73485 -35238 -73165 -35210
rect -73485 -35862 -73477 -35238
rect -73173 -35862 -73165 -35238
rect -73485 -35890 -73165 -35862
rect -72485 -35238 -72165 -35210
rect -72485 -35862 -72477 -35238
rect -72173 -35862 -72165 -35238
rect -72485 -35890 -72165 -35862
rect -71485 -35238 -71165 -35210
rect -71485 -35862 -71477 -35238
rect -71173 -35862 -71165 -35238
rect -71485 -35890 -71165 -35862
rect -70485 -35238 -70165 -35210
rect -70485 -35862 -70477 -35238
rect -70173 -35862 -70165 -35238
rect -70485 -35890 -70165 -35862
rect -69485 -35238 -69165 -35210
rect -69485 -35862 -69477 -35238
rect -69173 -35862 -69165 -35238
rect -69485 -35890 -69165 -35862
rect -68485 -35238 -68165 -35210
rect -68485 -35862 -68477 -35238
rect -68173 -35862 -68165 -35238
rect -68485 -35890 -68165 -35862
rect -67485 -35238 -67165 -35210
rect -67485 -35862 -67477 -35238
rect -67173 -35862 -67165 -35238
rect -67485 -35890 -67165 -35862
rect -66485 -35238 -66165 -35210
rect -66485 -35862 -66477 -35238
rect -66173 -35862 -66165 -35238
rect -66485 -35890 -66165 -35862
rect -65485 -35238 -65165 -35210
rect -65485 -35862 -65477 -35238
rect -65173 -35862 -65165 -35238
rect -65485 -35890 -65165 -35862
rect -64485 -35238 -64165 -35210
rect -64485 -35862 -64477 -35238
rect -64173 -35862 -64165 -35238
rect -64485 -35890 -64165 -35862
rect -63485 -35238 -63165 -35210
rect -63485 -35862 -63477 -35238
rect -63173 -35862 -63165 -35238
rect -63485 -35890 -63165 -35862
rect -62485 -35238 -62165 -35210
rect -62485 -35862 -62477 -35238
rect -62173 -35862 -62165 -35238
rect -62485 -35890 -62165 -35862
rect -61485 -35238 -61165 -35210
rect -61485 -35862 -61477 -35238
rect -61173 -35862 -61165 -35238
rect -61485 -35890 -61165 -35862
rect -60485 -35238 -60165 -35210
rect -60485 -35862 -60477 -35238
rect -60173 -35862 -60165 -35238
rect -60485 -35890 -60165 -35862
rect -59485 -35238 -59165 -35210
rect -59485 -35862 -59477 -35238
rect -59173 -35862 -59165 -35238
rect -59485 -35890 -59165 -35862
rect -58485 -35238 -58165 -35210
rect -58485 -35862 -58477 -35238
rect -58173 -35862 -58165 -35238
rect -58485 -35890 -58165 -35862
rect -57485 -35238 -57165 -35210
rect -57485 -35862 -57477 -35238
rect -57173 -35862 -57165 -35238
rect -57485 -35890 -57165 -35862
rect -56485 -35238 -56165 -35210
rect -56485 -35862 -56477 -35238
rect -56173 -35862 -56165 -35238
rect -56485 -35890 -56165 -35862
rect -55485 -35238 -55165 -35210
rect -55485 -35862 -55477 -35238
rect -55173 -35862 -55165 -35238
rect -55485 -35890 -55165 -35862
rect -54485 -35238 -54165 -35210
rect -54485 -35862 -54477 -35238
rect -54173 -35862 -54165 -35238
rect -54485 -35890 -54165 -35862
rect -53485 -35238 -53165 -35210
rect -53485 -35862 -53477 -35238
rect -53173 -35862 -53165 -35238
rect -53485 -35890 -53165 -35862
rect -52485 -35238 -52165 -35210
rect -52485 -35862 -52477 -35238
rect -52173 -35862 -52165 -35238
rect -52485 -35890 -52165 -35862
rect -51485 -35238 -51165 -35210
rect -51485 -35862 -51477 -35238
rect -51173 -35862 -51165 -35238
rect -51485 -35890 -51165 -35862
rect -50485 -35238 -50165 -35210
rect -50485 -35862 -50477 -35238
rect -50173 -35862 -50165 -35238
rect -50485 -35890 -50165 -35862
rect -49485 -35238 -49165 -35210
rect -49485 -35862 -49477 -35238
rect -49173 -35862 -49165 -35238
rect -49485 -35890 -49165 -35862
rect -74825 -35898 -48825 -35890
rect -74825 -36202 -74817 -35898
rect -74513 -36202 -74477 -35898
rect -74173 -36202 -74137 -35898
rect -73513 -36202 -73477 -35898
rect -73173 -36202 -73137 -35898
rect -72513 -36202 -72477 -35898
rect -72173 -36202 -72137 -35898
rect -71513 -36202 -71477 -35898
rect -71173 -36202 -71137 -35898
rect -70513 -36202 -70477 -35898
rect -70173 -36202 -70137 -35898
rect -69513 -36202 -69477 -35898
rect -69173 -36202 -69137 -35898
rect -68513 -36202 -68477 -35898
rect -68173 -36202 -68137 -35898
rect -67513 -36202 -67477 -35898
rect -67173 -36202 -67137 -35898
rect -66513 -36202 -66477 -35898
rect -66173 -36202 -66137 -35898
rect -65513 -36202 -65477 -35898
rect -65173 -36202 -65137 -35898
rect -64513 -36202 -64477 -35898
rect -64173 -36202 -64137 -35898
rect -63513 -36202 -63477 -35898
rect -63173 -36202 -63137 -35898
rect -62513 -36202 -62477 -35898
rect -62173 -36202 -62137 -35898
rect -61513 -36202 -61477 -35898
rect -61173 -36202 -61137 -35898
rect -60513 -36202 -60477 -35898
rect -60173 -36202 -60137 -35898
rect -59513 -36202 -59477 -35898
rect -59173 -36202 -59137 -35898
rect -58513 -36202 -58477 -35898
rect -58173 -36202 -58137 -35898
rect -57513 -36202 -57477 -35898
rect -57173 -36202 -57137 -35898
rect -56513 -36202 -56477 -35898
rect -56173 -36202 -56137 -35898
rect -55513 -36202 -55477 -35898
rect -55173 -36202 -55137 -35898
rect -54513 -36202 -54477 -35898
rect -54173 -36202 -54137 -35898
rect -53513 -36202 -53477 -35898
rect -53173 -36202 -53137 -35898
rect -52513 -36202 -52477 -35898
rect -52173 -36202 -52137 -35898
rect -51513 -36202 -51477 -35898
rect -51173 -36202 -51137 -35898
rect -50513 -36202 -50477 -35898
rect -50173 -36202 -50137 -35898
rect -49513 -36202 -49477 -35898
rect -49173 -36202 -49137 -35898
rect -48833 -36202 -48825 -35898
rect -74825 -36210 -48825 -36202
rect -74485 -36238 -74165 -36210
rect -74485 -36862 -74477 -36238
rect -74173 -36862 -74165 -36238
rect -74485 -36890 -74165 -36862
rect -73485 -36238 -73165 -36210
rect -73485 -36862 -73477 -36238
rect -73173 -36862 -73165 -36238
rect -73485 -36890 -73165 -36862
rect -72485 -36238 -72165 -36210
rect -72485 -36862 -72477 -36238
rect -72173 -36862 -72165 -36238
rect -72485 -36890 -72165 -36862
rect -71485 -36238 -71165 -36210
rect -71485 -36862 -71477 -36238
rect -71173 -36862 -71165 -36238
rect -71485 -36890 -71165 -36862
rect -70485 -36238 -70165 -36210
rect -70485 -36862 -70477 -36238
rect -70173 -36862 -70165 -36238
rect -70485 -36890 -70165 -36862
rect -69485 -36238 -69165 -36210
rect -69485 -36862 -69477 -36238
rect -69173 -36862 -69165 -36238
rect -69485 -36890 -69165 -36862
rect -68485 -36238 -68165 -36210
rect -68485 -36862 -68477 -36238
rect -68173 -36862 -68165 -36238
rect -68485 -36890 -68165 -36862
rect -67485 -36238 -67165 -36210
rect -67485 -36862 -67477 -36238
rect -67173 -36862 -67165 -36238
rect -67485 -36890 -67165 -36862
rect -66485 -36238 -66165 -36210
rect -66485 -36862 -66477 -36238
rect -66173 -36862 -66165 -36238
rect -66485 -36890 -66165 -36862
rect -65485 -36238 -65165 -36210
rect -65485 -36862 -65477 -36238
rect -65173 -36862 -65165 -36238
rect -65485 -36890 -65165 -36862
rect -64485 -36238 -64165 -36210
rect -64485 -36862 -64477 -36238
rect -64173 -36862 -64165 -36238
rect -64485 -36890 -64165 -36862
rect -63485 -36238 -63165 -36210
rect -63485 -36862 -63477 -36238
rect -63173 -36862 -63165 -36238
rect -63485 -36890 -63165 -36862
rect -62485 -36238 -62165 -36210
rect -62485 -36862 -62477 -36238
rect -62173 -36862 -62165 -36238
rect -62485 -36890 -62165 -36862
rect -61485 -36238 -61165 -36210
rect -61485 -36862 -61477 -36238
rect -61173 -36862 -61165 -36238
rect -61485 -36890 -61165 -36862
rect -60485 -36238 -60165 -36210
rect -60485 -36862 -60477 -36238
rect -60173 -36862 -60165 -36238
rect -60485 -36890 -60165 -36862
rect -59485 -36238 -59165 -36210
rect -59485 -36862 -59477 -36238
rect -59173 -36862 -59165 -36238
rect -59485 -36890 -59165 -36862
rect -58485 -36238 -58165 -36210
rect -58485 -36862 -58477 -36238
rect -58173 -36862 -58165 -36238
rect -58485 -36890 -58165 -36862
rect -57485 -36238 -57165 -36210
rect -57485 -36862 -57477 -36238
rect -57173 -36862 -57165 -36238
rect -57485 -36890 -57165 -36862
rect -56485 -36238 -56165 -36210
rect -56485 -36862 -56477 -36238
rect -56173 -36862 -56165 -36238
rect -56485 -36890 -56165 -36862
rect -55485 -36238 -55165 -36210
rect -55485 -36862 -55477 -36238
rect -55173 -36862 -55165 -36238
rect -55485 -36890 -55165 -36862
rect -54485 -36238 -54165 -36210
rect -54485 -36862 -54477 -36238
rect -54173 -36862 -54165 -36238
rect -54485 -36890 -54165 -36862
rect -53485 -36238 -53165 -36210
rect -53485 -36862 -53477 -36238
rect -53173 -36862 -53165 -36238
rect -53485 -36890 -53165 -36862
rect -52485 -36238 -52165 -36210
rect -52485 -36862 -52477 -36238
rect -52173 -36862 -52165 -36238
rect -52485 -36890 -52165 -36862
rect -51485 -36238 -51165 -36210
rect -51485 -36862 -51477 -36238
rect -51173 -36862 -51165 -36238
rect -51485 -36890 -51165 -36862
rect -50485 -36238 -50165 -36210
rect -50485 -36862 -50477 -36238
rect -50173 -36862 -50165 -36238
rect -50485 -36890 -50165 -36862
rect -49485 -36238 -49165 -36210
rect -49485 -36862 -49477 -36238
rect -49173 -36862 -49165 -36238
rect -49485 -36890 -49165 -36862
rect -74825 -36898 -48825 -36890
rect -74825 -37202 -74817 -36898
rect -74513 -37202 -74477 -36898
rect -74173 -37202 -74137 -36898
rect -73513 -37202 -73477 -36898
rect -73173 -37202 -73137 -36898
rect -72513 -37202 -72477 -36898
rect -72173 -37202 -72137 -36898
rect -71513 -37202 -71477 -36898
rect -71173 -37202 -71137 -36898
rect -70513 -37202 -70477 -36898
rect -70173 -37202 -70137 -36898
rect -69513 -37202 -69477 -36898
rect -69173 -37202 -69137 -36898
rect -68513 -37202 -68477 -36898
rect -68173 -37202 -68137 -36898
rect -67513 -37202 -67477 -36898
rect -67173 -37202 -67137 -36898
rect -66513 -37202 -66477 -36898
rect -66173 -37202 -66137 -36898
rect -65513 -37202 -65477 -36898
rect -65173 -37202 -65137 -36898
rect -64513 -37202 -64477 -36898
rect -64173 -37202 -64137 -36898
rect -63513 -37202 -63477 -36898
rect -63173 -37202 -63137 -36898
rect -62513 -37202 -62477 -36898
rect -62173 -37202 -62137 -36898
rect -61513 -37202 -61477 -36898
rect -61173 -37202 -61137 -36898
rect -60513 -37202 -60477 -36898
rect -60173 -37202 -60137 -36898
rect -59513 -37202 -59477 -36898
rect -59173 -37202 -59137 -36898
rect -58513 -37202 -58477 -36898
rect -58173 -37202 -58137 -36898
rect -57513 -37202 -57477 -36898
rect -57173 -37202 -57137 -36898
rect -56513 -37202 -56477 -36898
rect -56173 -37202 -56137 -36898
rect -55513 -37202 -55477 -36898
rect -55173 -37202 -55137 -36898
rect -54513 -37202 -54477 -36898
rect -54173 -37202 -54137 -36898
rect -53513 -37202 -53477 -36898
rect -53173 -37202 -53137 -36898
rect -52513 -37202 -52477 -36898
rect -52173 -37202 -52137 -36898
rect -51513 -37202 -51477 -36898
rect -51173 -37202 -51137 -36898
rect -50513 -37202 -50477 -36898
rect -50173 -37202 -50137 -36898
rect -49513 -37202 -49477 -36898
rect -49173 -37202 -49137 -36898
rect -48833 -37202 -48825 -36898
rect -74825 -37210 -48825 -37202
rect -74485 -37238 -74165 -37210
rect -74485 -37862 -74477 -37238
rect -74173 -37862 -74165 -37238
rect -74485 -37890 -74165 -37862
rect -73485 -37238 -73165 -37210
rect -73485 -37862 -73477 -37238
rect -73173 -37862 -73165 -37238
rect -73485 -37890 -73165 -37862
rect -72485 -37238 -72165 -37210
rect -72485 -37862 -72477 -37238
rect -72173 -37862 -72165 -37238
rect -72485 -37890 -72165 -37862
rect -71485 -37238 -71165 -37210
rect -71485 -37862 -71477 -37238
rect -71173 -37862 -71165 -37238
rect -71485 -37890 -71165 -37862
rect -70485 -37238 -70165 -37210
rect -70485 -37862 -70477 -37238
rect -70173 -37862 -70165 -37238
rect -70485 -37890 -70165 -37862
rect -69485 -37238 -69165 -37210
rect -69485 -37862 -69477 -37238
rect -69173 -37862 -69165 -37238
rect -69485 -37890 -69165 -37862
rect -68485 -37238 -68165 -37210
rect -68485 -37862 -68477 -37238
rect -68173 -37862 -68165 -37238
rect -68485 -37890 -68165 -37862
rect -67485 -37238 -67165 -37210
rect -67485 -37862 -67477 -37238
rect -67173 -37862 -67165 -37238
rect -67485 -37890 -67165 -37862
rect -66485 -37238 -66165 -37210
rect -66485 -37862 -66477 -37238
rect -66173 -37862 -66165 -37238
rect -66485 -37890 -66165 -37862
rect -65485 -37238 -65165 -37210
rect -65485 -37862 -65477 -37238
rect -65173 -37862 -65165 -37238
rect -65485 -37890 -65165 -37862
rect -64485 -37238 -64165 -37210
rect -64485 -37862 -64477 -37238
rect -64173 -37862 -64165 -37238
rect -64485 -37890 -64165 -37862
rect -63485 -37238 -63165 -37210
rect -63485 -37862 -63477 -37238
rect -63173 -37862 -63165 -37238
rect -63485 -37890 -63165 -37862
rect -62485 -37238 -62165 -37210
rect -62485 -37862 -62477 -37238
rect -62173 -37862 -62165 -37238
rect -62485 -37890 -62165 -37862
rect -61485 -37238 -61165 -37210
rect -61485 -37862 -61477 -37238
rect -61173 -37862 -61165 -37238
rect -61485 -37890 -61165 -37862
rect -60485 -37238 -60165 -37210
rect -60485 -37862 -60477 -37238
rect -60173 -37862 -60165 -37238
rect -60485 -37890 -60165 -37862
rect -59485 -37238 -59165 -37210
rect -59485 -37862 -59477 -37238
rect -59173 -37862 -59165 -37238
rect -59485 -37890 -59165 -37862
rect -58485 -37238 -58165 -37210
rect -58485 -37862 -58477 -37238
rect -58173 -37862 -58165 -37238
rect -58485 -37890 -58165 -37862
rect -57485 -37238 -57165 -37210
rect -57485 -37862 -57477 -37238
rect -57173 -37862 -57165 -37238
rect -57485 -37890 -57165 -37862
rect -56485 -37238 -56165 -37210
rect -56485 -37862 -56477 -37238
rect -56173 -37862 -56165 -37238
rect -56485 -37890 -56165 -37862
rect -55485 -37238 -55165 -37210
rect -55485 -37862 -55477 -37238
rect -55173 -37862 -55165 -37238
rect -55485 -37890 -55165 -37862
rect -54485 -37238 -54165 -37210
rect -54485 -37862 -54477 -37238
rect -54173 -37862 -54165 -37238
rect -54485 -37890 -54165 -37862
rect -53485 -37238 -53165 -37210
rect -53485 -37862 -53477 -37238
rect -53173 -37862 -53165 -37238
rect -53485 -37890 -53165 -37862
rect -52485 -37238 -52165 -37210
rect -52485 -37862 -52477 -37238
rect -52173 -37862 -52165 -37238
rect -52485 -37890 -52165 -37862
rect -51485 -37238 -51165 -37210
rect -51485 -37862 -51477 -37238
rect -51173 -37862 -51165 -37238
rect -51485 -37890 -51165 -37862
rect -50485 -37238 -50165 -37210
rect -50485 -37862 -50477 -37238
rect -50173 -37862 -50165 -37238
rect -50485 -37890 -50165 -37862
rect -49485 -37238 -49165 -37210
rect -49485 -37862 -49477 -37238
rect -49173 -37862 -49165 -37238
rect -49485 -37890 -49165 -37862
rect -74825 -37898 -48825 -37890
rect -74825 -38202 -74817 -37898
rect -74513 -38202 -74477 -37898
rect -74173 -38202 -74137 -37898
rect -73513 -38202 -73477 -37898
rect -73173 -38202 -73137 -37898
rect -72513 -38202 -72477 -37898
rect -72173 -38202 -72137 -37898
rect -71513 -38202 -71477 -37898
rect -71173 -38202 -71137 -37898
rect -70513 -38202 -70477 -37898
rect -70173 -38202 -70137 -37898
rect -69513 -38202 -69477 -37898
rect -69173 -38202 -69137 -37898
rect -68513 -38202 -68477 -37898
rect -68173 -38202 -68137 -37898
rect -67513 -38202 -67477 -37898
rect -67173 -38202 -67137 -37898
rect -66513 -38202 -66477 -37898
rect -66173 -38202 -66137 -37898
rect -65513 -38202 -65477 -37898
rect -65173 -38202 -65137 -37898
rect -64513 -38202 -64477 -37898
rect -64173 -38202 -64137 -37898
rect -63513 -38202 -63477 -37898
rect -63173 -38202 -63137 -37898
rect -62513 -38202 -62477 -37898
rect -62173 -38202 -62137 -37898
rect -61513 -38202 -61477 -37898
rect -61173 -38202 -61137 -37898
rect -60513 -38202 -60477 -37898
rect -60173 -38202 -60137 -37898
rect -59513 -38202 -59477 -37898
rect -59173 -38202 -59137 -37898
rect -58513 -38202 -58477 -37898
rect -58173 -38202 -58137 -37898
rect -57513 -38202 -57477 -37898
rect -57173 -38202 -57137 -37898
rect -56513 -38202 -56477 -37898
rect -56173 -38202 -56137 -37898
rect -55513 -38202 -55477 -37898
rect -55173 -38202 -55137 -37898
rect -54513 -38202 -54477 -37898
rect -54173 -38202 -54137 -37898
rect -53513 -38202 -53477 -37898
rect -53173 -38202 -53137 -37898
rect -52513 -38202 -52477 -37898
rect -52173 -38202 -52137 -37898
rect -51513 -38202 -51477 -37898
rect -51173 -38202 -51137 -37898
rect -50513 -38202 -50477 -37898
rect -50173 -38202 -50137 -37898
rect -49513 -38202 -49477 -37898
rect -49173 -38202 -49137 -37898
rect -48833 -38202 -48825 -37898
rect -74825 -38210 -48825 -38202
rect -74485 -38238 -74165 -38210
rect -74485 -38862 -74477 -38238
rect -74173 -38862 -74165 -38238
rect -74485 -38890 -74165 -38862
rect -73485 -38238 -73165 -38210
rect -73485 -38862 -73477 -38238
rect -73173 -38862 -73165 -38238
rect -73485 -38890 -73165 -38862
rect -72485 -38238 -72165 -38210
rect -72485 -38862 -72477 -38238
rect -72173 -38862 -72165 -38238
rect -72485 -38890 -72165 -38862
rect -71485 -38238 -71165 -38210
rect -71485 -38862 -71477 -38238
rect -71173 -38862 -71165 -38238
rect -71485 -38890 -71165 -38862
rect -70485 -38238 -70165 -38210
rect -70485 -38862 -70477 -38238
rect -70173 -38862 -70165 -38238
rect -70485 -38890 -70165 -38862
rect -69485 -38238 -69165 -38210
rect -69485 -38862 -69477 -38238
rect -69173 -38862 -69165 -38238
rect -69485 -38890 -69165 -38862
rect -68485 -38238 -68165 -38210
rect -68485 -38862 -68477 -38238
rect -68173 -38862 -68165 -38238
rect -68485 -38890 -68165 -38862
rect -67485 -38238 -67165 -38210
rect -67485 -38862 -67477 -38238
rect -67173 -38862 -67165 -38238
rect -67485 -38890 -67165 -38862
rect -66485 -38238 -66165 -38210
rect -66485 -38862 -66477 -38238
rect -66173 -38862 -66165 -38238
rect -66485 -38890 -66165 -38862
rect -65485 -38238 -65165 -38210
rect -65485 -38862 -65477 -38238
rect -65173 -38862 -65165 -38238
rect -65485 -38890 -65165 -38862
rect -64485 -38238 -64165 -38210
rect -64485 -38862 -64477 -38238
rect -64173 -38862 -64165 -38238
rect -64485 -38890 -64165 -38862
rect -63485 -38238 -63165 -38210
rect -63485 -38862 -63477 -38238
rect -63173 -38862 -63165 -38238
rect -63485 -38890 -63165 -38862
rect -62485 -38238 -62165 -38210
rect -62485 -38862 -62477 -38238
rect -62173 -38862 -62165 -38238
rect -62485 -38890 -62165 -38862
rect -61485 -38238 -61165 -38210
rect -61485 -38862 -61477 -38238
rect -61173 -38862 -61165 -38238
rect -61485 -38890 -61165 -38862
rect -60485 -38238 -60165 -38210
rect -60485 -38862 -60477 -38238
rect -60173 -38862 -60165 -38238
rect -60485 -38890 -60165 -38862
rect -59485 -38238 -59165 -38210
rect -59485 -38862 -59477 -38238
rect -59173 -38862 -59165 -38238
rect -59485 -38890 -59165 -38862
rect -58485 -38238 -58165 -38210
rect -58485 -38862 -58477 -38238
rect -58173 -38862 -58165 -38238
rect -58485 -38890 -58165 -38862
rect -57485 -38238 -57165 -38210
rect -57485 -38862 -57477 -38238
rect -57173 -38862 -57165 -38238
rect -57485 -38890 -57165 -38862
rect -56485 -38238 -56165 -38210
rect -56485 -38862 -56477 -38238
rect -56173 -38862 -56165 -38238
rect -56485 -38890 -56165 -38862
rect -55485 -38238 -55165 -38210
rect -55485 -38862 -55477 -38238
rect -55173 -38862 -55165 -38238
rect -55485 -38890 -55165 -38862
rect -54485 -38238 -54165 -38210
rect -54485 -38862 -54477 -38238
rect -54173 -38862 -54165 -38238
rect -54485 -38890 -54165 -38862
rect -53485 -38238 -53165 -38210
rect -53485 -38862 -53477 -38238
rect -53173 -38862 -53165 -38238
rect -53485 -38890 -53165 -38862
rect -52485 -38238 -52165 -38210
rect -52485 -38862 -52477 -38238
rect -52173 -38862 -52165 -38238
rect -52485 -38890 -52165 -38862
rect -51485 -38238 -51165 -38210
rect -51485 -38862 -51477 -38238
rect -51173 -38862 -51165 -38238
rect -51485 -38890 -51165 -38862
rect -50485 -38238 -50165 -38210
rect -50485 -38862 -50477 -38238
rect -50173 -38862 -50165 -38238
rect -50485 -38890 -50165 -38862
rect -49485 -38238 -49165 -38210
rect -49485 -38862 -49477 -38238
rect -49173 -38862 -49165 -38238
rect -49485 -38890 -49165 -38862
rect -74825 -38898 -48825 -38890
rect -74825 -39202 -74817 -38898
rect -74513 -39202 -74477 -38898
rect -74173 -39202 -74137 -38898
rect -73513 -39202 -73477 -38898
rect -73173 -39202 -73137 -38898
rect -72513 -39202 -72477 -38898
rect -72173 -39202 -72137 -38898
rect -71513 -39202 -71477 -38898
rect -71173 -39202 -71137 -38898
rect -70513 -39202 -70477 -38898
rect -70173 -39202 -70137 -38898
rect -69513 -39202 -69477 -38898
rect -69173 -39202 -69137 -38898
rect -68513 -39202 -68477 -38898
rect -68173 -39202 -68137 -38898
rect -67513 -39202 -67477 -38898
rect -67173 -39202 -67137 -38898
rect -66513 -39202 -66477 -38898
rect -66173 -39202 -66137 -38898
rect -65513 -39202 -65477 -38898
rect -65173 -39202 -65137 -38898
rect -64513 -39202 -64477 -38898
rect -64173 -39202 -64137 -38898
rect -63513 -39202 -63477 -38898
rect -63173 -39202 -63137 -38898
rect -62513 -39202 -62477 -38898
rect -62173 -39202 -62137 -38898
rect -61513 -39202 -61477 -38898
rect -61173 -39202 -61137 -38898
rect -60513 -39202 -60477 -38898
rect -60173 -39202 -60137 -38898
rect -59513 -39202 -59477 -38898
rect -59173 -39202 -59137 -38898
rect -58513 -39202 -58477 -38898
rect -58173 -39202 -58137 -38898
rect -57513 -39202 -57477 -38898
rect -57173 -39202 -57137 -38898
rect -56513 -39202 -56477 -38898
rect -56173 -39202 -56137 -38898
rect -55513 -39202 -55477 -38898
rect -55173 -39202 -55137 -38898
rect -54513 -39202 -54477 -38898
rect -54173 -39202 -54137 -38898
rect -53513 -39202 -53477 -38898
rect -53173 -39202 -53137 -38898
rect -52513 -39202 -52477 -38898
rect -52173 -39202 -52137 -38898
rect -51513 -39202 -51477 -38898
rect -51173 -39202 -51137 -38898
rect -50513 -39202 -50477 -38898
rect -50173 -39202 -50137 -38898
rect -49513 -39202 -49477 -38898
rect -49173 -39202 -49137 -38898
rect -48833 -39202 -48825 -38898
rect -74825 -39210 -48825 -39202
rect -74485 -39238 -74165 -39210
rect -74485 -39862 -74477 -39238
rect -74173 -39862 -74165 -39238
rect -74485 -39890 -74165 -39862
rect -73485 -39238 -73165 -39210
rect -73485 -39862 -73477 -39238
rect -73173 -39862 -73165 -39238
rect -73485 -39890 -73165 -39862
rect -72485 -39238 -72165 -39210
rect -72485 -39862 -72477 -39238
rect -72173 -39862 -72165 -39238
rect -72485 -39890 -72165 -39862
rect -71485 -39238 -71165 -39210
rect -71485 -39862 -71477 -39238
rect -71173 -39862 -71165 -39238
rect -71485 -39890 -71165 -39862
rect -70485 -39238 -70165 -39210
rect -70485 -39862 -70477 -39238
rect -70173 -39862 -70165 -39238
rect -70485 -39890 -70165 -39862
rect -69485 -39238 -69165 -39210
rect -69485 -39862 -69477 -39238
rect -69173 -39862 -69165 -39238
rect -69485 -39890 -69165 -39862
rect -68485 -39238 -68165 -39210
rect -68485 -39862 -68477 -39238
rect -68173 -39862 -68165 -39238
rect -68485 -39890 -68165 -39862
rect -67485 -39238 -67165 -39210
rect -67485 -39862 -67477 -39238
rect -67173 -39862 -67165 -39238
rect -67485 -39890 -67165 -39862
rect -66485 -39238 -66165 -39210
rect -66485 -39862 -66477 -39238
rect -66173 -39862 -66165 -39238
rect -66485 -39890 -66165 -39862
rect -65485 -39238 -65165 -39210
rect -65485 -39862 -65477 -39238
rect -65173 -39862 -65165 -39238
rect -65485 -39890 -65165 -39862
rect -64485 -39238 -64165 -39210
rect -64485 -39862 -64477 -39238
rect -64173 -39862 -64165 -39238
rect -64485 -39890 -64165 -39862
rect -63485 -39238 -63165 -39210
rect -63485 -39862 -63477 -39238
rect -63173 -39862 -63165 -39238
rect -63485 -39890 -63165 -39862
rect -62485 -39238 -62165 -39210
rect -62485 -39862 -62477 -39238
rect -62173 -39862 -62165 -39238
rect -62485 -39890 -62165 -39862
rect -61485 -39238 -61165 -39210
rect -61485 -39862 -61477 -39238
rect -61173 -39862 -61165 -39238
rect -61485 -39890 -61165 -39862
rect -60485 -39238 -60165 -39210
rect -60485 -39862 -60477 -39238
rect -60173 -39862 -60165 -39238
rect -60485 -39890 -60165 -39862
rect -59485 -39238 -59165 -39210
rect -59485 -39862 -59477 -39238
rect -59173 -39862 -59165 -39238
rect -59485 -39890 -59165 -39862
rect -58485 -39238 -58165 -39210
rect -58485 -39862 -58477 -39238
rect -58173 -39862 -58165 -39238
rect -58485 -39890 -58165 -39862
rect -57485 -39238 -57165 -39210
rect -57485 -39862 -57477 -39238
rect -57173 -39862 -57165 -39238
rect -57485 -39890 -57165 -39862
rect -56485 -39238 -56165 -39210
rect -56485 -39862 -56477 -39238
rect -56173 -39862 -56165 -39238
rect -56485 -39890 -56165 -39862
rect -55485 -39238 -55165 -39210
rect -55485 -39862 -55477 -39238
rect -55173 -39862 -55165 -39238
rect -55485 -39890 -55165 -39862
rect -54485 -39238 -54165 -39210
rect -54485 -39862 -54477 -39238
rect -54173 -39862 -54165 -39238
rect -54485 -39890 -54165 -39862
rect -53485 -39238 -53165 -39210
rect -53485 -39862 -53477 -39238
rect -53173 -39862 -53165 -39238
rect -53485 -39890 -53165 -39862
rect -52485 -39238 -52165 -39210
rect -52485 -39862 -52477 -39238
rect -52173 -39862 -52165 -39238
rect -52485 -39890 -52165 -39862
rect -51485 -39238 -51165 -39210
rect -51485 -39862 -51477 -39238
rect -51173 -39862 -51165 -39238
rect -51485 -39890 -51165 -39862
rect -50485 -39238 -50165 -39210
rect -50485 -39862 -50477 -39238
rect -50173 -39862 -50165 -39238
rect -50485 -39890 -50165 -39862
rect -49485 -39238 -49165 -39210
rect -49485 -39862 -49477 -39238
rect -49173 -39862 -49165 -39238
rect -49485 -39890 -49165 -39862
rect -74825 -39898 -48825 -39890
rect -74825 -40202 -74817 -39898
rect -74513 -40202 -74477 -39898
rect -74173 -40202 -74137 -39898
rect -73513 -40202 -73477 -39898
rect -73173 -40202 -73137 -39898
rect -72513 -40202 -72477 -39898
rect -72173 -40202 -72137 -39898
rect -71513 -40202 -71477 -39898
rect -71173 -40202 -71137 -39898
rect -70513 -40202 -70477 -39898
rect -70173 -40202 -70137 -39898
rect -69513 -40202 -69477 -39898
rect -69173 -40202 -69137 -39898
rect -68513 -40202 -68477 -39898
rect -68173 -40202 -68137 -39898
rect -67513 -40202 -67477 -39898
rect -67173 -40202 -67137 -39898
rect -66513 -40202 -66477 -39898
rect -66173 -40202 -66137 -39898
rect -65513 -40202 -65477 -39898
rect -65173 -40202 -65137 -39898
rect -64513 -40202 -64477 -39898
rect -64173 -40202 -64137 -39898
rect -63513 -40202 -63477 -39898
rect -63173 -40202 -63137 -39898
rect -62513 -40202 -62477 -39898
rect -62173 -40202 -62137 -39898
rect -61513 -40202 -61477 -39898
rect -61173 -40202 -61137 -39898
rect -60513 -40202 -60477 -39898
rect -60173 -40202 -60137 -39898
rect -59513 -40202 -59477 -39898
rect -59173 -40202 -59137 -39898
rect -58513 -40202 -58477 -39898
rect -58173 -40202 -58137 -39898
rect -57513 -40202 -57477 -39898
rect -57173 -40202 -57137 -39898
rect -56513 -40202 -56477 -39898
rect -56173 -40202 -56137 -39898
rect -55513 -40202 -55477 -39898
rect -55173 -40202 -55137 -39898
rect -54513 -40202 -54477 -39898
rect -54173 -40202 -54137 -39898
rect -53513 -40202 -53477 -39898
rect -53173 -40202 -53137 -39898
rect -52513 -40202 -52477 -39898
rect -52173 -40202 -52137 -39898
rect -51513 -40202 -51477 -39898
rect -51173 -40202 -51137 -39898
rect -50513 -40202 -50477 -39898
rect -50173 -40202 -50137 -39898
rect -49513 -40202 -49477 -39898
rect -49173 -40202 -49137 -39898
rect -48833 -40202 -48825 -39898
rect -74825 -40210 -48825 -40202
rect -74485 -40238 -74165 -40210
rect -74485 -40862 -74477 -40238
rect -74173 -40862 -74165 -40238
rect -74485 -40890 -74165 -40862
rect -73485 -40238 -73165 -40210
rect -73485 -40862 -73477 -40238
rect -73173 -40862 -73165 -40238
rect -73485 -40890 -73165 -40862
rect -72485 -40238 -72165 -40210
rect -72485 -40862 -72477 -40238
rect -72173 -40862 -72165 -40238
rect -72485 -40890 -72165 -40862
rect -71485 -40238 -71165 -40210
rect -71485 -40862 -71477 -40238
rect -71173 -40862 -71165 -40238
rect -71485 -40890 -71165 -40862
rect -70485 -40238 -70165 -40210
rect -70485 -40862 -70477 -40238
rect -70173 -40862 -70165 -40238
rect -70485 -40890 -70165 -40862
rect -69485 -40238 -69165 -40210
rect -69485 -40862 -69477 -40238
rect -69173 -40862 -69165 -40238
rect -69485 -40890 -69165 -40862
rect -68485 -40238 -68165 -40210
rect -68485 -40862 -68477 -40238
rect -68173 -40862 -68165 -40238
rect -68485 -40890 -68165 -40862
rect -67485 -40238 -67165 -40210
rect -67485 -40862 -67477 -40238
rect -67173 -40862 -67165 -40238
rect -67485 -40890 -67165 -40862
rect -66485 -40238 -66165 -40210
rect -66485 -40862 -66477 -40238
rect -66173 -40862 -66165 -40238
rect -66485 -40890 -66165 -40862
rect -65485 -40238 -65165 -40210
rect -65485 -40862 -65477 -40238
rect -65173 -40862 -65165 -40238
rect -65485 -40890 -65165 -40862
rect -64485 -40238 -64165 -40210
rect -64485 -40862 -64477 -40238
rect -64173 -40862 -64165 -40238
rect -64485 -40890 -64165 -40862
rect -63485 -40238 -63165 -40210
rect -63485 -40862 -63477 -40238
rect -63173 -40862 -63165 -40238
rect -63485 -40890 -63165 -40862
rect -62485 -40238 -62165 -40210
rect -62485 -40862 -62477 -40238
rect -62173 -40862 -62165 -40238
rect -62485 -40890 -62165 -40862
rect -61485 -40238 -61165 -40210
rect -61485 -40862 -61477 -40238
rect -61173 -40862 -61165 -40238
rect -61485 -40890 -61165 -40862
rect -60485 -40238 -60165 -40210
rect -60485 -40862 -60477 -40238
rect -60173 -40862 -60165 -40238
rect -60485 -40890 -60165 -40862
rect -59485 -40238 -59165 -40210
rect -59485 -40862 -59477 -40238
rect -59173 -40862 -59165 -40238
rect -59485 -40890 -59165 -40862
rect -58485 -40238 -58165 -40210
rect -58485 -40862 -58477 -40238
rect -58173 -40862 -58165 -40238
rect -58485 -40890 -58165 -40862
rect -57485 -40238 -57165 -40210
rect -57485 -40862 -57477 -40238
rect -57173 -40862 -57165 -40238
rect -57485 -40890 -57165 -40862
rect -56485 -40238 -56165 -40210
rect -56485 -40862 -56477 -40238
rect -56173 -40862 -56165 -40238
rect -56485 -40890 -56165 -40862
rect -55485 -40238 -55165 -40210
rect -55485 -40862 -55477 -40238
rect -55173 -40862 -55165 -40238
rect -55485 -40890 -55165 -40862
rect -54485 -40238 -54165 -40210
rect -54485 -40862 -54477 -40238
rect -54173 -40862 -54165 -40238
rect -54485 -40890 -54165 -40862
rect -53485 -40238 -53165 -40210
rect -53485 -40862 -53477 -40238
rect -53173 -40862 -53165 -40238
rect -53485 -40890 -53165 -40862
rect -52485 -40238 -52165 -40210
rect -52485 -40862 -52477 -40238
rect -52173 -40862 -52165 -40238
rect -52485 -40890 -52165 -40862
rect -51485 -40238 -51165 -40210
rect -51485 -40862 -51477 -40238
rect -51173 -40862 -51165 -40238
rect -51485 -40890 -51165 -40862
rect -50485 -40238 -50165 -40210
rect -50485 -40862 -50477 -40238
rect -50173 -40862 -50165 -40238
rect -50485 -40890 -50165 -40862
rect -49485 -40238 -49165 -40210
rect -49485 -40862 -49477 -40238
rect -49173 -40862 -49165 -40238
rect -49485 -40890 -49165 -40862
rect -74825 -40898 -48825 -40890
rect -74825 -41202 -74817 -40898
rect -74513 -41202 -74477 -40898
rect -74173 -41202 -74137 -40898
rect -73513 -41202 -73477 -40898
rect -73173 -41202 -73137 -40898
rect -72513 -41202 -72477 -40898
rect -72173 -41202 -72137 -40898
rect -71513 -41202 -71477 -40898
rect -71173 -41202 -71137 -40898
rect -70513 -41202 -70477 -40898
rect -70173 -41202 -70137 -40898
rect -69513 -41202 -69477 -40898
rect -69173 -41202 -69137 -40898
rect -68513 -41202 -68477 -40898
rect -68173 -41202 -68137 -40898
rect -67513 -41202 -67477 -40898
rect -67173 -41202 -67137 -40898
rect -66513 -41202 -66477 -40898
rect -66173 -41202 -66137 -40898
rect -65513 -41202 -65477 -40898
rect -65173 -41202 -65137 -40898
rect -64513 -41202 -64477 -40898
rect -64173 -41202 -64137 -40898
rect -63513 -41202 -63477 -40898
rect -63173 -41202 -63137 -40898
rect -62513 -41202 -62477 -40898
rect -62173 -41202 -62137 -40898
rect -61513 -41202 -61477 -40898
rect -61173 -41202 -61137 -40898
rect -60513 -41202 -60477 -40898
rect -60173 -41202 -60137 -40898
rect -59513 -41202 -59477 -40898
rect -59173 -41202 -59137 -40898
rect -58513 -41202 -58477 -40898
rect -58173 -41202 -58137 -40898
rect -57513 -41202 -57477 -40898
rect -57173 -41202 -57137 -40898
rect -56513 -41202 -56477 -40898
rect -56173 -41202 -56137 -40898
rect -55513 -41202 -55477 -40898
rect -55173 -41202 -55137 -40898
rect -54513 -41202 -54477 -40898
rect -54173 -41202 -54137 -40898
rect -53513 -41202 -53477 -40898
rect -53173 -41202 -53137 -40898
rect -52513 -41202 -52477 -40898
rect -52173 -41202 -52137 -40898
rect -51513 -41202 -51477 -40898
rect -51173 -41202 -51137 -40898
rect -50513 -41202 -50477 -40898
rect -50173 -41202 -50137 -40898
rect -49513 -41202 -49477 -40898
rect -49173 -41202 -49137 -40898
rect -48833 -41202 -48825 -40898
rect -74825 -41210 -48825 -41202
rect -74485 -41238 -74165 -41210
rect -74485 -41862 -74477 -41238
rect -74173 -41862 -74165 -41238
rect -74485 -41890 -74165 -41862
rect -73485 -41238 -73165 -41210
rect -73485 -41862 -73477 -41238
rect -73173 -41862 -73165 -41238
rect -73485 -41890 -73165 -41862
rect -72485 -41238 -72165 -41210
rect -72485 -41862 -72477 -41238
rect -72173 -41862 -72165 -41238
rect -72485 -41890 -72165 -41862
rect -71485 -41238 -71165 -41210
rect -71485 -41862 -71477 -41238
rect -71173 -41862 -71165 -41238
rect -71485 -41890 -71165 -41862
rect -70485 -41238 -70165 -41210
rect -70485 -41862 -70477 -41238
rect -70173 -41862 -70165 -41238
rect -70485 -41890 -70165 -41862
rect -69485 -41238 -69165 -41210
rect -69485 -41862 -69477 -41238
rect -69173 -41862 -69165 -41238
rect -69485 -41890 -69165 -41862
rect -68485 -41238 -68165 -41210
rect -68485 -41862 -68477 -41238
rect -68173 -41862 -68165 -41238
rect -68485 -41890 -68165 -41862
rect -67485 -41238 -67165 -41210
rect -67485 -41862 -67477 -41238
rect -67173 -41862 -67165 -41238
rect -67485 -41890 -67165 -41862
rect -66485 -41238 -66165 -41210
rect -66485 -41862 -66477 -41238
rect -66173 -41862 -66165 -41238
rect -66485 -41890 -66165 -41862
rect -65485 -41238 -65165 -41210
rect -65485 -41862 -65477 -41238
rect -65173 -41862 -65165 -41238
rect -65485 -41890 -65165 -41862
rect -64485 -41238 -64165 -41210
rect -64485 -41862 -64477 -41238
rect -64173 -41862 -64165 -41238
rect -64485 -41890 -64165 -41862
rect -63485 -41238 -63165 -41210
rect -63485 -41862 -63477 -41238
rect -63173 -41862 -63165 -41238
rect -63485 -41890 -63165 -41862
rect -62485 -41238 -62165 -41210
rect -62485 -41862 -62477 -41238
rect -62173 -41862 -62165 -41238
rect -62485 -41890 -62165 -41862
rect -61485 -41238 -61165 -41210
rect -61485 -41862 -61477 -41238
rect -61173 -41862 -61165 -41238
rect -61485 -41890 -61165 -41862
rect -60485 -41238 -60165 -41210
rect -60485 -41862 -60477 -41238
rect -60173 -41862 -60165 -41238
rect -60485 -41890 -60165 -41862
rect -59485 -41238 -59165 -41210
rect -59485 -41862 -59477 -41238
rect -59173 -41862 -59165 -41238
rect -59485 -41890 -59165 -41862
rect -58485 -41238 -58165 -41210
rect -58485 -41862 -58477 -41238
rect -58173 -41862 -58165 -41238
rect -58485 -41890 -58165 -41862
rect -57485 -41238 -57165 -41210
rect -57485 -41862 -57477 -41238
rect -57173 -41862 -57165 -41238
rect -57485 -41890 -57165 -41862
rect -56485 -41238 -56165 -41210
rect -56485 -41862 -56477 -41238
rect -56173 -41862 -56165 -41238
rect -56485 -41890 -56165 -41862
rect -55485 -41238 -55165 -41210
rect -55485 -41862 -55477 -41238
rect -55173 -41862 -55165 -41238
rect -55485 -41890 -55165 -41862
rect -54485 -41238 -54165 -41210
rect -54485 -41862 -54477 -41238
rect -54173 -41862 -54165 -41238
rect -54485 -41890 -54165 -41862
rect -53485 -41238 -53165 -41210
rect -53485 -41862 -53477 -41238
rect -53173 -41862 -53165 -41238
rect -53485 -41890 -53165 -41862
rect -52485 -41238 -52165 -41210
rect -52485 -41862 -52477 -41238
rect -52173 -41862 -52165 -41238
rect -52485 -41890 -52165 -41862
rect -51485 -41238 -51165 -41210
rect -51485 -41862 -51477 -41238
rect -51173 -41862 -51165 -41238
rect -51485 -41890 -51165 -41862
rect -50485 -41238 -50165 -41210
rect -50485 -41862 -50477 -41238
rect -50173 -41862 -50165 -41238
rect -50485 -41890 -50165 -41862
rect -49485 -41238 -49165 -41210
rect -49485 -41862 -49477 -41238
rect -49173 -41862 -49165 -41238
rect -49485 -41890 -49165 -41862
rect -74825 -41898 -48825 -41890
rect -74825 -42202 -74817 -41898
rect -74513 -42202 -74477 -41898
rect -74173 -42202 -74137 -41898
rect -73513 -42202 -73477 -41898
rect -73173 -42202 -73137 -41898
rect -72513 -42202 -72477 -41898
rect -72173 -42202 -72137 -41898
rect -71513 -42202 -71477 -41898
rect -71173 -42202 -71137 -41898
rect -70513 -42202 -70477 -41898
rect -70173 -42202 -70137 -41898
rect -69513 -42202 -69477 -41898
rect -69173 -42202 -69137 -41898
rect -68513 -42202 -68477 -41898
rect -68173 -42202 -68137 -41898
rect -67513 -42202 -67477 -41898
rect -67173 -42202 -67137 -41898
rect -66513 -42202 -66477 -41898
rect -66173 -42202 -66137 -41898
rect -65513 -42202 -65477 -41898
rect -65173 -42202 -65137 -41898
rect -64513 -42202 -64477 -41898
rect -64173 -42202 -64137 -41898
rect -63513 -42202 -63477 -41898
rect -63173 -42202 -63137 -41898
rect -62513 -42202 -62477 -41898
rect -62173 -42202 -62137 -41898
rect -61513 -42202 -61477 -41898
rect -61173 -42202 -61137 -41898
rect -60513 -42202 -60477 -41898
rect -60173 -42202 -60137 -41898
rect -59513 -42202 -59477 -41898
rect -59173 -42202 -59137 -41898
rect -58513 -42202 -58477 -41898
rect -58173 -42202 -58137 -41898
rect -57513 -42202 -57477 -41898
rect -57173 -42202 -57137 -41898
rect -56513 -42202 -56477 -41898
rect -56173 -42202 -56137 -41898
rect -55513 -42202 -55477 -41898
rect -55173 -42202 -55137 -41898
rect -54513 -42202 -54477 -41898
rect -54173 -42202 -54137 -41898
rect -53513 -42202 -53477 -41898
rect -53173 -42202 -53137 -41898
rect -52513 -42202 -52477 -41898
rect -52173 -42202 -52137 -41898
rect -51513 -42202 -51477 -41898
rect -51173 -42202 -51137 -41898
rect -50513 -42202 -50477 -41898
rect -50173 -42202 -50137 -41898
rect -49513 -42202 -49477 -41898
rect -49173 -42202 -49137 -41898
rect -48833 -42202 -48825 -41898
rect -74825 -42210 -48825 -42202
rect -74485 -42238 -74165 -42210
rect -74485 -42862 -74477 -42238
rect -74173 -42862 -74165 -42238
rect -74485 -42890 -74165 -42862
rect -73485 -42238 -73165 -42210
rect -73485 -42862 -73477 -42238
rect -73173 -42862 -73165 -42238
rect -73485 -42890 -73165 -42862
rect -72485 -42238 -72165 -42210
rect -72485 -42862 -72477 -42238
rect -72173 -42862 -72165 -42238
rect -72485 -42890 -72165 -42862
rect -71485 -42238 -71165 -42210
rect -71485 -42862 -71477 -42238
rect -71173 -42862 -71165 -42238
rect -71485 -42890 -71165 -42862
rect -70485 -42238 -70165 -42210
rect -70485 -42862 -70477 -42238
rect -70173 -42862 -70165 -42238
rect -70485 -42890 -70165 -42862
rect -69485 -42238 -69165 -42210
rect -69485 -42862 -69477 -42238
rect -69173 -42862 -69165 -42238
rect -69485 -42890 -69165 -42862
rect -68485 -42238 -68165 -42210
rect -68485 -42862 -68477 -42238
rect -68173 -42862 -68165 -42238
rect -68485 -42890 -68165 -42862
rect -67485 -42238 -67165 -42210
rect -67485 -42862 -67477 -42238
rect -67173 -42862 -67165 -42238
rect -67485 -42890 -67165 -42862
rect -66485 -42238 -66165 -42210
rect -66485 -42862 -66477 -42238
rect -66173 -42862 -66165 -42238
rect -66485 -42890 -66165 -42862
rect -65485 -42238 -65165 -42210
rect -65485 -42862 -65477 -42238
rect -65173 -42862 -65165 -42238
rect -65485 -42890 -65165 -42862
rect -64485 -42238 -64165 -42210
rect -64485 -42862 -64477 -42238
rect -64173 -42862 -64165 -42238
rect -64485 -42890 -64165 -42862
rect -63485 -42238 -63165 -42210
rect -63485 -42862 -63477 -42238
rect -63173 -42862 -63165 -42238
rect -63485 -42890 -63165 -42862
rect -62485 -42238 -62165 -42210
rect -62485 -42862 -62477 -42238
rect -62173 -42862 -62165 -42238
rect -62485 -42890 -62165 -42862
rect -61485 -42238 -61165 -42210
rect -61485 -42862 -61477 -42238
rect -61173 -42862 -61165 -42238
rect -61485 -42890 -61165 -42862
rect -60485 -42238 -60165 -42210
rect -60485 -42862 -60477 -42238
rect -60173 -42862 -60165 -42238
rect -60485 -42890 -60165 -42862
rect -59485 -42238 -59165 -42210
rect -59485 -42862 -59477 -42238
rect -59173 -42862 -59165 -42238
rect -59485 -42890 -59165 -42862
rect -58485 -42238 -58165 -42210
rect -58485 -42862 -58477 -42238
rect -58173 -42862 -58165 -42238
rect -58485 -42890 -58165 -42862
rect -57485 -42238 -57165 -42210
rect -57485 -42862 -57477 -42238
rect -57173 -42862 -57165 -42238
rect -57485 -42890 -57165 -42862
rect -56485 -42238 -56165 -42210
rect -56485 -42862 -56477 -42238
rect -56173 -42862 -56165 -42238
rect -56485 -42890 -56165 -42862
rect -55485 -42238 -55165 -42210
rect -55485 -42862 -55477 -42238
rect -55173 -42862 -55165 -42238
rect -55485 -42890 -55165 -42862
rect -54485 -42238 -54165 -42210
rect -54485 -42862 -54477 -42238
rect -54173 -42862 -54165 -42238
rect -54485 -42890 -54165 -42862
rect -53485 -42238 -53165 -42210
rect -53485 -42862 -53477 -42238
rect -53173 -42862 -53165 -42238
rect -53485 -42890 -53165 -42862
rect -52485 -42238 -52165 -42210
rect -52485 -42862 -52477 -42238
rect -52173 -42862 -52165 -42238
rect -52485 -42890 -52165 -42862
rect -51485 -42238 -51165 -42210
rect -51485 -42862 -51477 -42238
rect -51173 -42862 -51165 -42238
rect -51485 -42890 -51165 -42862
rect -50485 -42238 -50165 -42210
rect -50485 -42862 -50477 -42238
rect -50173 -42862 -50165 -42238
rect -50485 -42890 -50165 -42862
rect -49485 -42238 -49165 -42210
rect -49485 -42862 -49477 -42238
rect -49173 -42862 -49165 -42238
rect -49485 -42890 -49165 -42862
rect -74825 -42898 -48825 -42890
rect -74825 -43202 -74817 -42898
rect -74513 -43202 -74477 -42898
rect -74173 -43202 -74137 -42898
rect -73513 -43202 -73477 -42898
rect -73173 -43202 -73137 -42898
rect -72513 -43202 -72477 -42898
rect -72173 -43202 -72137 -42898
rect -71513 -43202 -71477 -42898
rect -71173 -43202 -71137 -42898
rect -70513 -43202 -70477 -42898
rect -70173 -43202 -70137 -42898
rect -69513 -43202 -69477 -42898
rect -69173 -43202 -69137 -42898
rect -68513 -43202 -68477 -42898
rect -68173 -43202 -68137 -42898
rect -67513 -43202 -67477 -42898
rect -67173 -43202 -67137 -42898
rect -66513 -43202 -66477 -42898
rect -66173 -43202 -66137 -42898
rect -65513 -43202 -65477 -42898
rect -65173 -43202 -65137 -42898
rect -64513 -43202 -64477 -42898
rect -64173 -43202 -64137 -42898
rect -63513 -43202 -63477 -42898
rect -63173 -43202 -63137 -42898
rect -62513 -43202 -62477 -42898
rect -62173 -43202 -62137 -42898
rect -61513 -43202 -61477 -42898
rect -61173 -43202 -61137 -42898
rect -60513 -43202 -60477 -42898
rect -60173 -43202 -60137 -42898
rect -59513 -43202 -59477 -42898
rect -59173 -43202 -59137 -42898
rect -58513 -43202 -58477 -42898
rect -58173 -43202 -58137 -42898
rect -57513 -43202 -57477 -42898
rect -57173 -43202 -57137 -42898
rect -56513 -43202 -56477 -42898
rect -56173 -43202 -56137 -42898
rect -55513 -43202 -55477 -42898
rect -55173 -43202 -55137 -42898
rect -54513 -43202 -54477 -42898
rect -54173 -43202 -54137 -42898
rect -53513 -43202 -53477 -42898
rect -53173 -43202 -53137 -42898
rect -52513 -43202 -52477 -42898
rect -52173 -43202 -52137 -42898
rect -51513 -43202 -51477 -42898
rect -51173 -43202 -51137 -42898
rect -50513 -43202 -50477 -42898
rect -50173 -43202 -50137 -42898
rect -49513 -43202 -49477 -42898
rect -49173 -43202 -49137 -42898
rect -48833 -43202 -48825 -42898
rect -74825 -43210 -48825 -43202
rect -74485 -43238 -74165 -43210
rect -74485 -43862 -74477 -43238
rect -74173 -43862 -74165 -43238
rect -74485 -43890 -74165 -43862
rect -73485 -43238 -73165 -43210
rect -73485 -43862 -73477 -43238
rect -73173 -43862 -73165 -43238
rect -73485 -43890 -73165 -43862
rect -72485 -43238 -72165 -43210
rect -72485 -43862 -72477 -43238
rect -72173 -43862 -72165 -43238
rect -72485 -43890 -72165 -43862
rect -71485 -43238 -71165 -43210
rect -71485 -43862 -71477 -43238
rect -71173 -43862 -71165 -43238
rect -71485 -43890 -71165 -43862
rect -70485 -43238 -70165 -43210
rect -70485 -43862 -70477 -43238
rect -70173 -43862 -70165 -43238
rect -70485 -43890 -70165 -43862
rect -69485 -43238 -69165 -43210
rect -69485 -43862 -69477 -43238
rect -69173 -43862 -69165 -43238
rect -69485 -43890 -69165 -43862
rect -68485 -43238 -68165 -43210
rect -68485 -43862 -68477 -43238
rect -68173 -43862 -68165 -43238
rect -68485 -43890 -68165 -43862
rect -67485 -43238 -67165 -43210
rect -67485 -43862 -67477 -43238
rect -67173 -43862 -67165 -43238
rect -67485 -43890 -67165 -43862
rect -66485 -43238 -66165 -43210
rect -66485 -43862 -66477 -43238
rect -66173 -43862 -66165 -43238
rect -66485 -43890 -66165 -43862
rect -65485 -43238 -65165 -43210
rect -65485 -43862 -65477 -43238
rect -65173 -43862 -65165 -43238
rect -65485 -43890 -65165 -43862
rect -64485 -43238 -64165 -43210
rect -64485 -43862 -64477 -43238
rect -64173 -43862 -64165 -43238
rect -64485 -43890 -64165 -43862
rect -63485 -43238 -63165 -43210
rect -63485 -43862 -63477 -43238
rect -63173 -43862 -63165 -43238
rect -63485 -43890 -63165 -43862
rect -62485 -43238 -62165 -43210
rect -62485 -43862 -62477 -43238
rect -62173 -43862 -62165 -43238
rect -62485 -43890 -62165 -43862
rect -61485 -43238 -61165 -43210
rect -61485 -43862 -61477 -43238
rect -61173 -43862 -61165 -43238
rect -61485 -43890 -61165 -43862
rect -60485 -43238 -60165 -43210
rect -60485 -43862 -60477 -43238
rect -60173 -43862 -60165 -43238
rect -60485 -43890 -60165 -43862
rect -59485 -43238 -59165 -43210
rect -59485 -43862 -59477 -43238
rect -59173 -43862 -59165 -43238
rect -59485 -43890 -59165 -43862
rect -58485 -43238 -58165 -43210
rect -58485 -43862 -58477 -43238
rect -58173 -43862 -58165 -43238
rect -58485 -43890 -58165 -43862
rect -57485 -43238 -57165 -43210
rect -57485 -43862 -57477 -43238
rect -57173 -43862 -57165 -43238
rect -57485 -43890 -57165 -43862
rect -56485 -43238 -56165 -43210
rect -56485 -43862 -56477 -43238
rect -56173 -43862 -56165 -43238
rect -56485 -43890 -56165 -43862
rect -55485 -43238 -55165 -43210
rect -55485 -43862 -55477 -43238
rect -55173 -43862 -55165 -43238
rect -55485 -43890 -55165 -43862
rect -54485 -43238 -54165 -43210
rect -54485 -43862 -54477 -43238
rect -54173 -43862 -54165 -43238
rect -54485 -43890 -54165 -43862
rect -53485 -43238 -53165 -43210
rect -53485 -43862 -53477 -43238
rect -53173 -43862 -53165 -43238
rect -53485 -43890 -53165 -43862
rect -52485 -43238 -52165 -43210
rect -52485 -43862 -52477 -43238
rect -52173 -43862 -52165 -43238
rect -52485 -43890 -52165 -43862
rect -51485 -43238 -51165 -43210
rect -51485 -43862 -51477 -43238
rect -51173 -43862 -51165 -43238
rect -51485 -43890 -51165 -43862
rect -50485 -43238 -50165 -43210
rect -50485 -43862 -50477 -43238
rect -50173 -43862 -50165 -43238
rect -50485 -43890 -50165 -43862
rect -49485 -43238 -49165 -43210
rect -49485 -43862 -49477 -43238
rect -49173 -43862 -49165 -43238
rect -49485 -43890 -49165 -43862
rect -74825 -43898 -48825 -43890
rect -74825 -44202 -74817 -43898
rect -74513 -44202 -74477 -43898
rect -74173 -44202 -74137 -43898
rect -73513 -44202 -73477 -43898
rect -73173 -44202 -73137 -43898
rect -72513 -44202 -72477 -43898
rect -72173 -44202 -72137 -43898
rect -71513 -44202 -71477 -43898
rect -71173 -44202 -71137 -43898
rect -70513 -44202 -70477 -43898
rect -70173 -44202 -70137 -43898
rect -69513 -44202 -69477 -43898
rect -69173 -44202 -69137 -43898
rect -68513 -44202 -68477 -43898
rect -68173 -44202 -68137 -43898
rect -67513 -44202 -67477 -43898
rect -67173 -44202 -67137 -43898
rect -66513 -44202 -66477 -43898
rect -66173 -44202 -66137 -43898
rect -65513 -44202 -65477 -43898
rect -65173 -44202 -65137 -43898
rect -64513 -44202 -64477 -43898
rect -64173 -44202 -64137 -43898
rect -63513 -44202 -63477 -43898
rect -63173 -44202 -63137 -43898
rect -62513 -44202 -62477 -43898
rect -62173 -44202 -62137 -43898
rect -61513 -44202 -61477 -43898
rect -61173 -44202 -61137 -43898
rect -60513 -44202 -60477 -43898
rect -60173 -44202 -60137 -43898
rect -59513 -44202 -59477 -43898
rect -59173 -44202 -59137 -43898
rect -58513 -44202 -58477 -43898
rect -58173 -44202 -58137 -43898
rect -57513 -44202 -57477 -43898
rect -57173 -44202 -57137 -43898
rect -56513 -44202 -56477 -43898
rect -56173 -44202 -56137 -43898
rect -55513 -44202 -55477 -43898
rect -55173 -44202 -55137 -43898
rect -54513 -44202 -54477 -43898
rect -54173 -44202 -54137 -43898
rect -53513 -44202 -53477 -43898
rect -53173 -44202 -53137 -43898
rect -52513 -44202 -52477 -43898
rect -52173 -44202 -52137 -43898
rect -51513 -44202 -51477 -43898
rect -51173 -44202 -51137 -43898
rect -50513 -44202 -50477 -43898
rect -50173 -44202 -50137 -43898
rect -49513 -44202 -49477 -43898
rect -49173 -44202 -49137 -43898
rect -48833 -44202 -48825 -43898
rect -74825 -44210 -48825 -44202
rect -74485 -44238 -74165 -44210
rect -74485 -44862 -74477 -44238
rect -74173 -44862 -74165 -44238
rect -74485 -44890 -74165 -44862
rect -73485 -44238 -73165 -44210
rect -73485 -44862 -73477 -44238
rect -73173 -44862 -73165 -44238
rect -73485 -44890 -73165 -44862
rect -72485 -44238 -72165 -44210
rect -72485 -44862 -72477 -44238
rect -72173 -44862 -72165 -44238
rect -72485 -44890 -72165 -44862
rect -71485 -44238 -71165 -44210
rect -71485 -44862 -71477 -44238
rect -71173 -44862 -71165 -44238
rect -71485 -44890 -71165 -44862
rect -70485 -44238 -70165 -44210
rect -70485 -44862 -70477 -44238
rect -70173 -44862 -70165 -44238
rect -70485 -44890 -70165 -44862
rect -69485 -44238 -69165 -44210
rect -69485 -44862 -69477 -44238
rect -69173 -44862 -69165 -44238
rect -69485 -44890 -69165 -44862
rect -68485 -44238 -68165 -44210
rect -68485 -44862 -68477 -44238
rect -68173 -44862 -68165 -44238
rect -68485 -44890 -68165 -44862
rect -67485 -44238 -67165 -44210
rect -67485 -44862 -67477 -44238
rect -67173 -44862 -67165 -44238
rect -67485 -44890 -67165 -44862
rect -66485 -44238 -66165 -44210
rect -66485 -44862 -66477 -44238
rect -66173 -44862 -66165 -44238
rect -66485 -44890 -66165 -44862
rect -65485 -44238 -65165 -44210
rect -65485 -44862 -65477 -44238
rect -65173 -44862 -65165 -44238
rect -65485 -44890 -65165 -44862
rect -64485 -44238 -64165 -44210
rect -64485 -44862 -64477 -44238
rect -64173 -44862 -64165 -44238
rect -64485 -44890 -64165 -44862
rect -63485 -44238 -63165 -44210
rect -63485 -44862 -63477 -44238
rect -63173 -44862 -63165 -44238
rect -63485 -44890 -63165 -44862
rect -62485 -44238 -62165 -44210
rect -62485 -44862 -62477 -44238
rect -62173 -44862 -62165 -44238
rect -62485 -44890 -62165 -44862
rect -61485 -44238 -61165 -44210
rect -61485 -44862 -61477 -44238
rect -61173 -44862 -61165 -44238
rect -61485 -44890 -61165 -44862
rect -60485 -44238 -60165 -44210
rect -60485 -44862 -60477 -44238
rect -60173 -44862 -60165 -44238
rect -60485 -44890 -60165 -44862
rect -59485 -44238 -59165 -44210
rect -59485 -44862 -59477 -44238
rect -59173 -44862 -59165 -44238
rect -59485 -44890 -59165 -44862
rect -58485 -44238 -58165 -44210
rect -58485 -44862 -58477 -44238
rect -58173 -44862 -58165 -44238
rect -58485 -44890 -58165 -44862
rect -57485 -44238 -57165 -44210
rect -57485 -44862 -57477 -44238
rect -57173 -44862 -57165 -44238
rect -57485 -44890 -57165 -44862
rect -56485 -44238 -56165 -44210
rect -56485 -44862 -56477 -44238
rect -56173 -44862 -56165 -44238
rect -56485 -44890 -56165 -44862
rect -55485 -44238 -55165 -44210
rect -55485 -44862 -55477 -44238
rect -55173 -44862 -55165 -44238
rect -55485 -44890 -55165 -44862
rect -54485 -44238 -54165 -44210
rect -54485 -44862 -54477 -44238
rect -54173 -44862 -54165 -44238
rect -54485 -44890 -54165 -44862
rect -53485 -44238 -53165 -44210
rect -53485 -44862 -53477 -44238
rect -53173 -44862 -53165 -44238
rect -53485 -44890 -53165 -44862
rect -52485 -44238 -52165 -44210
rect -52485 -44862 -52477 -44238
rect -52173 -44862 -52165 -44238
rect -52485 -44890 -52165 -44862
rect -51485 -44238 -51165 -44210
rect -51485 -44862 -51477 -44238
rect -51173 -44862 -51165 -44238
rect -51485 -44890 -51165 -44862
rect -50485 -44238 -50165 -44210
rect -50485 -44862 -50477 -44238
rect -50173 -44862 -50165 -44238
rect -50485 -44890 -50165 -44862
rect -49485 -44238 -49165 -44210
rect -49485 -44862 -49477 -44238
rect -49173 -44862 -49165 -44238
rect -46275 -44502 -46232 -32598
rect -36328 -44502 -36275 -32598
rect -46275 -44550 -36275 -44502
rect -4275 -32598 5725 -32550
rect -4275 -44502 -4232 -32598
rect 5672 -44502 5725 -32598
rect 8615 -32862 8623 -32238
rect 8927 -32862 8935 -32238
rect 8615 -32890 8935 -32862
rect 9615 -32238 9935 -32210
rect 9615 -32862 9623 -32238
rect 9927 -32862 9935 -32238
rect 9615 -32890 9935 -32862
rect 10615 -32238 10935 -32210
rect 10615 -32862 10623 -32238
rect 10927 -32862 10935 -32238
rect 10615 -32890 10935 -32862
rect 11615 -32238 11935 -32210
rect 11615 -32862 11623 -32238
rect 11927 -32862 11935 -32238
rect 11615 -32890 11935 -32862
rect 12615 -32238 12935 -32210
rect 12615 -32862 12623 -32238
rect 12927 -32862 12935 -32238
rect 12615 -32890 12935 -32862
rect 13615 -32238 13935 -32210
rect 13615 -32862 13623 -32238
rect 13927 -32862 13935 -32238
rect 13615 -32890 13935 -32862
rect 14615 -32238 14935 -32210
rect 14615 -32862 14623 -32238
rect 14927 -32862 14935 -32238
rect 14615 -32890 14935 -32862
rect 15615 -32238 15935 -32210
rect 15615 -32862 15623 -32238
rect 15927 -32862 15935 -32238
rect 15615 -32890 15935 -32862
rect 16615 -32238 16935 -32210
rect 16615 -32862 16623 -32238
rect 16927 -32862 16935 -32238
rect 16615 -32890 16935 -32862
rect 17615 -32238 17935 -32210
rect 17615 -32862 17623 -32238
rect 17927 -32862 17935 -32238
rect 17615 -32890 17935 -32862
rect 18615 -32238 18935 -32210
rect 18615 -32862 18623 -32238
rect 18927 -32862 18935 -32238
rect 18615 -32890 18935 -32862
rect 19615 -32238 19935 -32210
rect 19615 -32862 19623 -32238
rect 19927 -32862 19935 -32238
rect 19615 -32890 19935 -32862
rect 20615 -32238 20935 -32210
rect 20615 -32862 20623 -32238
rect 20927 -32862 20935 -32238
rect 20615 -32890 20935 -32862
rect 21615 -32238 21935 -32210
rect 21615 -32862 21623 -32238
rect 21927 -32862 21935 -32238
rect 21615 -32890 21935 -32862
rect 22615 -32238 22935 -32210
rect 22615 -32862 22623 -32238
rect 22927 -32862 22935 -32238
rect 22615 -32890 22935 -32862
rect 23615 -32238 23935 -32210
rect 23615 -32862 23623 -32238
rect 23927 -32862 23935 -32238
rect 23615 -32890 23935 -32862
rect 24615 -32238 24935 -32210
rect 24615 -32862 24623 -32238
rect 24927 -32862 24935 -32238
rect 24615 -32890 24935 -32862
rect 25615 -32238 25935 -32210
rect 25615 -32862 25623 -32238
rect 25927 -32862 25935 -32238
rect 25615 -32890 25935 -32862
rect 26615 -32238 26935 -32210
rect 26615 -32862 26623 -32238
rect 26927 -32862 26935 -32238
rect 26615 -32890 26935 -32862
rect 27615 -32238 27935 -32210
rect 27615 -32862 27623 -32238
rect 27927 -32862 27935 -32238
rect 27615 -32890 27935 -32862
rect 28615 -32238 28935 -32210
rect 28615 -32862 28623 -32238
rect 28927 -32862 28935 -32238
rect 28615 -32890 28935 -32862
rect 29615 -32238 29935 -32210
rect 29615 -32862 29623 -32238
rect 29927 -32862 29935 -32238
rect 29615 -32890 29935 -32862
rect 30615 -32238 30935 -32210
rect 30615 -32862 30623 -32238
rect 30927 -32862 30935 -32238
rect 30615 -32890 30935 -32862
rect 31615 -32238 31935 -32210
rect 31615 -32862 31623 -32238
rect 31927 -32862 31935 -32238
rect 31615 -32890 31935 -32862
rect 32615 -32238 32935 -32210
rect 32615 -32862 32623 -32238
rect 32927 -32862 32935 -32238
rect 32615 -32890 32935 -32862
rect 33615 -32238 33935 -32210
rect 33615 -32862 33623 -32238
rect 33927 -32862 33935 -32238
rect 33615 -32890 33935 -32862
rect 8275 -32898 34275 -32890
rect 8275 -33202 8283 -32898
rect 8587 -33202 8623 -32898
rect 8927 -33202 8963 -32898
rect 9587 -33202 9623 -32898
rect 9927 -33202 9963 -32898
rect 10587 -33202 10623 -32898
rect 10927 -33202 10963 -32898
rect 11587 -33202 11623 -32898
rect 11927 -33202 11963 -32898
rect 12587 -33202 12623 -32898
rect 12927 -33202 12963 -32898
rect 13587 -33202 13623 -32898
rect 13927 -33202 13963 -32898
rect 14587 -33202 14623 -32898
rect 14927 -33202 14963 -32898
rect 15587 -33202 15623 -32898
rect 15927 -33202 15963 -32898
rect 16587 -33202 16623 -32898
rect 16927 -33202 16963 -32898
rect 17587 -33202 17623 -32898
rect 17927 -33202 17963 -32898
rect 18587 -33202 18623 -32898
rect 18927 -33202 18963 -32898
rect 19587 -33202 19623 -32898
rect 19927 -33202 19963 -32898
rect 20587 -33202 20623 -32898
rect 20927 -33202 20963 -32898
rect 21587 -33202 21623 -32898
rect 21927 -33202 21963 -32898
rect 22587 -33202 22623 -32898
rect 22927 -33202 22963 -32898
rect 23587 -33202 23623 -32898
rect 23927 -33202 23963 -32898
rect 24587 -33202 24623 -32898
rect 24927 -33202 24963 -32898
rect 25587 -33202 25623 -32898
rect 25927 -33202 25963 -32898
rect 26587 -33202 26623 -32898
rect 26927 -33202 26963 -32898
rect 27587 -33202 27623 -32898
rect 27927 -33202 27963 -32898
rect 28587 -33202 28623 -32898
rect 28927 -33202 28963 -32898
rect 29587 -33202 29623 -32898
rect 29927 -33202 29963 -32898
rect 30587 -33202 30623 -32898
rect 30927 -33202 30963 -32898
rect 31587 -33202 31623 -32898
rect 31927 -33202 31963 -32898
rect 32587 -33202 32623 -32898
rect 32927 -33202 32963 -32898
rect 33587 -33202 33623 -32898
rect 33927 -33202 33963 -32898
rect 34267 -33202 34275 -32898
rect 8275 -33210 34275 -33202
rect 8615 -33238 8935 -33210
rect 8615 -33862 8623 -33238
rect 8927 -33862 8935 -33238
rect 8615 -33890 8935 -33862
rect 9615 -33238 9935 -33210
rect 9615 -33862 9623 -33238
rect 9927 -33862 9935 -33238
rect 9615 -33890 9935 -33862
rect 10615 -33238 10935 -33210
rect 10615 -33862 10623 -33238
rect 10927 -33862 10935 -33238
rect 10615 -33890 10935 -33862
rect 11615 -33238 11935 -33210
rect 11615 -33862 11623 -33238
rect 11927 -33862 11935 -33238
rect 11615 -33890 11935 -33862
rect 12615 -33238 12935 -33210
rect 12615 -33862 12623 -33238
rect 12927 -33862 12935 -33238
rect 12615 -33890 12935 -33862
rect 13615 -33238 13935 -33210
rect 13615 -33862 13623 -33238
rect 13927 -33862 13935 -33238
rect 13615 -33890 13935 -33862
rect 14615 -33238 14935 -33210
rect 14615 -33862 14623 -33238
rect 14927 -33862 14935 -33238
rect 14615 -33890 14935 -33862
rect 15615 -33238 15935 -33210
rect 15615 -33862 15623 -33238
rect 15927 -33862 15935 -33238
rect 15615 -33890 15935 -33862
rect 16615 -33238 16935 -33210
rect 16615 -33862 16623 -33238
rect 16927 -33862 16935 -33238
rect 16615 -33890 16935 -33862
rect 17615 -33238 17935 -33210
rect 17615 -33862 17623 -33238
rect 17927 -33862 17935 -33238
rect 17615 -33890 17935 -33862
rect 18615 -33238 18935 -33210
rect 18615 -33862 18623 -33238
rect 18927 -33862 18935 -33238
rect 18615 -33890 18935 -33862
rect 19615 -33238 19935 -33210
rect 19615 -33862 19623 -33238
rect 19927 -33862 19935 -33238
rect 19615 -33890 19935 -33862
rect 20615 -33238 20935 -33210
rect 20615 -33862 20623 -33238
rect 20927 -33862 20935 -33238
rect 20615 -33890 20935 -33862
rect 21615 -33238 21935 -33210
rect 21615 -33862 21623 -33238
rect 21927 -33862 21935 -33238
rect 21615 -33890 21935 -33862
rect 22615 -33238 22935 -33210
rect 22615 -33862 22623 -33238
rect 22927 -33862 22935 -33238
rect 22615 -33890 22935 -33862
rect 23615 -33238 23935 -33210
rect 23615 -33862 23623 -33238
rect 23927 -33862 23935 -33238
rect 23615 -33890 23935 -33862
rect 24615 -33238 24935 -33210
rect 24615 -33862 24623 -33238
rect 24927 -33862 24935 -33238
rect 24615 -33890 24935 -33862
rect 25615 -33238 25935 -33210
rect 25615 -33862 25623 -33238
rect 25927 -33862 25935 -33238
rect 25615 -33890 25935 -33862
rect 26615 -33238 26935 -33210
rect 26615 -33862 26623 -33238
rect 26927 -33862 26935 -33238
rect 26615 -33890 26935 -33862
rect 27615 -33238 27935 -33210
rect 27615 -33862 27623 -33238
rect 27927 -33862 27935 -33238
rect 27615 -33890 27935 -33862
rect 28615 -33238 28935 -33210
rect 28615 -33862 28623 -33238
rect 28927 -33862 28935 -33238
rect 28615 -33890 28935 -33862
rect 29615 -33238 29935 -33210
rect 29615 -33862 29623 -33238
rect 29927 -33862 29935 -33238
rect 29615 -33890 29935 -33862
rect 30615 -33238 30935 -33210
rect 30615 -33862 30623 -33238
rect 30927 -33862 30935 -33238
rect 30615 -33890 30935 -33862
rect 31615 -33238 31935 -33210
rect 31615 -33862 31623 -33238
rect 31927 -33862 31935 -33238
rect 31615 -33890 31935 -33862
rect 32615 -33238 32935 -33210
rect 32615 -33862 32623 -33238
rect 32927 -33862 32935 -33238
rect 32615 -33890 32935 -33862
rect 33615 -33238 33935 -33210
rect 33615 -33862 33623 -33238
rect 33927 -33862 33935 -33238
rect 33615 -33890 33935 -33862
rect 8275 -33898 34275 -33890
rect 8275 -34202 8283 -33898
rect 8587 -34202 8623 -33898
rect 8927 -34202 8963 -33898
rect 9587 -34202 9623 -33898
rect 9927 -34202 9963 -33898
rect 10587 -34202 10623 -33898
rect 10927 -34202 10963 -33898
rect 11587 -34202 11623 -33898
rect 11927 -34202 11963 -33898
rect 12587 -34202 12623 -33898
rect 12927 -34202 12963 -33898
rect 13587 -34202 13623 -33898
rect 13927 -34202 13963 -33898
rect 14587 -34202 14623 -33898
rect 14927 -34202 14963 -33898
rect 15587 -34202 15623 -33898
rect 15927 -34202 15963 -33898
rect 16587 -34202 16623 -33898
rect 16927 -34202 16963 -33898
rect 17587 -34202 17623 -33898
rect 17927 -34202 17963 -33898
rect 18587 -34202 18623 -33898
rect 18927 -34202 18963 -33898
rect 19587 -34202 19623 -33898
rect 19927 -34202 19963 -33898
rect 20587 -34202 20623 -33898
rect 20927 -34202 20963 -33898
rect 21587 -34202 21623 -33898
rect 21927 -34202 21963 -33898
rect 22587 -34202 22623 -33898
rect 22927 -34202 22963 -33898
rect 23587 -34202 23623 -33898
rect 23927 -34202 23963 -33898
rect 24587 -34202 24623 -33898
rect 24927 -34202 24963 -33898
rect 25587 -34202 25623 -33898
rect 25927 -34202 25963 -33898
rect 26587 -34202 26623 -33898
rect 26927 -34202 26963 -33898
rect 27587 -34202 27623 -33898
rect 27927 -34202 27963 -33898
rect 28587 -34202 28623 -33898
rect 28927 -34202 28963 -33898
rect 29587 -34202 29623 -33898
rect 29927 -34202 29963 -33898
rect 30587 -34202 30623 -33898
rect 30927 -34202 30963 -33898
rect 31587 -34202 31623 -33898
rect 31927 -34202 31963 -33898
rect 32587 -34202 32623 -33898
rect 32927 -34202 32963 -33898
rect 33587 -34202 33623 -33898
rect 33927 -34202 33963 -33898
rect 34267 -34202 34275 -33898
rect 8275 -34210 34275 -34202
rect 8615 -34238 8935 -34210
rect 8615 -34862 8623 -34238
rect 8927 -34862 8935 -34238
rect 8615 -34890 8935 -34862
rect 9615 -34238 9935 -34210
rect 9615 -34862 9623 -34238
rect 9927 -34862 9935 -34238
rect 9615 -34890 9935 -34862
rect 10615 -34238 10935 -34210
rect 10615 -34862 10623 -34238
rect 10927 -34862 10935 -34238
rect 10615 -34890 10935 -34862
rect 11615 -34238 11935 -34210
rect 11615 -34862 11623 -34238
rect 11927 -34862 11935 -34238
rect 11615 -34890 11935 -34862
rect 12615 -34238 12935 -34210
rect 12615 -34862 12623 -34238
rect 12927 -34862 12935 -34238
rect 12615 -34890 12935 -34862
rect 13615 -34238 13935 -34210
rect 13615 -34862 13623 -34238
rect 13927 -34862 13935 -34238
rect 13615 -34890 13935 -34862
rect 14615 -34238 14935 -34210
rect 14615 -34862 14623 -34238
rect 14927 -34862 14935 -34238
rect 14615 -34890 14935 -34862
rect 15615 -34238 15935 -34210
rect 15615 -34862 15623 -34238
rect 15927 -34862 15935 -34238
rect 15615 -34890 15935 -34862
rect 16615 -34238 16935 -34210
rect 16615 -34862 16623 -34238
rect 16927 -34862 16935 -34238
rect 16615 -34890 16935 -34862
rect 17615 -34238 17935 -34210
rect 17615 -34862 17623 -34238
rect 17927 -34862 17935 -34238
rect 17615 -34890 17935 -34862
rect 18615 -34238 18935 -34210
rect 18615 -34862 18623 -34238
rect 18927 -34862 18935 -34238
rect 18615 -34890 18935 -34862
rect 19615 -34238 19935 -34210
rect 19615 -34862 19623 -34238
rect 19927 -34862 19935 -34238
rect 19615 -34890 19935 -34862
rect 20615 -34238 20935 -34210
rect 20615 -34862 20623 -34238
rect 20927 -34862 20935 -34238
rect 20615 -34890 20935 -34862
rect 21615 -34238 21935 -34210
rect 21615 -34862 21623 -34238
rect 21927 -34862 21935 -34238
rect 21615 -34890 21935 -34862
rect 22615 -34238 22935 -34210
rect 22615 -34862 22623 -34238
rect 22927 -34862 22935 -34238
rect 22615 -34890 22935 -34862
rect 23615 -34238 23935 -34210
rect 23615 -34862 23623 -34238
rect 23927 -34862 23935 -34238
rect 23615 -34890 23935 -34862
rect 24615 -34238 24935 -34210
rect 24615 -34862 24623 -34238
rect 24927 -34862 24935 -34238
rect 24615 -34890 24935 -34862
rect 25615 -34238 25935 -34210
rect 25615 -34862 25623 -34238
rect 25927 -34862 25935 -34238
rect 25615 -34890 25935 -34862
rect 26615 -34238 26935 -34210
rect 26615 -34862 26623 -34238
rect 26927 -34862 26935 -34238
rect 26615 -34890 26935 -34862
rect 27615 -34238 27935 -34210
rect 27615 -34862 27623 -34238
rect 27927 -34862 27935 -34238
rect 27615 -34890 27935 -34862
rect 28615 -34238 28935 -34210
rect 28615 -34862 28623 -34238
rect 28927 -34862 28935 -34238
rect 28615 -34890 28935 -34862
rect 29615 -34238 29935 -34210
rect 29615 -34862 29623 -34238
rect 29927 -34862 29935 -34238
rect 29615 -34890 29935 -34862
rect 30615 -34238 30935 -34210
rect 30615 -34862 30623 -34238
rect 30927 -34862 30935 -34238
rect 30615 -34890 30935 -34862
rect 31615 -34238 31935 -34210
rect 31615 -34862 31623 -34238
rect 31927 -34862 31935 -34238
rect 31615 -34890 31935 -34862
rect 32615 -34238 32935 -34210
rect 32615 -34862 32623 -34238
rect 32927 -34862 32935 -34238
rect 32615 -34890 32935 -34862
rect 33615 -34238 33935 -34210
rect 33615 -34862 33623 -34238
rect 33927 -34862 33935 -34238
rect 33615 -34890 33935 -34862
rect 8275 -34898 34275 -34890
rect 8275 -35202 8283 -34898
rect 8587 -35202 8623 -34898
rect 8927 -35202 8963 -34898
rect 9587 -35202 9623 -34898
rect 9927 -35202 9963 -34898
rect 10587 -35202 10623 -34898
rect 10927 -35202 10963 -34898
rect 11587 -35202 11623 -34898
rect 11927 -35202 11963 -34898
rect 12587 -35202 12623 -34898
rect 12927 -35202 12963 -34898
rect 13587 -35202 13623 -34898
rect 13927 -35202 13963 -34898
rect 14587 -35202 14623 -34898
rect 14927 -35202 14963 -34898
rect 15587 -35202 15623 -34898
rect 15927 -35202 15963 -34898
rect 16587 -35202 16623 -34898
rect 16927 -35202 16963 -34898
rect 17587 -35202 17623 -34898
rect 17927 -35202 17963 -34898
rect 18587 -35202 18623 -34898
rect 18927 -35202 18963 -34898
rect 19587 -35202 19623 -34898
rect 19927 -35202 19963 -34898
rect 20587 -35202 20623 -34898
rect 20927 -35202 20963 -34898
rect 21587 -35202 21623 -34898
rect 21927 -35202 21963 -34898
rect 22587 -35202 22623 -34898
rect 22927 -35202 22963 -34898
rect 23587 -35202 23623 -34898
rect 23927 -35202 23963 -34898
rect 24587 -35202 24623 -34898
rect 24927 -35202 24963 -34898
rect 25587 -35202 25623 -34898
rect 25927 -35202 25963 -34898
rect 26587 -35202 26623 -34898
rect 26927 -35202 26963 -34898
rect 27587 -35202 27623 -34898
rect 27927 -35202 27963 -34898
rect 28587 -35202 28623 -34898
rect 28927 -35202 28963 -34898
rect 29587 -35202 29623 -34898
rect 29927 -35202 29963 -34898
rect 30587 -35202 30623 -34898
rect 30927 -35202 30963 -34898
rect 31587 -35202 31623 -34898
rect 31927 -35202 31963 -34898
rect 32587 -35202 32623 -34898
rect 32927 -35202 32963 -34898
rect 33587 -35202 33623 -34898
rect 33927 -35202 33963 -34898
rect 34267 -35202 34275 -34898
rect 8275 -35210 34275 -35202
rect 8615 -35238 8935 -35210
rect 8615 -35862 8623 -35238
rect 8927 -35862 8935 -35238
rect 8615 -35890 8935 -35862
rect 9615 -35238 9935 -35210
rect 9615 -35862 9623 -35238
rect 9927 -35862 9935 -35238
rect 9615 -35890 9935 -35862
rect 10615 -35238 10935 -35210
rect 10615 -35862 10623 -35238
rect 10927 -35862 10935 -35238
rect 10615 -35890 10935 -35862
rect 11615 -35238 11935 -35210
rect 11615 -35862 11623 -35238
rect 11927 -35862 11935 -35238
rect 11615 -35890 11935 -35862
rect 12615 -35238 12935 -35210
rect 12615 -35862 12623 -35238
rect 12927 -35862 12935 -35238
rect 12615 -35890 12935 -35862
rect 13615 -35238 13935 -35210
rect 13615 -35862 13623 -35238
rect 13927 -35862 13935 -35238
rect 13615 -35890 13935 -35862
rect 14615 -35238 14935 -35210
rect 14615 -35862 14623 -35238
rect 14927 -35862 14935 -35238
rect 14615 -35890 14935 -35862
rect 15615 -35238 15935 -35210
rect 15615 -35862 15623 -35238
rect 15927 -35862 15935 -35238
rect 15615 -35890 15935 -35862
rect 16615 -35238 16935 -35210
rect 16615 -35862 16623 -35238
rect 16927 -35862 16935 -35238
rect 16615 -35890 16935 -35862
rect 17615 -35238 17935 -35210
rect 17615 -35862 17623 -35238
rect 17927 -35862 17935 -35238
rect 17615 -35890 17935 -35862
rect 18615 -35238 18935 -35210
rect 18615 -35862 18623 -35238
rect 18927 -35862 18935 -35238
rect 18615 -35890 18935 -35862
rect 19615 -35238 19935 -35210
rect 19615 -35862 19623 -35238
rect 19927 -35862 19935 -35238
rect 19615 -35890 19935 -35862
rect 20615 -35238 20935 -35210
rect 20615 -35862 20623 -35238
rect 20927 -35862 20935 -35238
rect 20615 -35890 20935 -35862
rect 21615 -35238 21935 -35210
rect 21615 -35862 21623 -35238
rect 21927 -35862 21935 -35238
rect 21615 -35890 21935 -35862
rect 22615 -35238 22935 -35210
rect 22615 -35862 22623 -35238
rect 22927 -35862 22935 -35238
rect 22615 -35890 22935 -35862
rect 23615 -35238 23935 -35210
rect 23615 -35862 23623 -35238
rect 23927 -35862 23935 -35238
rect 23615 -35890 23935 -35862
rect 24615 -35238 24935 -35210
rect 24615 -35862 24623 -35238
rect 24927 -35862 24935 -35238
rect 24615 -35890 24935 -35862
rect 25615 -35238 25935 -35210
rect 25615 -35862 25623 -35238
rect 25927 -35862 25935 -35238
rect 25615 -35890 25935 -35862
rect 26615 -35238 26935 -35210
rect 26615 -35862 26623 -35238
rect 26927 -35862 26935 -35238
rect 26615 -35890 26935 -35862
rect 27615 -35238 27935 -35210
rect 27615 -35862 27623 -35238
rect 27927 -35862 27935 -35238
rect 27615 -35890 27935 -35862
rect 28615 -35238 28935 -35210
rect 28615 -35862 28623 -35238
rect 28927 -35862 28935 -35238
rect 28615 -35890 28935 -35862
rect 29615 -35238 29935 -35210
rect 29615 -35862 29623 -35238
rect 29927 -35862 29935 -35238
rect 29615 -35890 29935 -35862
rect 30615 -35238 30935 -35210
rect 30615 -35862 30623 -35238
rect 30927 -35862 30935 -35238
rect 30615 -35890 30935 -35862
rect 31615 -35238 31935 -35210
rect 31615 -35862 31623 -35238
rect 31927 -35862 31935 -35238
rect 31615 -35890 31935 -35862
rect 32615 -35238 32935 -35210
rect 32615 -35862 32623 -35238
rect 32927 -35862 32935 -35238
rect 32615 -35890 32935 -35862
rect 33615 -35238 33935 -35210
rect 33615 -35862 33623 -35238
rect 33927 -35862 33935 -35238
rect 33615 -35890 33935 -35862
rect 8275 -35898 34275 -35890
rect 8275 -36202 8283 -35898
rect 8587 -36202 8623 -35898
rect 8927 -36202 8963 -35898
rect 9587 -36202 9623 -35898
rect 9927 -36202 9963 -35898
rect 10587 -36202 10623 -35898
rect 10927 -36202 10963 -35898
rect 11587 -36202 11623 -35898
rect 11927 -36202 11963 -35898
rect 12587 -36202 12623 -35898
rect 12927 -36202 12963 -35898
rect 13587 -36202 13623 -35898
rect 13927 -36202 13963 -35898
rect 14587 -36202 14623 -35898
rect 14927 -36202 14963 -35898
rect 15587 -36202 15623 -35898
rect 15927 -36202 15963 -35898
rect 16587 -36202 16623 -35898
rect 16927 -36202 16963 -35898
rect 17587 -36202 17623 -35898
rect 17927 -36202 17963 -35898
rect 18587 -36202 18623 -35898
rect 18927 -36202 18963 -35898
rect 19587 -36202 19623 -35898
rect 19927 -36202 19963 -35898
rect 20587 -36202 20623 -35898
rect 20927 -36202 20963 -35898
rect 21587 -36202 21623 -35898
rect 21927 -36202 21963 -35898
rect 22587 -36202 22623 -35898
rect 22927 -36202 22963 -35898
rect 23587 -36202 23623 -35898
rect 23927 -36202 23963 -35898
rect 24587 -36202 24623 -35898
rect 24927 -36202 24963 -35898
rect 25587 -36202 25623 -35898
rect 25927 -36202 25963 -35898
rect 26587 -36202 26623 -35898
rect 26927 -36202 26963 -35898
rect 27587 -36202 27623 -35898
rect 27927 -36202 27963 -35898
rect 28587 -36202 28623 -35898
rect 28927 -36202 28963 -35898
rect 29587 -36202 29623 -35898
rect 29927 -36202 29963 -35898
rect 30587 -36202 30623 -35898
rect 30927 -36202 30963 -35898
rect 31587 -36202 31623 -35898
rect 31927 -36202 31963 -35898
rect 32587 -36202 32623 -35898
rect 32927 -36202 32963 -35898
rect 33587 -36202 33623 -35898
rect 33927 -36202 33963 -35898
rect 34267 -36202 34275 -35898
rect 8275 -36210 34275 -36202
rect 8615 -36238 8935 -36210
rect 8615 -36862 8623 -36238
rect 8927 -36862 8935 -36238
rect 8615 -36890 8935 -36862
rect 9615 -36238 9935 -36210
rect 9615 -36862 9623 -36238
rect 9927 -36862 9935 -36238
rect 9615 -36890 9935 -36862
rect 10615 -36238 10935 -36210
rect 10615 -36862 10623 -36238
rect 10927 -36862 10935 -36238
rect 10615 -36890 10935 -36862
rect 11615 -36238 11935 -36210
rect 11615 -36862 11623 -36238
rect 11927 -36862 11935 -36238
rect 11615 -36890 11935 -36862
rect 12615 -36238 12935 -36210
rect 12615 -36862 12623 -36238
rect 12927 -36862 12935 -36238
rect 12615 -36890 12935 -36862
rect 13615 -36238 13935 -36210
rect 13615 -36862 13623 -36238
rect 13927 -36862 13935 -36238
rect 13615 -36890 13935 -36862
rect 14615 -36238 14935 -36210
rect 14615 -36862 14623 -36238
rect 14927 -36862 14935 -36238
rect 14615 -36890 14935 -36862
rect 15615 -36238 15935 -36210
rect 15615 -36862 15623 -36238
rect 15927 -36862 15935 -36238
rect 15615 -36890 15935 -36862
rect 16615 -36238 16935 -36210
rect 16615 -36862 16623 -36238
rect 16927 -36862 16935 -36238
rect 16615 -36890 16935 -36862
rect 17615 -36238 17935 -36210
rect 17615 -36862 17623 -36238
rect 17927 -36862 17935 -36238
rect 17615 -36890 17935 -36862
rect 18615 -36238 18935 -36210
rect 18615 -36862 18623 -36238
rect 18927 -36862 18935 -36238
rect 18615 -36890 18935 -36862
rect 19615 -36238 19935 -36210
rect 19615 -36862 19623 -36238
rect 19927 -36862 19935 -36238
rect 19615 -36890 19935 -36862
rect 20615 -36238 20935 -36210
rect 20615 -36862 20623 -36238
rect 20927 -36862 20935 -36238
rect 20615 -36890 20935 -36862
rect 21615 -36238 21935 -36210
rect 21615 -36862 21623 -36238
rect 21927 -36862 21935 -36238
rect 21615 -36890 21935 -36862
rect 22615 -36238 22935 -36210
rect 22615 -36862 22623 -36238
rect 22927 -36862 22935 -36238
rect 22615 -36890 22935 -36862
rect 23615 -36238 23935 -36210
rect 23615 -36862 23623 -36238
rect 23927 -36862 23935 -36238
rect 23615 -36890 23935 -36862
rect 24615 -36238 24935 -36210
rect 24615 -36862 24623 -36238
rect 24927 -36862 24935 -36238
rect 24615 -36890 24935 -36862
rect 25615 -36238 25935 -36210
rect 25615 -36862 25623 -36238
rect 25927 -36862 25935 -36238
rect 25615 -36890 25935 -36862
rect 26615 -36238 26935 -36210
rect 26615 -36862 26623 -36238
rect 26927 -36862 26935 -36238
rect 26615 -36890 26935 -36862
rect 27615 -36238 27935 -36210
rect 27615 -36862 27623 -36238
rect 27927 -36862 27935 -36238
rect 27615 -36890 27935 -36862
rect 28615 -36238 28935 -36210
rect 28615 -36862 28623 -36238
rect 28927 -36862 28935 -36238
rect 28615 -36890 28935 -36862
rect 29615 -36238 29935 -36210
rect 29615 -36862 29623 -36238
rect 29927 -36862 29935 -36238
rect 29615 -36890 29935 -36862
rect 30615 -36238 30935 -36210
rect 30615 -36862 30623 -36238
rect 30927 -36862 30935 -36238
rect 30615 -36890 30935 -36862
rect 31615 -36238 31935 -36210
rect 31615 -36862 31623 -36238
rect 31927 -36862 31935 -36238
rect 31615 -36890 31935 -36862
rect 32615 -36238 32935 -36210
rect 32615 -36862 32623 -36238
rect 32927 -36862 32935 -36238
rect 32615 -36890 32935 -36862
rect 33615 -36238 33935 -36210
rect 33615 -36862 33623 -36238
rect 33927 -36862 33935 -36238
rect 33615 -36890 33935 -36862
rect 8275 -36898 34275 -36890
rect 8275 -37202 8283 -36898
rect 8587 -37202 8623 -36898
rect 8927 -37202 8963 -36898
rect 9587 -37202 9623 -36898
rect 9927 -37202 9963 -36898
rect 10587 -37202 10623 -36898
rect 10927 -37202 10963 -36898
rect 11587 -37202 11623 -36898
rect 11927 -37202 11963 -36898
rect 12587 -37202 12623 -36898
rect 12927 -37202 12963 -36898
rect 13587 -37202 13623 -36898
rect 13927 -37202 13963 -36898
rect 14587 -37202 14623 -36898
rect 14927 -37202 14963 -36898
rect 15587 -37202 15623 -36898
rect 15927 -37202 15963 -36898
rect 16587 -37202 16623 -36898
rect 16927 -37202 16963 -36898
rect 17587 -37202 17623 -36898
rect 17927 -37202 17963 -36898
rect 18587 -37202 18623 -36898
rect 18927 -37202 18963 -36898
rect 19587 -37202 19623 -36898
rect 19927 -37202 19963 -36898
rect 20587 -37202 20623 -36898
rect 20927 -37202 20963 -36898
rect 21587 -37202 21623 -36898
rect 21927 -37202 21963 -36898
rect 22587 -37202 22623 -36898
rect 22927 -37202 22963 -36898
rect 23587 -37202 23623 -36898
rect 23927 -37202 23963 -36898
rect 24587 -37202 24623 -36898
rect 24927 -37202 24963 -36898
rect 25587 -37202 25623 -36898
rect 25927 -37202 25963 -36898
rect 26587 -37202 26623 -36898
rect 26927 -37202 26963 -36898
rect 27587 -37202 27623 -36898
rect 27927 -37202 27963 -36898
rect 28587 -37202 28623 -36898
rect 28927 -37202 28963 -36898
rect 29587 -37202 29623 -36898
rect 29927 -37202 29963 -36898
rect 30587 -37202 30623 -36898
rect 30927 -37202 30963 -36898
rect 31587 -37202 31623 -36898
rect 31927 -37202 31963 -36898
rect 32587 -37202 32623 -36898
rect 32927 -37202 32963 -36898
rect 33587 -37202 33623 -36898
rect 33927 -37202 33963 -36898
rect 34267 -37202 34275 -36898
rect 8275 -37210 34275 -37202
rect 8615 -37238 8935 -37210
rect 8615 -37862 8623 -37238
rect 8927 -37862 8935 -37238
rect 8615 -37890 8935 -37862
rect 9615 -37238 9935 -37210
rect 9615 -37862 9623 -37238
rect 9927 -37862 9935 -37238
rect 9615 -37890 9935 -37862
rect 10615 -37238 10935 -37210
rect 10615 -37862 10623 -37238
rect 10927 -37862 10935 -37238
rect 10615 -37890 10935 -37862
rect 11615 -37238 11935 -37210
rect 11615 -37862 11623 -37238
rect 11927 -37862 11935 -37238
rect 11615 -37890 11935 -37862
rect 12615 -37238 12935 -37210
rect 12615 -37862 12623 -37238
rect 12927 -37862 12935 -37238
rect 12615 -37890 12935 -37862
rect 13615 -37238 13935 -37210
rect 13615 -37862 13623 -37238
rect 13927 -37862 13935 -37238
rect 13615 -37890 13935 -37862
rect 14615 -37238 14935 -37210
rect 14615 -37862 14623 -37238
rect 14927 -37862 14935 -37238
rect 14615 -37890 14935 -37862
rect 15615 -37238 15935 -37210
rect 15615 -37862 15623 -37238
rect 15927 -37862 15935 -37238
rect 15615 -37890 15935 -37862
rect 16615 -37238 16935 -37210
rect 16615 -37862 16623 -37238
rect 16927 -37862 16935 -37238
rect 16615 -37890 16935 -37862
rect 17615 -37238 17935 -37210
rect 17615 -37862 17623 -37238
rect 17927 -37862 17935 -37238
rect 17615 -37890 17935 -37862
rect 18615 -37238 18935 -37210
rect 18615 -37862 18623 -37238
rect 18927 -37862 18935 -37238
rect 18615 -37890 18935 -37862
rect 19615 -37238 19935 -37210
rect 19615 -37862 19623 -37238
rect 19927 -37862 19935 -37238
rect 19615 -37890 19935 -37862
rect 20615 -37238 20935 -37210
rect 20615 -37862 20623 -37238
rect 20927 -37862 20935 -37238
rect 20615 -37890 20935 -37862
rect 21615 -37238 21935 -37210
rect 21615 -37862 21623 -37238
rect 21927 -37862 21935 -37238
rect 21615 -37890 21935 -37862
rect 22615 -37238 22935 -37210
rect 22615 -37862 22623 -37238
rect 22927 -37862 22935 -37238
rect 22615 -37890 22935 -37862
rect 23615 -37238 23935 -37210
rect 23615 -37862 23623 -37238
rect 23927 -37862 23935 -37238
rect 23615 -37890 23935 -37862
rect 24615 -37238 24935 -37210
rect 24615 -37862 24623 -37238
rect 24927 -37862 24935 -37238
rect 24615 -37890 24935 -37862
rect 25615 -37238 25935 -37210
rect 25615 -37862 25623 -37238
rect 25927 -37862 25935 -37238
rect 25615 -37890 25935 -37862
rect 26615 -37238 26935 -37210
rect 26615 -37862 26623 -37238
rect 26927 -37862 26935 -37238
rect 26615 -37890 26935 -37862
rect 27615 -37238 27935 -37210
rect 27615 -37862 27623 -37238
rect 27927 -37862 27935 -37238
rect 27615 -37890 27935 -37862
rect 28615 -37238 28935 -37210
rect 28615 -37862 28623 -37238
rect 28927 -37862 28935 -37238
rect 28615 -37890 28935 -37862
rect 29615 -37238 29935 -37210
rect 29615 -37862 29623 -37238
rect 29927 -37862 29935 -37238
rect 29615 -37890 29935 -37862
rect 30615 -37238 30935 -37210
rect 30615 -37862 30623 -37238
rect 30927 -37862 30935 -37238
rect 30615 -37890 30935 -37862
rect 31615 -37238 31935 -37210
rect 31615 -37862 31623 -37238
rect 31927 -37862 31935 -37238
rect 31615 -37890 31935 -37862
rect 32615 -37238 32935 -37210
rect 32615 -37862 32623 -37238
rect 32927 -37862 32935 -37238
rect 32615 -37890 32935 -37862
rect 33615 -37238 33935 -37210
rect 33615 -37862 33623 -37238
rect 33927 -37862 33935 -37238
rect 33615 -37890 33935 -37862
rect 8275 -37898 34275 -37890
rect 8275 -38202 8283 -37898
rect 8587 -38202 8623 -37898
rect 8927 -38202 8963 -37898
rect 9587 -38202 9623 -37898
rect 9927 -38202 9963 -37898
rect 10587 -38202 10623 -37898
rect 10927 -38202 10963 -37898
rect 11587 -38202 11623 -37898
rect 11927 -38202 11963 -37898
rect 12587 -38202 12623 -37898
rect 12927 -38202 12963 -37898
rect 13587 -38202 13623 -37898
rect 13927 -38202 13963 -37898
rect 14587 -38202 14623 -37898
rect 14927 -38202 14963 -37898
rect 15587 -38202 15623 -37898
rect 15927 -38202 15963 -37898
rect 16587 -38202 16623 -37898
rect 16927 -38202 16963 -37898
rect 17587 -38202 17623 -37898
rect 17927 -38202 17963 -37898
rect 18587 -38202 18623 -37898
rect 18927 -38202 18963 -37898
rect 19587 -38202 19623 -37898
rect 19927 -38202 19963 -37898
rect 20587 -38202 20623 -37898
rect 20927 -38202 20963 -37898
rect 21587 -38202 21623 -37898
rect 21927 -38202 21963 -37898
rect 22587 -38202 22623 -37898
rect 22927 -38202 22963 -37898
rect 23587 -38202 23623 -37898
rect 23927 -38202 23963 -37898
rect 24587 -38202 24623 -37898
rect 24927 -38202 24963 -37898
rect 25587 -38202 25623 -37898
rect 25927 -38202 25963 -37898
rect 26587 -38202 26623 -37898
rect 26927 -38202 26963 -37898
rect 27587 -38202 27623 -37898
rect 27927 -38202 27963 -37898
rect 28587 -38202 28623 -37898
rect 28927 -38202 28963 -37898
rect 29587 -38202 29623 -37898
rect 29927 -38202 29963 -37898
rect 30587 -38202 30623 -37898
rect 30927 -38202 30963 -37898
rect 31587 -38202 31623 -37898
rect 31927 -38202 31963 -37898
rect 32587 -38202 32623 -37898
rect 32927 -38202 32963 -37898
rect 33587 -38202 33623 -37898
rect 33927 -38202 33963 -37898
rect 34267 -38202 34275 -37898
rect 8275 -38210 34275 -38202
rect 8615 -38238 8935 -38210
rect 8615 -38862 8623 -38238
rect 8927 -38862 8935 -38238
rect 8615 -38890 8935 -38862
rect 9615 -38238 9935 -38210
rect 9615 -38862 9623 -38238
rect 9927 -38862 9935 -38238
rect 9615 -38890 9935 -38862
rect 10615 -38238 10935 -38210
rect 10615 -38862 10623 -38238
rect 10927 -38862 10935 -38238
rect 10615 -38890 10935 -38862
rect 11615 -38238 11935 -38210
rect 11615 -38862 11623 -38238
rect 11927 -38862 11935 -38238
rect 11615 -38890 11935 -38862
rect 12615 -38238 12935 -38210
rect 12615 -38862 12623 -38238
rect 12927 -38862 12935 -38238
rect 12615 -38890 12935 -38862
rect 13615 -38238 13935 -38210
rect 13615 -38862 13623 -38238
rect 13927 -38862 13935 -38238
rect 13615 -38890 13935 -38862
rect 14615 -38238 14935 -38210
rect 14615 -38862 14623 -38238
rect 14927 -38862 14935 -38238
rect 14615 -38890 14935 -38862
rect 15615 -38238 15935 -38210
rect 15615 -38862 15623 -38238
rect 15927 -38862 15935 -38238
rect 15615 -38890 15935 -38862
rect 16615 -38238 16935 -38210
rect 16615 -38862 16623 -38238
rect 16927 -38862 16935 -38238
rect 16615 -38890 16935 -38862
rect 17615 -38238 17935 -38210
rect 17615 -38862 17623 -38238
rect 17927 -38862 17935 -38238
rect 17615 -38890 17935 -38862
rect 18615 -38238 18935 -38210
rect 18615 -38862 18623 -38238
rect 18927 -38862 18935 -38238
rect 18615 -38890 18935 -38862
rect 19615 -38238 19935 -38210
rect 19615 -38862 19623 -38238
rect 19927 -38862 19935 -38238
rect 19615 -38890 19935 -38862
rect 20615 -38238 20935 -38210
rect 20615 -38862 20623 -38238
rect 20927 -38862 20935 -38238
rect 20615 -38890 20935 -38862
rect 21615 -38238 21935 -38210
rect 21615 -38862 21623 -38238
rect 21927 -38862 21935 -38238
rect 21615 -38890 21935 -38862
rect 22615 -38238 22935 -38210
rect 22615 -38862 22623 -38238
rect 22927 -38862 22935 -38238
rect 22615 -38890 22935 -38862
rect 23615 -38238 23935 -38210
rect 23615 -38862 23623 -38238
rect 23927 -38862 23935 -38238
rect 23615 -38890 23935 -38862
rect 24615 -38238 24935 -38210
rect 24615 -38862 24623 -38238
rect 24927 -38862 24935 -38238
rect 24615 -38890 24935 -38862
rect 25615 -38238 25935 -38210
rect 25615 -38862 25623 -38238
rect 25927 -38862 25935 -38238
rect 25615 -38890 25935 -38862
rect 26615 -38238 26935 -38210
rect 26615 -38862 26623 -38238
rect 26927 -38862 26935 -38238
rect 26615 -38890 26935 -38862
rect 27615 -38238 27935 -38210
rect 27615 -38862 27623 -38238
rect 27927 -38862 27935 -38238
rect 27615 -38890 27935 -38862
rect 28615 -38238 28935 -38210
rect 28615 -38862 28623 -38238
rect 28927 -38862 28935 -38238
rect 28615 -38890 28935 -38862
rect 29615 -38238 29935 -38210
rect 29615 -38862 29623 -38238
rect 29927 -38862 29935 -38238
rect 29615 -38890 29935 -38862
rect 30615 -38238 30935 -38210
rect 30615 -38862 30623 -38238
rect 30927 -38862 30935 -38238
rect 30615 -38890 30935 -38862
rect 31615 -38238 31935 -38210
rect 31615 -38862 31623 -38238
rect 31927 -38862 31935 -38238
rect 31615 -38890 31935 -38862
rect 32615 -38238 32935 -38210
rect 32615 -38862 32623 -38238
rect 32927 -38862 32935 -38238
rect 32615 -38890 32935 -38862
rect 33615 -38238 33935 -38210
rect 33615 -38862 33623 -38238
rect 33927 -38862 33935 -38238
rect 33615 -38890 33935 -38862
rect 8275 -38898 34275 -38890
rect 8275 -39202 8283 -38898
rect 8587 -39202 8623 -38898
rect 8927 -39202 8963 -38898
rect 9587 -39202 9623 -38898
rect 9927 -39202 9963 -38898
rect 10587 -39202 10623 -38898
rect 10927 -39202 10963 -38898
rect 11587 -39202 11623 -38898
rect 11927 -39202 11963 -38898
rect 12587 -39202 12623 -38898
rect 12927 -39202 12963 -38898
rect 13587 -39202 13623 -38898
rect 13927 -39202 13963 -38898
rect 14587 -39202 14623 -38898
rect 14927 -39202 14963 -38898
rect 15587 -39202 15623 -38898
rect 15927 -39202 15963 -38898
rect 16587 -39202 16623 -38898
rect 16927 -39202 16963 -38898
rect 17587 -39202 17623 -38898
rect 17927 -39202 17963 -38898
rect 18587 -39202 18623 -38898
rect 18927 -39202 18963 -38898
rect 19587 -39202 19623 -38898
rect 19927 -39202 19963 -38898
rect 20587 -39202 20623 -38898
rect 20927 -39202 20963 -38898
rect 21587 -39202 21623 -38898
rect 21927 -39202 21963 -38898
rect 22587 -39202 22623 -38898
rect 22927 -39202 22963 -38898
rect 23587 -39202 23623 -38898
rect 23927 -39202 23963 -38898
rect 24587 -39202 24623 -38898
rect 24927 -39202 24963 -38898
rect 25587 -39202 25623 -38898
rect 25927 -39202 25963 -38898
rect 26587 -39202 26623 -38898
rect 26927 -39202 26963 -38898
rect 27587 -39202 27623 -38898
rect 27927 -39202 27963 -38898
rect 28587 -39202 28623 -38898
rect 28927 -39202 28963 -38898
rect 29587 -39202 29623 -38898
rect 29927 -39202 29963 -38898
rect 30587 -39202 30623 -38898
rect 30927 -39202 30963 -38898
rect 31587 -39202 31623 -38898
rect 31927 -39202 31963 -38898
rect 32587 -39202 32623 -38898
rect 32927 -39202 32963 -38898
rect 33587 -39202 33623 -38898
rect 33927 -39202 33963 -38898
rect 34267 -39202 34275 -38898
rect 8275 -39210 34275 -39202
rect 8615 -39238 8935 -39210
rect 8615 -39862 8623 -39238
rect 8927 -39862 8935 -39238
rect 8615 -39890 8935 -39862
rect 9615 -39238 9935 -39210
rect 9615 -39862 9623 -39238
rect 9927 -39862 9935 -39238
rect 9615 -39890 9935 -39862
rect 10615 -39238 10935 -39210
rect 10615 -39862 10623 -39238
rect 10927 -39862 10935 -39238
rect 10615 -39890 10935 -39862
rect 11615 -39238 11935 -39210
rect 11615 -39862 11623 -39238
rect 11927 -39862 11935 -39238
rect 11615 -39890 11935 -39862
rect 12615 -39238 12935 -39210
rect 12615 -39862 12623 -39238
rect 12927 -39862 12935 -39238
rect 12615 -39890 12935 -39862
rect 13615 -39238 13935 -39210
rect 13615 -39862 13623 -39238
rect 13927 -39862 13935 -39238
rect 13615 -39890 13935 -39862
rect 14615 -39238 14935 -39210
rect 14615 -39862 14623 -39238
rect 14927 -39862 14935 -39238
rect 14615 -39890 14935 -39862
rect 15615 -39238 15935 -39210
rect 15615 -39862 15623 -39238
rect 15927 -39862 15935 -39238
rect 15615 -39890 15935 -39862
rect 16615 -39238 16935 -39210
rect 16615 -39862 16623 -39238
rect 16927 -39862 16935 -39238
rect 16615 -39890 16935 -39862
rect 17615 -39238 17935 -39210
rect 17615 -39862 17623 -39238
rect 17927 -39862 17935 -39238
rect 17615 -39890 17935 -39862
rect 18615 -39238 18935 -39210
rect 18615 -39862 18623 -39238
rect 18927 -39862 18935 -39238
rect 18615 -39890 18935 -39862
rect 19615 -39238 19935 -39210
rect 19615 -39862 19623 -39238
rect 19927 -39862 19935 -39238
rect 19615 -39890 19935 -39862
rect 20615 -39238 20935 -39210
rect 20615 -39862 20623 -39238
rect 20927 -39862 20935 -39238
rect 20615 -39890 20935 -39862
rect 21615 -39238 21935 -39210
rect 21615 -39862 21623 -39238
rect 21927 -39862 21935 -39238
rect 21615 -39890 21935 -39862
rect 22615 -39238 22935 -39210
rect 22615 -39862 22623 -39238
rect 22927 -39862 22935 -39238
rect 22615 -39890 22935 -39862
rect 23615 -39238 23935 -39210
rect 23615 -39862 23623 -39238
rect 23927 -39862 23935 -39238
rect 23615 -39890 23935 -39862
rect 24615 -39238 24935 -39210
rect 24615 -39862 24623 -39238
rect 24927 -39862 24935 -39238
rect 24615 -39890 24935 -39862
rect 25615 -39238 25935 -39210
rect 25615 -39862 25623 -39238
rect 25927 -39862 25935 -39238
rect 25615 -39890 25935 -39862
rect 26615 -39238 26935 -39210
rect 26615 -39862 26623 -39238
rect 26927 -39862 26935 -39238
rect 26615 -39890 26935 -39862
rect 27615 -39238 27935 -39210
rect 27615 -39862 27623 -39238
rect 27927 -39862 27935 -39238
rect 27615 -39890 27935 -39862
rect 28615 -39238 28935 -39210
rect 28615 -39862 28623 -39238
rect 28927 -39862 28935 -39238
rect 28615 -39890 28935 -39862
rect 29615 -39238 29935 -39210
rect 29615 -39862 29623 -39238
rect 29927 -39862 29935 -39238
rect 29615 -39890 29935 -39862
rect 30615 -39238 30935 -39210
rect 30615 -39862 30623 -39238
rect 30927 -39862 30935 -39238
rect 30615 -39890 30935 -39862
rect 31615 -39238 31935 -39210
rect 31615 -39862 31623 -39238
rect 31927 -39862 31935 -39238
rect 31615 -39890 31935 -39862
rect 32615 -39238 32935 -39210
rect 32615 -39862 32623 -39238
rect 32927 -39862 32935 -39238
rect 32615 -39890 32935 -39862
rect 33615 -39238 33935 -39210
rect 33615 -39862 33623 -39238
rect 33927 -39862 33935 -39238
rect 33615 -39890 33935 -39862
rect 8275 -39898 34275 -39890
rect 8275 -40202 8283 -39898
rect 8587 -40202 8623 -39898
rect 8927 -40202 8963 -39898
rect 9587 -40202 9623 -39898
rect 9927 -40202 9963 -39898
rect 10587 -40202 10623 -39898
rect 10927 -40202 10963 -39898
rect 11587 -40202 11623 -39898
rect 11927 -40202 11963 -39898
rect 12587 -40202 12623 -39898
rect 12927 -40202 12963 -39898
rect 13587 -40202 13623 -39898
rect 13927 -40202 13963 -39898
rect 14587 -40202 14623 -39898
rect 14927 -40202 14963 -39898
rect 15587 -40202 15623 -39898
rect 15927 -40202 15963 -39898
rect 16587 -40202 16623 -39898
rect 16927 -40202 16963 -39898
rect 17587 -40202 17623 -39898
rect 17927 -40202 17963 -39898
rect 18587 -40202 18623 -39898
rect 18927 -40202 18963 -39898
rect 19587 -40202 19623 -39898
rect 19927 -40202 19963 -39898
rect 20587 -40202 20623 -39898
rect 20927 -40202 20963 -39898
rect 21587 -40202 21623 -39898
rect 21927 -40202 21963 -39898
rect 22587 -40202 22623 -39898
rect 22927 -40202 22963 -39898
rect 23587 -40202 23623 -39898
rect 23927 -40202 23963 -39898
rect 24587 -40202 24623 -39898
rect 24927 -40202 24963 -39898
rect 25587 -40202 25623 -39898
rect 25927 -40202 25963 -39898
rect 26587 -40202 26623 -39898
rect 26927 -40202 26963 -39898
rect 27587 -40202 27623 -39898
rect 27927 -40202 27963 -39898
rect 28587 -40202 28623 -39898
rect 28927 -40202 28963 -39898
rect 29587 -40202 29623 -39898
rect 29927 -40202 29963 -39898
rect 30587 -40202 30623 -39898
rect 30927 -40202 30963 -39898
rect 31587 -40202 31623 -39898
rect 31927 -40202 31963 -39898
rect 32587 -40202 32623 -39898
rect 32927 -40202 32963 -39898
rect 33587 -40202 33623 -39898
rect 33927 -40202 33963 -39898
rect 34267 -40202 34275 -39898
rect 8275 -40210 34275 -40202
rect 8615 -40238 8935 -40210
rect 8615 -40862 8623 -40238
rect 8927 -40862 8935 -40238
rect 8615 -40890 8935 -40862
rect 9615 -40238 9935 -40210
rect 9615 -40862 9623 -40238
rect 9927 -40862 9935 -40238
rect 9615 -40890 9935 -40862
rect 10615 -40238 10935 -40210
rect 10615 -40862 10623 -40238
rect 10927 -40862 10935 -40238
rect 10615 -40890 10935 -40862
rect 11615 -40238 11935 -40210
rect 11615 -40862 11623 -40238
rect 11927 -40862 11935 -40238
rect 11615 -40890 11935 -40862
rect 12615 -40238 12935 -40210
rect 12615 -40862 12623 -40238
rect 12927 -40862 12935 -40238
rect 12615 -40890 12935 -40862
rect 13615 -40238 13935 -40210
rect 13615 -40862 13623 -40238
rect 13927 -40862 13935 -40238
rect 13615 -40890 13935 -40862
rect 14615 -40238 14935 -40210
rect 14615 -40862 14623 -40238
rect 14927 -40862 14935 -40238
rect 14615 -40890 14935 -40862
rect 15615 -40238 15935 -40210
rect 15615 -40862 15623 -40238
rect 15927 -40862 15935 -40238
rect 15615 -40890 15935 -40862
rect 16615 -40238 16935 -40210
rect 16615 -40862 16623 -40238
rect 16927 -40862 16935 -40238
rect 16615 -40890 16935 -40862
rect 17615 -40238 17935 -40210
rect 17615 -40862 17623 -40238
rect 17927 -40862 17935 -40238
rect 17615 -40890 17935 -40862
rect 18615 -40238 18935 -40210
rect 18615 -40862 18623 -40238
rect 18927 -40862 18935 -40238
rect 18615 -40890 18935 -40862
rect 19615 -40238 19935 -40210
rect 19615 -40862 19623 -40238
rect 19927 -40862 19935 -40238
rect 19615 -40890 19935 -40862
rect 20615 -40238 20935 -40210
rect 20615 -40862 20623 -40238
rect 20927 -40862 20935 -40238
rect 20615 -40890 20935 -40862
rect 21615 -40238 21935 -40210
rect 21615 -40862 21623 -40238
rect 21927 -40862 21935 -40238
rect 21615 -40890 21935 -40862
rect 22615 -40238 22935 -40210
rect 22615 -40862 22623 -40238
rect 22927 -40862 22935 -40238
rect 22615 -40890 22935 -40862
rect 23615 -40238 23935 -40210
rect 23615 -40862 23623 -40238
rect 23927 -40862 23935 -40238
rect 23615 -40890 23935 -40862
rect 24615 -40238 24935 -40210
rect 24615 -40862 24623 -40238
rect 24927 -40862 24935 -40238
rect 24615 -40890 24935 -40862
rect 25615 -40238 25935 -40210
rect 25615 -40862 25623 -40238
rect 25927 -40862 25935 -40238
rect 25615 -40890 25935 -40862
rect 26615 -40238 26935 -40210
rect 26615 -40862 26623 -40238
rect 26927 -40862 26935 -40238
rect 26615 -40890 26935 -40862
rect 27615 -40238 27935 -40210
rect 27615 -40862 27623 -40238
rect 27927 -40862 27935 -40238
rect 27615 -40890 27935 -40862
rect 28615 -40238 28935 -40210
rect 28615 -40862 28623 -40238
rect 28927 -40862 28935 -40238
rect 28615 -40890 28935 -40862
rect 29615 -40238 29935 -40210
rect 29615 -40862 29623 -40238
rect 29927 -40862 29935 -40238
rect 29615 -40890 29935 -40862
rect 30615 -40238 30935 -40210
rect 30615 -40862 30623 -40238
rect 30927 -40862 30935 -40238
rect 30615 -40890 30935 -40862
rect 31615 -40238 31935 -40210
rect 31615 -40862 31623 -40238
rect 31927 -40862 31935 -40238
rect 31615 -40890 31935 -40862
rect 32615 -40238 32935 -40210
rect 32615 -40862 32623 -40238
rect 32927 -40862 32935 -40238
rect 32615 -40890 32935 -40862
rect 33615 -40238 33935 -40210
rect 33615 -40862 33623 -40238
rect 33927 -40862 33935 -40238
rect 33615 -40890 33935 -40862
rect 8275 -40898 34275 -40890
rect 8275 -41202 8283 -40898
rect 8587 -41202 8623 -40898
rect 8927 -41202 8963 -40898
rect 9587 -41202 9623 -40898
rect 9927 -41202 9963 -40898
rect 10587 -41202 10623 -40898
rect 10927 -41202 10963 -40898
rect 11587 -41202 11623 -40898
rect 11927 -41202 11963 -40898
rect 12587 -41202 12623 -40898
rect 12927 -41202 12963 -40898
rect 13587 -41202 13623 -40898
rect 13927 -41202 13963 -40898
rect 14587 -41202 14623 -40898
rect 14927 -41202 14963 -40898
rect 15587 -41202 15623 -40898
rect 15927 -41202 15963 -40898
rect 16587 -41202 16623 -40898
rect 16927 -41202 16963 -40898
rect 17587 -41202 17623 -40898
rect 17927 -41202 17963 -40898
rect 18587 -41202 18623 -40898
rect 18927 -41202 18963 -40898
rect 19587 -41202 19623 -40898
rect 19927 -41202 19963 -40898
rect 20587 -41202 20623 -40898
rect 20927 -41202 20963 -40898
rect 21587 -41202 21623 -40898
rect 21927 -41202 21963 -40898
rect 22587 -41202 22623 -40898
rect 22927 -41202 22963 -40898
rect 23587 -41202 23623 -40898
rect 23927 -41202 23963 -40898
rect 24587 -41202 24623 -40898
rect 24927 -41202 24963 -40898
rect 25587 -41202 25623 -40898
rect 25927 -41202 25963 -40898
rect 26587 -41202 26623 -40898
rect 26927 -41202 26963 -40898
rect 27587 -41202 27623 -40898
rect 27927 -41202 27963 -40898
rect 28587 -41202 28623 -40898
rect 28927 -41202 28963 -40898
rect 29587 -41202 29623 -40898
rect 29927 -41202 29963 -40898
rect 30587 -41202 30623 -40898
rect 30927 -41202 30963 -40898
rect 31587 -41202 31623 -40898
rect 31927 -41202 31963 -40898
rect 32587 -41202 32623 -40898
rect 32927 -41202 32963 -40898
rect 33587 -41202 33623 -40898
rect 33927 -41202 33963 -40898
rect 34267 -41202 34275 -40898
rect 8275 -41210 34275 -41202
rect 8615 -41238 8935 -41210
rect 8615 -41862 8623 -41238
rect 8927 -41862 8935 -41238
rect 8615 -41890 8935 -41862
rect 9615 -41238 9935 -41210
rect 9615 -41862 9623 -41238
rect 9927 -41862 9935 -41238
rect 9615 -41890 9935 -41862
rect 10615 -41238 10935 -41210
rect 10615 -41862 10623 -41238
rect 10927 -41862 10935 -41238
rect 10615 -41890 10935 -41862
rect 11615 -41238 11935 -41210
rect 11615 -41862 11623 -41238
rect 11927 -41862 11935 -41238
rect 11615 -41890 11935 -41862
rect 12615 -41238 12935 -41210
rect 12615 -41862 12623 -41238
rect 12927 -41862 12935 -41238
rect 12615 -41890 12935 -41862
rect 13615 -41238 13935 -41210
rect 13615 -41862 13623 -41238
rect 13927 -41862 13935 -41238
rect 13615 -41890 13935 -41862
rect 14615 -41238 14935 -41210
rect 14615 -41862 14623 -41238
rect 14927 -41862 14935 -41238
rect 14615 -41890 14935 -41862
rect 15615 -41238 15935 -41210
rect 15615 -41862 15623 -41238
rect 15927 -41862 15935 -41238
rect 15615 -41890 15935 -41862
rect 16615 -41238 16935 -41210
rect 16615 -41862 16623 -41238
rect 16927 -41862 16935 -41238
rect 16615 -41890 16935 -41862
rect 17615 -41238 17935 -41210
rect 17615 -41862 17623 -41238
rect 17927 -41862 17935 -41238
rect 17615 -41890 17935 -41862
rect 18615 -41238 18935 -41210
rect 18615 -41862 18623 -41238
rect 18927 -41862 18935 -41238
rect 18615 -41890 18935 -41862
rect 19615 -41238 19935 -41210
rect 19615 -41862 19623 -41238
rect 19927 -41862 19935 -41238
rect 19615 -41890 19935 -41862
rect 20615 -41238 20935 -41210
rect 20615 -41862 20623 -41238
rect 20927 -41862 20935 -41238
rect 20615 -41890 20935 -41862
rect 21615 -41238 21935 -41210
rect 21615 -41862 21623 -41238
rect 21927 -41862 21935 -41238
rect 21615 -41890 21935 -41862
rect 22615 -41238 22935 -41210
rect 22615 -41862 22623 -41238
rect 22927 -41862 22935 -41238
rect 22615 -41890 22935 -41862
rect 23615 -41238 23935 -41210
rect 23615 -41862 23623 -41238
rect 23927 -41862 23935 -41238
rect 23615 -41890 23935 -41862
rect 24615 -41238 24935 -41210
rect 24615 -41862 24623 -41238
rect 24927 -41862 24935 -41238
rect 24615 -41890 24935 -41862
rect 25615 -41238 25935 -41210
rect 25615 -41862 25623 -41238
rect 25927 -41862 25935 -41238
rect 25615 -41890 25935 -41862
rect 26615 -41238 26935 -41210
rect 26615 -41862 26623 -41238
rect 26927 -41862 26935 -41238
rect 26615 -41890 26935 -41862
rect 27615 -41238 27935 -41210
rect 27615 -41862 27623 -41238
rect 27927 -41862 27935 -41238
rect 27615 -41890 27935 -41862
rect 28615 -41238 28935 -41210
rect 28615 -41862 28623 -41238
rect 28927 -41862 28935 -41238
rect 28615 -41890 28935 -41862
rect 29615 -41238 29935 -41210
rect 29615 -41862 29623 -41238
rect 29927 -41862 29935 -41238
rect 29615 -41890 29935 -41862
rect 30615 -41238 30935 -41210
rect 30615 -41862 30623 -41238
rect 30927 -41862 30935 -41238
rect 30615 -41890 30935 -41862
rect 31615 -41238 31935 -41210
rect 31615 -41862 31623 -41238
rect 31927 -41862 31935 -41238
rect 31615 -41890 31935 -41862
rect 32615 -41238 32935 -41210
rect 32615 -41862 32623 -41238
rect 32927 -41862 32935 -41238
rect 32615 -41890 32935 -41862
rect 33615 -41238 33935 -41210
rect 33615 -41862 33623 -41238
rect 33927 -41862 33935 -41238
rect 33615 -41890 33935 -41862
rect 8275 -41898 34275 -41890
rect 8275 -42202 8283 -41898
rect 8587 -42202 8623 -41898
rect 8927 -42202 8963 -41898
rect 9587 -42202 9623 -41898
rect 9927 -42202 9963 -41898
rect 10587 -42202 10623 -41898
rect 10927 -42202 10963 -41898
rect 11587 -42202 11623 -41898
rect 11927 -42202 11963 -41898
rect 12587 -42202 12623 -41898
rect 12927 -42202 12963 -41898
rect 13587 -42202 13623 -41898
rect 13927 -42202 13963 -41898
rect 14587 -42202 14623 -41898
rect 14927 -42202 14963 -41898
rect 15587 -42202 15623 -41898
rect 15927 -42202 15963 -41898
rect 16587 -42202 16623 -41898
rect 16927 -42202 16963 -41898
rect 17587 -42202 17623 -41898
rect 17927 -42202 17963 -41898
rect 18587 -42202 18623 -41898
rect 18927 -42202 18963 -41898
rect 19587 -42202 19623 -41898
rect 19927 -42202 19963 -41898
rect 20587 -42202 20623 -41898
rect 20927 -42202 20963 -41898
rect 21587 -42202 21623 -41898
rect 21927 -42202 21963 -41898
rect 22587 -42202 22623 -41898
rect 22927 -42202 22963 -41898
rect 23587 -42202 23623 -41898
rect 23927 -42202 23963 -41898
rect 24587 -42202 24623 -41898
rect 24927 -42202 24963 -41898
rect 25587 -42202 25623 -41898
rect 25927 -42202 25963 -41898
rect 26587 -42202 26623 -41898
rect 26927 -42202 26963 -41898
rect 27587 -42202 27623 -41898
rect 27927 -42202 27963 -41898
rect 28587 -42202 28623 -41898
rect 28927 -42202 28963 -41898
rect 29587 -42202 29623 -41898
rect 29927 -42202 29963 -41898
rect 30587 -42202 30623 -41898
rect 30927 -42202 30963 -41898
rect 31587 -42202 31623 -41898
rect 31927 -42202 31963 -41898
rect 32587 -42202 32623 -41898
rect 32927 -42202 32963 -41898
rect 33587 -42202 33623 -41898
rect 33927 -42202 33963 -41898
rect 34267 -42202 34275 -41898
rect 8275 -42210 34275 -42202
rect 8615 -42238 8935 -42210
rect 8615 -42862 8623 -42238
rect 8927 -42862 8935 -42238
rect 8615 -42890 8935 -42862
rect 9615 -42238 9935 -42210
rect 9615 -42862 9623 -42238
rect 9927 -42862 9935 -42238
rect 9615 -42890 9935 -42862
rect 10615 -42238 10935 -42210
rect 10615 -42862 10623 -42238
rect 10927 -42862 10935 -42238
rect 10615 -42890 10935 -42862
rect 11615 -42238 11935 -42210
rect 11615 -42862 11623 -42238
rect 11927 -42862 11935 -42238
rect 11615 -42890 11935 -42862
rect 12615 -42238 12935 -42210
rect 12615 -42862 12623 -42238
rect 12927 -42862 12935 -42238
rect 12615 -42890 12935 -42862
rect 13615 -42238 13935 -42210
rect 13615 -42862 13623 -42238
rect 13927 -42862 13935 -42238
rect 13615 -42890 13935 -42862
rect 14615 -42238 14935 -42210
rect 14615 -42862 14623 -42238
rect 14927 -42862 14935 -42238
rect 14615 -42890 14935 -42862
rect 15615 -42238 15935 -42210
rect 15615 -42862 15623 -42238
rect 15927 -42862 15935 -42238
rect 15615 -42890 15935 -42862
rect 16615 -42238 16935 -42210
rect 16615 -42862 16623 -42238
rect 16927 -42862 16935 -42238
rect 16615 -42890 16935 -42862
rect 17615 -42238 17935 -42210
rect 17615 -42862 17623 -42238
rect 17927 -42862 17935 -42238
rect 17615 -42890 17935 -42862
rect 18615 -42238 18935 -42210
rect 18615 -42862 18623 -42238
rect 18927 -42862 18935 -42238
rect 18615 -42890 18935 -42862
rect 19615 -42238 19935 -42210
rect 19615 -42862 19623 -42238
rect 19927 -42862 19935 -42238
rect 19615 -42890 19935 -42862
rect 20615 -42238 20935 -42210
rect 20615 -42862 20623 -42238
rect 20927 -42862 20935 -42238
rect 20615 -42890 20935 -42862
rect 21615 -42238 21935 -42210
rect 21615 -42862 21623 -42238
rect 21927 -42862 21935 -42238
rect 21615 -42890 21935 -42862
rect 22615 -42238 22935 -42210
rect 22615 -42862 22623 -42238
rect 22927 -42862 22935 -42238
rect 22615 -42890 22935 -42862
rect 23615 -42238 23935 -42210
rect 23615 -42862 23623 -42238
rect 23927 -42862 23935 -42238
rect 23615 -42890 23935 -42862
rect 24615 -42238 24935 -42210
rect 24615 -42862 24623 -42238
rect 24927 -42862 24935 -42238
rect 24615 -42890 24935 -42862
rect 25615 -42238 25935 -42210
rect 25615 -42862 25623 -42238
rect 25927 -42862 25935 -42238
rect 25615 -42890 25935 -42862
rect 26615 -42238 26935 -42210
rect 26615 -42862 26623 -42238
rect 26927 -42862 26935 -42238
rect 26615 -42890 26935 -42862
rect 27615 -42238 27935 -42210
rect 27615 -42862 27623 -42238
rect 27927 -42862 27935 -42238
rect 27615 -42890 27935 -42862
rect 28615 -42238 28935 -42210
rect 28615 -42862 28623 -42238
rect 28927 -42862 28935 -42238
rect 28615 -42890 28935 -42862
rect 29615 -42238 29935 -42210
rect 29615 -42862 29623 -42238
rect 29927 -42862 29935 -42238
rect 29615 -42890 29935 -42862
rect 30615 -42238 30935 -42210
rect 30615 -42862 30623 -42238
rect 30927 -42862 30935 -42238
rect 30615 -42890 30935 -42862
rect 31615 -42238 31935 -42210
rect 31615 -42862 31623 -42238
rect 31927 -42862 31935 -42238
rect 31615 -42890 31935 -42862
rect 32615 -42238 32935 -42210
rect 32615 -42862 32623 -42238
rect 32927 -42862 32935 -42238
rect 32615 -42890 32935 -42862
rect 33615 -42238 33935 -42210
rect 33615 -42862 33623 -42238
rect 33927 -42862 33935 -42238
rect 33615 -42890 33935 -42862
rect 8275 -42898 34275 -42890
rect 8275 -43202 8283 -42898
rect 8587 -43202 8623 -42898
rect 8927 -43202 8963 -42898
rect 9587 -43202 9623 -42898
rect 9927 -43202 9963 -42898
rect 10587 -43202 10623 -42898
rect 10927 -43202 10963 -42898
rect 11587 -43202 11623 -42898
rect 11927 -43202 11963 -42898
rect 12587 -43202 12623 -42898
rect 12927 -43202 12963 -42898
rect 13587 -43202 13623 -42898
rect 13927 -43202 13963 -42898
rect 14587 -43202 14623 -42898
rect 14927 -43202 14963 -42898
rect 15587 -43202 15623 -42898
rect 15927 -43202 15963 -42898
rect 16587 -43202 16623 -42898
rect 16927 -43202 16963 -42898
rect 17587 -43202 17623 -42898
rect 17927 -43202 17963 -42898
rect 18587 -43202 18623 -42898
rect 18927 -43202 18963 -42898
rect 19587 -43202 19623 -42898
rect 19927 -43202 19963 -42898
rect 20587 -43202 20623 -42898
rect 20927 -43202 20963 -42898
rect 21587 -43202 21623 -42898
rect 21927 -43202 21963 -42898
rect 22587 -43202 22623 -42898
rect 22927 -43202 22963 -42898
rect 23587 -43202 23623 -42898
rect 23927 -43202 23963 -42898
rect 24587 -43202 24623 -42898
rect 24927 -43202 24963 -42898
rect 25587 -43202 25623 -42898
rect 25927 -43202 25963 -42898
rect 26587 -43202 26623 -42898
rect 26927 -43202 26963 -42898
rect 27587 -43202 27623 -42898
rect 27927 -43202 27963 -42898
rect 28587 -43202 28623 -42898
rect 28927 -43202 28963 -42898
rect 29587 -43202 29623 -42898
rect 29927 -43202 29963 -42898
rect 30587 -43202 30623 -42898
rect 30927 -43202 30963 -42898
rect 31587 -43202 31623 -42898
rect 31927 -43202 31963 -42898
rect 32587 -43202 32623 -42898
rect 32927 -43202 32963 -42898
rect 33587 -43202 33623 -42898
rect 33927 -43202 33963 -42898
rect 34267 -43202 34275 -42898
rect 8275 -43210 34275 -43202
rect 8615 -43238 8935 -43210
rect 8615 -43862 8623 -43238
rect 8927 -43862 8935 -43238
rect 8615 -43890 8935 -43862
rect 9615 -43238 9935 -43210
rect 9615 -43862 9623 -43238
rect 9927 -43862 9935 -43238
rect 9615 -43890 9935 -43862
rect 10615 -43238 10935 -43210
rect 10615 -43862 10623 -43238
rect 10927 -43862 10935 -43238
rect 10615 -43890 10935 -43862
rect 11615 -43238 11935 -43210
rect 11615 -43862 11623 -43238
rect 11927 -43862 11935 -43238
rect 11615 -43890 11935 -43862
rect 12615 -43238 12935 -43210
rect 12615 -43862 12623 -43238
rect 12927 -43862 12935 -43238
rect 12615 -43890 12935 -43862
rect 13615 -43238 13935 -43210
rect 13615 -43862 13623 -43238
rect 13927 -43862 13935 -43238
rect 13615 -43890 13935 -43862
rect 14615 -43238 14935 -43210
rect 14615 -43862 14623 -43238
rect 14927 -43862 14935 -43238
rect 14615 -43890 14935 -43862
rect 15615 -43238 15935 -43210
rect 15615 -43862 15623 -43238
rect 15927 -43862 15935 -43238
rect 15615 -43890 15935 -43862
rect 16615 -43238 16935 -43210
rect 16615 -43862 16623 -43238
rect 16927 -43862 16935 -43238
rect 16615 -43890 16935 -43862
rect 17615 -43238 17935 -43210
rect 17615 -43862 17623 -43238
rect 17927 -43862 17935 -43238
rect 17615 -43890 17935 -43862
rect 18615 -43238 18935 -43210
rect 18615 -43862 18623 -43238
rect 18927 -43862 18935 -43238
rect 18615 -43890 18935 -43862
rect 19615 -43238 19935 -43210
rect 19615 -43862 19623 -43238
rect 19927 -43862 19935 -43238
rect 19615 -43890 19935 -43862
rect 20615 -43238 20935 -43210
rect 20615 -43862 20623 -43238
rect 20927 -43862 20935 -43238
rect 20615 -43890 20935 -43862
rect 21615 -43238 21935 -43210
rect 21615 -43862 21623 -43238
rect 21927 -43862 21935 -43238
rect 21615 -43890 21935 -43862
rect 22615 -43238 22935 -43210
rect 22615 -43862 22623 -43238
rect 22927 -43862 22935 -43238
rect 22615 -43890 22935 -43862
rect 23615 -43238 23935 -43210
rect 23615 -43862 23623 -43238
rect 23927 -43862 23935 -43238
rect 23615 -43890 23935 -43862
rect 24615 -43238 24935 -43210
rect 24615 -43862 24623 -43238
rect 24927 -43862 24935 -43238
rect 24615 -43890 24935 -43862
rect 25615 -43238 25935 -43210
rect 25615 -43862 25623 -43238
rect 25927 -43862 25935 -43238
rect 25615 -43890 25935 -43862
rect 26615 -43238 26935 -43210
rect 26615 -43862 26623 -43238
rect 26927 -43862 26935 -43238
rect 26615 -43890 26935 -43862
rect 27615 -43238 27935 -43210
rect 27615 -43862 27623 -43238
rect 27927 -43862 27935 -43238
rect 27615 -43890 27935 -43862
rect 28615 -43238 28935 -43210
rect 28615 -43862 28623 -43238
rect 28927 -43862 28935 -43238
rect 28615 -43890 28935 -43862
rect 29615 -43238 29935 -43210
rect 29615 -43862 29623 -43238
rect 29927 -43862 29935 -43238
rect 29615 -43890 29935 -43862
rect 30615 -43238 30935 -43210
rect 30615 -43862 30623 -43238
rect 30927 -43862 30935 -43238
rect 30615 -43890 30935 -43862
rect 31615 -43238 31935 -43210
rect 31615 -43862 31623 -43238
rect 31927 -43862 31935 -43238
rect 31615 -43890 31935 -43862
rect 32615 -43238 32935 -43210
rect 32615 -43862 32623 -43238
rect 32927 -43862 32935 -43238
rect 32615 -43890 32935 -43862
rect 33615 -43238 33935 -43210
rect 33615 -43862 33623 -43238
rect 33927 -43862 33935 -43238
rect 33615 -43890 33935 -43862
rect 8275 -43898 34275 -43890
rect 8275 -44202 8283 -43898
rect 8587 -44202 8623 -43898
rect 8927 -44202 8963 -43898
rect 9587 -44202 9623 -43898
rect 9927 -44202 9963 -43898
rect 10587 -44202 10623 -43898
rect 10927 -44202 10963 -43898
rect 11587 -44202 11623 -43898
rect 11927 -44202 11963 -43898
rect 12587 -44202 12623 -43898
rect 12927 -44202 12963 -43898
rect 13587 -44202 13623 -43898
rect 13927 -44202 13963 -43898
rect 14587 -44202 14623 -43898
rect 14927 -44202 14963 -43898
rect 15587 -44202 15623 -43898
rect 15927 -44202 15963 -43898
rect 16587 -44202 16623 -43898
rect 16927 -44202 16963 -43898
rect 17587 -44202 17623 -43898
rect 17927 -44202 17963 -43898
rect 18587 -44202 18623 -43898
rect 18927 -44202 18963 -43898
rect 19587 -44202 19623 -43898
rect 19927 -44202 19963 -43898
rect 20587 -44202 20623 -43898
rect 20927 -44202 20963 -43898
rect 21587 -44202 21623 -43898
rect 21927 -44202 21963 -43898
rect 22587 -44202 22623 -43898
rect 22927 -44202 22963 -43898
rect 23587 -44202 23623 -43898
rect 23927 -44202 23963 -43898
rect 24587 -44202 24623 -43898
rect 24927 -44202 24963 -43898
rect 25587 -44202 25623 -43898
rect 25927 -44202 25963 -43898
rect 26587 -44202 26623 -43898
rect 26927 -44202 26963 -43898
rect 27587 -44202 27623 -43898
rect 27927 -44202 27963 -43898
rect 28587 -44202 28623 -43898
rect 28927 -44202 28963 -43898
rect 29587 -44202 29623 -43898
rect 29927 -44202 29963 -43898
rect 30587 -44202 30623 -43898
rect 30927 -44202 30963 -43898
rect 31587 -44202 31623 -43898
rect 31927 -44202 31963 -43898
rect 32587 -44202 32623 -43898
rect 32927 -44202 32963 -43898
rect 33587 -44202 33623 -43898
rect 33927 -44202 33963 -43898
rect 34267 -44202 34275 -43898
rect 8275 -44210 34275 -44202
rect -4275 -44550 5725 -44502
rect 8615 -44238 8935 -44210
rect -49485 -44890 -49165 -44862
rect 8615 -44862 8623 -44238
rect 8927 -44862 8935 -44238
rect 8615 -44890 8935 -44862
rect 9615 -44238 9935 -44210
rect 9615 -44862 9623 -44238
rect 9927 -44862 9935 -44238
rect 9615 -44890 9935 -44862
rect 10615 -44238 10935 -44210
rect 10615 -44862 10623 -44238
rect 10927 -44862 10935 -44238
rect 10615 -44890 10935 -44862
rect 11615 -44238 11935 -44210
rect 11615 -44862 11623 -44238
rect 11927 -44862 11935 -44238
rect 11615 -44890 11935 -44862
rect 12615 -44238 12935 -44210
rect 12615 -44862 12623 -44238
rect 12927 -44862 12935 -44238
rect 12615 -44890 12935 -44862
rect 13615 -44238 13935 -44210
rect 13615 -44862 13623 -44238
rect 13927 -44862 13935 -44238
rect 13615 -44890 13935 -44862
rect 14615 -44238 14935 -44210
rect 14615 -44862 14623 -44238
rect 14927 -44862 14935 -44238
rect 14615 -44890 14935 -44862
rect 15615 -44238 15935 -44210
rect 15615 -44862 15623 -44238
rect 15927 -44862 15935 -44238
rect 15615 -44890 15935 -44862
rect 16615 -44238 16935 -44210
rect 16615 -44862 16623 -44238
rect 16927 -44862 16935 -44238
rect 16615 -44890 16935 -44862
rect 17615 -44238 17935 -44210
rect 17615 -44862 17623 -44238
rect 17927 -44862 17935 -44238
rect 17615 -44890 17935 -44862
rect 18615 -44238 18935 -44210
rect 18615 -44862 18623 -44238
rect 18927 -44862 18935 -44238
rect 18615 -44890 18935 -44862
rect 19615 -44238 19935 -44210
rect 19615 -44862 19623 -44238
rect 19927 -44862 19935 -44238
rect 19615 -44890 19935 -44862
rect 20615 -44238 20935 -44210
rect 20615 -44862 20623 -44238
rect 20927 -44862 20935 -44238
rect 20615 -44890 20935 -44862
rect 21615 -44238 21935 -44210
rect 21615 -44862 21623 -44238
rect 21927 -44862 21935 -44238
rect 21615 -44890 21935 -44862
rect 22615 -44238 22935 -44210
rect 22615 -44862 22623 -44238
rect 22927 -44862 22935 -44238
rect 22615 -44890 22935 -44862
rect 23615 -44238 23935 -44210
rect 23615 -44862 23623 -44238
rect 23927 -44862 23935 -44238
rect 23615 -44890 23935 -44862
rect 24615 -44238 24935 -44210
rect 24615 -44862 24623 -44238
rect 24927 -44862 24935 -44238
rect 24615 -44890 24935 -44862
rect 25615 -44238 25935 -44210
rect 25615 -44862 25623 -44238
rect 25927 -44862 25935 -44238
rect 25615 -44890 25935 -44862
rect 26615 -44238 26935 -44210
rect 26615 -44862 26623 -44238
rect 26927 -44862 26935 -44238
rect 26615 -44890 26935 -44862
rect 27615 -44238 27935 -44210
rect 27615 -44862 27623 -44238
rect 27927 -44862 27935 -44238
rect 27615 -44890 27935 -44862
rect 28615 -44238 28935 -44210
rect 28615 -44862 28623 -44238
rect 28927 -44862 28935 -44238
rect 28615 -44890 28935 -44862
rect 29615 -44238 29935 -44210
rect 29615 -44862 29623 -44238
rect 29927 -44862 29935 -44238
rect 29615 -44890 29935 -44862
rect 30615 -44238 30935 -44210
rect 30615 -44862 30623 -44238
rect 30927 -44862 30935 -44238
rect 30615 -44890 30935 -44862
rect 31615 -44238 31935 -44210
rect 31615 -44862 31623 -44238
rect 31927 -44862 31935 -44238
rect 31615 -44890 31935 -44862
rect 32615 -44238 32935 -44210
rect 32615 -44862 32623 -44238
rect 32927 -44862 32935 -44238
rect 32615 -44890 32935 -44862
rect 33615 -44238 33935 -44210
rect 33615 -44862 33623 -44238
rect 33927 -44862 33935 -44238
rect 33615 -44890 33935 -44862
rect -74825 -44898 -48825 -44890
rect -74825 -45202 -74817 -44898
rect -74513 -45202 -74477 -44898
rect -74173 -45202 -74137 -44898
rect -73513 -45202 -73477 -44898
rect -73173 -45202 -73137 -44898
rect -72513 -45202 -72477 -44898
rect -72173 -45202 -72137 -44898
rect -71513 -45202 -71477 -44898
rect -71173 -45202 -71137 -44898
rect -70513 -45202 -70477 -44898
rect -70173 -45202 -70137 -44898
rect -69513 -45202 -69477 -44898
rect -69173 -45202 -69137 -44898
rect -68513 -45202 -68477 -44898
rect -68173 -45202 -68137 -44898
rect -67513 -45202 -67477 -44898
rect -67173 -45202 -67137 -44898
rect -66513 -45202 -66477 -44898
rect -66173 -45202 -66137 -44898
rect -65513 -45202 -65477 -44898
rect -65173 -45202 -65137 -44898
rect -64513 -45202 -64477 -44898
rect -64173 -45202 -64137 -44898
rect -63513 -45202 -63477 -44898
rect -63173 -45202 -63137 -44898
rect -62513 -45202 -62477 -44898
rect -62173 -45202 -62137 -44898
rect -61513 -45202 -61477 -44898
rect -61173 -45202 -61137 -44898
rect -60513 -45202 -60477 -44898
rect -60173 -45202 -60137 -44898
rect -59513 -45202 -59477 -44898
rect -59173 -45202 -59137 -44898
rect -58513 -45202 -58477 -44898
rect -58173 -45202 -58137 -44898
rect -57513 -45202 -57477 -44898
rect -57173 -45202 -57137 -44898
rect -56513 -45202 -56477 -44898
rect -56173 -45202 -56137 -44898
rect -55513 -45202 -55477 -44898
rect -55173 -45202 -55137 -44898
rect -54513 -45202 -54477 -44898
rect -54173 -45202 -54137 -44898
rect -53513 -45202 -53477 -44898
rect -53173 -45202 -53137 -44898
rect -52513 -45202 -52477 -44898
rect -52173 -45202 -52137 -44898
rect -51513 -45202 -51477 -44898
rect -51173 -45202 -51137 -44898
rect -50513 -45202 -50477 -44898
rect -50173 -45202 -50137 -44898
rect -49513 -45202 -49477 -44898
rect -49173 -45202 -49137 -44898
rect -48833 -45202 -48825 -44898
rect -74825 -45210 -48825 -45202
rect 8275 -44898 34275 -44890
rect 8275 -45202 8283 -44898
rect 8587 -45202 8623 -44898
rect 8927 -45202 8963 -44898
rect 9587 -45202 9623 -44898
rect 9927 -45202 9963 -44898
rect 10587 -45202 10623 -44898
rect 10927 -45202 10963 -44898
rect 11587 -45202 11623 -44898
rect 11927 -45202 11963 -44898
rect 12587 -45202 12623 -44898
rect 12927 -45202 12963 -44898
rect 13587 -45202 13623 -44898
rect 13927 -45202 13963 -44898
rect 14587 -45202 14623 -44898
rect 14927 -45202 14963 -44898
rect 15587 -45202 15623 -44898
rect 15927 -45202 15963 -44898
rect 16587 -45202 16623 -44898
rect 16927 -45202 16963 -44898
rect 17587 -45202 17623 -44898
rect 17927 -45202 17963 -44898
rect 18587 -45202 18623 -44898
rect 18927 -45202 18963 -44898
rect 19587 -45202 19623 -44898
rect 19927 -45202 19963 -44898
rect 20587 -45202 20623 -44898
rect 20927 -45202 20963 -44898
rect 21587 -45202 21623 -44898
rect 21927 -45202 21963 -44898
rect 22587 -45202 22623 -44898
rect 22927 -45202 22963 -44898
rect 23587 -45202 23623 -44898
rect 23927 -45202 23963 -44898
rect 24587 -45202 24623 -44898
rect 24927 -45202 24963 -44898
rect 25587 -45202 25623 -44898
rect 25927 -45202 25963 -44898
rect 26587 -45202 26623 -44898
rect 26927 -45202 26963 -44898
rect 27587 -45202 27623 -44898
rect 27927 -45202 27963 -44898
rect 28587 -45202 28623 -44898
rect 28927 -45202 28963 -44898
rect 29587 -45202 29623 -44898
rect 29927 -45202 29963 -44898
rect 30587 -45202 30623 -44898
rect 30927 -45202 30963 -44898
rect 31587 -45202 31623 -44898
rect 31927 -45202 31963 -44898
rect 32587 -45202 32623 -44898
rect 32927 -45202 32963 -44898
rect 33587 -45202 33623 -44898
rect 33927 -45202 33963 -44898
rect 34267 -45202 34275 -44898
rect 8275 -45210 34275 -45202
rect -74485 -45238 -74165 -45210
rect -74485 -45862 -74477 -45238
rect -74173 -45862 -74165 -45238
rect -74485 -45890 -74165 -45862
rect -73485 -45238 -73165 -45210
rect -73485 -45862 -73477 -45238
rect -73173 -45862 -73165 -45238
rect -73485 -45890 -73165 -45862
rect -72485 -45238 -72165 -45210
rect -72485 -45862 -72477 -45238
rect -72173 -45862 -72165 -45238
rect -72485 -45890 -72165 -45862
rect -71485 -45238 -71165 -45210
rect -71485 -45862 -71477 -45238
rect -71173 -45862 -71165 -45238
rect -71485 -45890 -71165 -45862
rect -70485 -45238 -70165 -45210
rect -70485 -45862 -70477 -45238
rect -70173 -45862 -70165 -45238
rect -70485 -45890 -70165 -45862
rect -69485 -45238 -69165 -45210
rect -69485 -45862 -69477 -45238
rect -69173 -45862 -69165 -45238
rect -69485 -45890 -69165 -45862
rect -68485 -45238 -68165 -45210
rect -68485 -45862 -68477 -45238
rect -68173 -45862 -68165 -45238
rect -68485 -45890 -68165 -45862
rect -67485 -45238 -67165 -45210
rect -67485 -45862 -67477 -45238
rect -67173 -45862 -67165 -45238
rect -67485 -45890 -67165 -45862
rect -66485 -45238 -66165 -45210
rect -66485 -45862 -66477 -45238
rect -66173 -45862 -66165 -45238
rect -66485 -45890 -66165 -45862
rect -65485 -45238 -65165 -45210
rect -65485 -45862 -65477 -45238
rect -65173 -45862 -65165 -45238
rect -65485 -45890 -65165 -45862
rect -64485 -45238 -64165 -45210
rect -64485 -45862 -64477 -45238
rect -64173 -45862 -64165 -45238
rect -64485 -45890 -64165 -45862
rect -63485 -45238 -63165 -45210
rect -63485 -45862 -63477 -45238
rect -63173 -45862 -63165 -45238
rect -63485 -45890 -63165 -45862
rect -62485 -45238 -62165 -45210
rect -62485 -45862 -62477 -45238
rect -62173 -45862 -62165 -45238
rect -62485 -45890 -62165 -45862
rect -61485 -45238 -61165 -45210
rect -61485 -45862 -61477 -45238
rect -61173 -45862 -61165 -45238
rect -61485 -45890 -61165 -45862
rect -60485 -45238 -60165 -45210
rect -60485 -45862 -60477 -45238
rect -60173 -45862 -60165 -45238
rect -60485 -45890 -60165 -45862
rect -59485 -45238 -59165 -45210
rect -59485 -45862 -59477 -45238
rect -59173 -45862 -59165 -45238
rect -59485 -45890 -59165 -45862
rect -58485 -45238 -58165 -45210
rect -58485 -45862 -58477 -45238
rect -58173 -45862 -58165 -45238
rect -58485 -45890 -58165 -45862
rect -57485 -45238 -57165 -45210
rect -57485 -45862 -57477 -45238
rect -57173 -45862 -57165 -45238
rect -57485 -45890 -57165 -45862
rect -56485 -45238 -56165 -45210
rect -56485 -45862 -56477 -45238
rect -56173 -45862 -56165 -45238
rect -56485 -45890 -56165 -45862
rect -55485 -45238 -55165 -45210
rect -55485 -45862 -55477 -45238
rect -55173 -45862 -55165 -45238
rect -55485 -45890 -55165 -45862
rect -54485 -45238 -54165 -45210
rect -54485 -45862 -54477 -45238
rect -54173 -45862 -54165 -45238
rect -54485 -45890 -54165 -45862
rect -53485 -45238 -53165 -45210
rect -53485 -45862 -53477 -45238
rect -53173 -45862 -53165 -45238
rect -53485 -45890 -53165 -45862
rect -52485 -45238 -52165 -45210
rect -52485 -45862 -52477 -45238
rect -52173 -45862 -52165 -45238
rect -52485 -45890 -52165 -45862
rect -51485 -45238 -51165 -45210
rect -51485 -45862 -51477 -45238
rect -51173 -45862 -51165 -45238
rect -51485 -45890 -51165 -45862
rect -50485 -45238 -50165 -45210
rect -50485 -45862 -50477 -45238
rect -50173 -45862 -50165 -45238
rect -50485 -45890 -50165 -45862
rect -49485 -45238 -49165 -45210
rect -49485 -45862 -49477 -45238
rect -49173 -45862 -49165 -45238
rect -49485 -45890 -49165 -45862
rect 8615 -45238 8935 -45210
rect 8615 -45862 8623 -45238
rect 8927 -45862 8935 -45238
rect 8615 -45890 8935 -45862
rect 9615 -45238 9935 -45210
rect 9615 -45862 9623 -45238
rect 9927 -45862 9935 -45238
rect 9615 -45890 9935 -45862
rect 10615 -45238 10935 -45210
rect 10615 -45862 10623 -45238
rect 10927 -45862 10935 -45238
rect 10615 -45890 10935 -45862
rect 11615 -45238 11935 -45210
rect 11615 -45862 11623 -45238
rect 11927 -45862 11935 -45238
rect 11615 -45890 11935 -45862
rect 12615 -45238 12935 -45210
rect 12615 -45862 12623 -45238
rect 12927 -45862 12935 -45238
rect 12615 -45890 12935 -45862
rect 13615 -45238 13935 -45210
rect 13615 -45862 13623 -45238
rect 13927 -45862 13935 -45238
rect 13615 -45890 13935 -45862
rect 14615 -45238 14935 -45210
rect 14615 -45862 14623 -45238
rect 14927 -45862 14935 -45238
rect 14615 -45890 14935 -45862
rect 15615 -45238 15935 -45210
rect 15615 -45862 15623 -45238
rect 15927 -45862 15935 -45238
rect 15615 -45890 15935 -45862
rect 16615 -45238 16935 -45210
rect 16615 -45862 16623 -45238
rect 16927 -45862 16935 -45238
rect 16615 -45890 16935 -45862
rect 17615 -45238 17935 -45210
rect 17615 -45862 17623 -45238
rect 17927 -45862 17935 -45238
rect 17615 -45890 17935 -45862
rect 18615 -45238 18935 -45210
rect 18615 -45862 18623 -45238
rect 18927 -45862 18935 -45238
rect 18615 -45890 18935 -45862
rect 19615 -45238 19935 -45210
rect 19615 -45862 19623 -45238
rect 19927 -45862 19935 -45238
rect 19615 -45890 19935 -45862
rect 20615 -45238 20935 -45210
rect 20615 -45862 20623 -45238
rect 20927 -45862 20935 -45238
rect 20615 -45890 20935 -45862
rect 21615 -45238 21935 -45210
rect 21615 -45862 21623 -45238
rect 21927 -45862 21935 -45238
rect 21615 -45890 21935 -45862
rect 22615 -45238 22935 -45210
rect 22615 -45862 22623 -45238
rect 22927 -45862 22935 -45238
rect 22615 -45890 22935 -45862
rect 23615 -45238 23935 -45210
rect 23615 -45862 23623 -45238
rect 23927 -45862 23935 -45238
rect 23615 -45890 23935 -45862
rect 24615 -45238 24935 -45210
rect 24615 -45862 24623 -45238
rect 24927 -45862 24935 -45238
rect 24615 -45890 24935 -45862
rect 25615 -45238 25935 -45210
rect 25615 -45862 25623 -45238
rect 25927 -45862 25935 -45238
rect 25615 -45890 25935 -45862
rect 26615 -45238 26935 -45210
rect 26615 -45862 26623 -45238
rect 26927 -45862 26935 -45238
rect 26615 -45890 26935 -45862
rect 27615 -45238 27935 -45210
rect 27615 -45862 27623 -45238
rect 27927 -45862 27935 -45238
rect 27615 -45890 27935 -45862
rect 28615 -45238 28935 -45210
rect 28615 -45862 28623 -45238
rect 28927 -45862 28935 -45238
rect 28615 -45890 28935 -45862
rect 29615 -45238 29935 -45210
rect 29615 -45862 29623 -45238
rect 29927 -45862 29935 -45238
rect 29615 -45890 29935 -45862
rect 30615 -45238 30935 -45210
rect 30615 -45862 30623 -45238
rect 30927 -45862 30935 -45238
rect 30615 -45890 30935 -45862
rect 31615 -45238 31935 -45210
rect 31615 -45862 31623 -45238
rect 31927 -45862 31935 -45238
rect 31615 -45890 31935 -45862
rect 32615 -45238 32935 -45210
rect 32615 -45862 32623 -45238
rect 32927 -45862 32935 -45238
rect 32615 -45890 32935 -45862
rect 33615 -45238 33935 -45210
rect 33615 -45862 33623 -45238
rect 33927 -45862 33935 -45238
rect 33615 -45890 33935 -45862
rect -74825 -45898 -48825 -45890
rect -74825 -46202 -74817 -45898
rect -74513 -46202 -74477 -45898
rect -74173 -46202 -74137 -45898
rect -73513 -46202 -73477 -45898
rect -73173 -46202 -73137 -45898
rect -72513 -46202 -72477 -45898
rect -72173 -46202 -72137 -45898
rect -71513 -46202 -71477 -45898
rect -71173 -46202 -71137 -45898
rect -70513 -46202 -70477 -45898
rect -70173 -46202 -70137 -45898
rect -69513 -46202 -69477 -45898
rect -69173 -46202 -69137 -45898
rect -68513 -46202 -68477 -45898
rect -68173 -46202 -68137 -45898
rect -67513 -46202 -67477 -45898
rect -67173 -46202 -67137 -45898
rect -66513 -46202 -66477 -45898
rect -66173 -46202 -66137 -45898
rect -65513 -46202 -65477 -45898
rect -65173 -46202 -65137 -45898
rect -64513 -46202 -64477 -45898
rect -64173 -46202 -64137 -45898
rect -63513 -46202 -63477 -45898
rect -63173 -46202 -63137 -45898
rect -62513 -46202 -62477 -45898
rect -62173 -46202 -62137 -45898
rect -61513 -46202 -61477 -45898
rect -61173 -46202 -61137 -45898
rect -60513 -46202 -60477 -45898
rect -60173 -46202 -60137 -45898
rect -59513 -46202 -59477 -45898
rect -59173 -46202 -59137 -45898
rect -58513 -46202 -58477 -45898
rect -58173 -46202 -58137 -45898
rect -57513 -46202 -57477 -45898
rect -57173 -46202 -57137 -45898
rect -56513 -46202 -56477 -45898
rect -56173 -46202 -56137 -45898
rect -55513 -46202 -55477 -45898
rect -55173 -46202 -55137 -45898
rect -54513 -46202 -54477 -45898
rect -54173 -46202 -54137 -45898
rect -53513 -46202 -53477 -45898
rect -53173 -46202 -53137 -45898
rect -52513 -46202 -52477 -45898
rect -52173 -46202 -52137 -45898
rect -51513 -46202 -51477 -45898
rect -51173 -46202 -51137 -45898
rect -50513 -46202 -50477 -45898
rect -50173 -46202 -50137 -45898
rect -49513 -46202 -49477 -45898
rect -49173 -46202 -49137 -45898
rect -48833 -46202 -48825 -45898
rect -74825 -46210 -48825 -46202
rect 8275 -45898 34275 -45890
rect 8275 -46202 8283 -45898
rect 8587 -46202 8623 -45898
rect 8927 -46202 8963 -45898
rect 9587 -46202 9623 -45898
rect 9927 -46202 9963 -45898
rect 10587 -46202 10623 -45898
rect 10927 -46202 10963 -45898
rect 11587 -46202 11623 -45898
rect 11927 -46202 11963 -45898
rect 12587 -46202 12623 -45898
rect 12927 -46202 12963 -45898
rect 13587 -46202 13623 -45898
rect 13927 -46202 13963 -45898
rect 14587 -46202 14623 -45898
rect 14927 -46202 14963 -45898
rect 15587 -46202 15623 -45898
rect 15927 -46202 15963 -45898
rect 16587 -46202 16623 -45898
rect 16927 -46202 16963 -45898
rect 17587 -46202 17623 -45898
rect 17927 -46202 17963 -45898
rect 18587 -46202 18623 -45898
rect 18927 -46202 18963 -45898
rect 19587 -46202 19623 -45898
rect 19927 -46202 19963 -45898
rect 20587 -46202 20623 -45898
rect 20927 -46202 20963 -45898
rect 21587 -46202 21623 -45898
rect 21927 -46202 21963 -45898
rect 22587 -46202 22623 -45898
rect 22927 -46202 22963 -45898
rect 23587 -46202 23623 -45898
rect 23927 -46202 23963 -45898
rect 24587 -46202 24623 -45898
rect 24927 -46202 24963 -45898
rect 25587 -46202 25623 -45898
rect 25927 -46202 25963 -45898
rect 26587 -46202 26623 -45898
rect 26927 -46202 26963 -45898
rect 27587 -46202 27623 -45898
rect 27927 -46202 27963 -45898
rect 28587 -46202 28623 -45898
rect 28927 -46202 28963 -45898
rect 29587 -46202 29623 -45898
rect 29927 -46202 29963 -45898
rect 30587 -46202 30623 -45898
rect 30927 -46202 30963 -45898
rect 31587 -46202 31623 -45898
rect 31927 -46202 31963 -45898
rect 32587 -46202 32623 -45898
rect 32927 -46202 32963 -45898
rect 33587 -46202 33623 -45898
rect 33927 -46202 33963 -45898
rect 34267 -46202 34275 -45898
rect 8275 -46210 34275 -46202
rect -74485 -46238 -74165 -46210
rect -74485 -46542 -74477 -46238
rect -74173 -46542 -74165 -46238
rect -74485 -46550 -74165 -46542
rect -73485 -46238 -73165 -46210
rect -73485 -46542 -73477 -46238
rect -73173 -46542 -73165 -46238
rect -73485 -46550 -73165 -46542
rect -72485 -46238 -72165 -46210
rect -72485 -46542 -72477 -46238
rect -72173 -46542 -72165 -46238
rect -72485 -46550 -72165 -46542
rect -71485 -46238 -71165 -46210
rect -71485 -46542 -71477 -46238
rect -71173 -46542 -71165 -46238
rect -71485 -46550 -71165 -46542
rect -70485 -46238 -70165 -46210
rect -70485 -46542 -70477 -46238
rect -70173 -46542 -70165 -46238
rect -70485 -46550 -70165 -46542
rect -69485 -46238 -69165 -46210
rect -69485 -46542 -69477 -46238
rect -69173 -46542 -69165 -46238
rect -69485 -46550 -69165 -46542
rect -68485 -46238 -68165 -46210
rect -68485 -46542 -68477 -46238
rect -68173 -46542 -68165 -46238
rect -68485 -46550 -68165 -46542
rect -67485 -46238 -67165 -46210
rect -67485 -46542 -67477 -46238
rect -67173 -46542 -67165 -46238
rect -67485 -46550 -67165 -46542
rect -66485 -46238 -66165 -46210
rect -66485 -46542 -66477 -46238
rect -66173 -46542 -66165 -46238
rect -66485 -46550 -66165 -46542
rect -65485 -46238 -65165 -46210
rect -65485 -46542 -65477 -46238
rect -65173 -46542 -65165 -46238
rect -65485 -46550 -65165 -46542
rect -64485 -46238 -64165 -46210
rect -64485 -46542 -64477 -46238
rect -64173 -46542 -64165 -46238
rect -64485 -46550 -64165 -46542
rect -63485 -46238 -63165 -46210
rect -63485 -46542 -63477 -46238
rect -63173 -46542 -63165 -46238
rect -63485 -46550 -63165 -46542
rect -62485 -46238 -62165 -46210
rect -62485 -46542 -62477 -46238
rect -62173 -46542 -62165 -46238
rect -62485 -46550 -62165 -46542
rect -61485 -46238 -61165 -46210
rect -61485 -46542 -61477 -46238
rect -61173 -46542 -61165 -46238
rect -61485 -46550 -61165 -46542
rect -60485 -46238 -60165 -46210
rect -60485 -46542 -60477 -46238
rect -60173 -46542 -60165 -46238
rect -60485 -46550 -60165 -46542
rect -59485 -46238 -59165 -46210
rect -59485 -46542 -59477 -46238
rect -59173 -46542 -59165 -46238
rect -59485 -46550 -59165 -46542
rect -58485 -46238 -58165 -46210
rect -58485 -46542 -58477 -46238
rect -58173 -46542 -58165 -46238
rect -58485 -46550 -58165 -46542
rect -57485 -46238 -57165 -46210
rect -57485 -46542 -57477 -46238
rect -57173 -46542 -57165 -46238
rect -57485 -46550 -57165 -46542
rect -56485 -46238 -56165 -46210
rect -56485 -46542 -56477 -46238
rect -56173 -46542 -56165 -46238
rect -56485 -46550 -56165 -46542
rect -55485 -46238 -55165 -46210
rect -55485 -46542 -55477 -46238
rect -55173 -46542 -55165 -46238
rect -55485 -46550 -55165 -46542
rect -54485 -46238 -54165 -46210
rect -54485 -46542 -54477 -46238
rect -54173 -46542 -54165 -46238
rect -54485 -46550 -54165 -46542
rect -53485 -46238 -53165 -46210
rect -53485 -46542 -53477 -46238
rect -53173 -46542 -53165 -46238
rect -53485 -46550 -53165 -46542
rect -52485 -46238 -52165 -46210
rect -52485 -46542 -52477 -46238
rect -52173 -46542 -52165 -46238
rect -52485 -46550 -52165 -46542
rect -51485 -46238 -51165 -46210
rect -51485 -46542 -51477 -46238
rect -51173 -46542 -51165 -46238
rect -51485 -46550 -51165 -46542
rect -50485 -46238 -50165 -46210
rect -50485 -46542 -50477 -46238
rect -50173 -46542 -50165 -46238
rect -50485 -46550 -50165 -46542
rect -49485 -46238 -49165 -46210
rect -49485 -46542 -49477 -46238
rect -49173 -46542 -49165 -46238
rect -49485 -46550 -49165 -46542
rect 8615 -46238 8935 -46210
rect 8615 -46542 8623 -46238
rect 8927 -46542 8935 -46238
rect 8615 -46550 8935 -46542
rect 9615 -46238 9935 -46210
rect 9615 -46542 9623 -46238
rect 9927 -46542 9935 -46238
rect 9615 -46550 9935 -46542
rect 10615 -46238 10935 -46210
rect 10615 -46542 10623 -46238
rect 10927 -46542 10935 -46238
rect 10615 -46550 10935 -46542
rect 11615 -46238 11935 -46210
rect 11615 -46542 11623 -46238
rect 11927 -46542 11935 -46238
rect 11615 -46550 11935 -46542
rect 12615 -46238 12935 -46210
rect 12615 -46542 12623 -46238
rect 12927 -46542 12935 -46238
rect 12615 -46550 12935 -46542
rect 13615 -46238 13935 -46210
rect 13615 -46542 13623 -46238
rect 13927 -46542 13935 -46238
rect 13615 -46550 13935 -46542
rect 14615 -46238 14935 -46210
rect 14615 -46542 14623 -46238
rect 14927 -46542 14935 -46238
rect 14615 -46550 14935 -46542
rect 15615 -46238 15935 -46210
rect 15615 -46542 15623 -46238
rect 15927 -46542 15935 -46238
rect 15615 -46550 15935 -46542
rect 16615 -46238 16935 -46210
rect 16615 -46542 16623 -46238
rect 16927 -46542 16935 -46238
rect 16615 -46550 16935 -46542
rect 17615 -46238 17935 -46210
rect 17615 -46542 17623 -46238
rect 17927 -46542 17935 -46238
rect 17615 -46550 17935 -46542
rect 18615 -46238 18935 -46210
rect 18615 -46542 18623 -46238
rect 18927 -46542 18935 -46238
rect 18615 -46550 18935 -46542
rect 19615 -46238 19935 -46210
rect 19615 -46542 19623 -46238
rect 19927 -46542 19935 -46238
rect 19615 -46550 19935 -46542
rect 20615 -46238 20935 -46210
rect 20615 -46542 20623 -46238
rect 20927 -46542 20935 -46238
rect 20615 -46550 20935 -46542
rect 21615 -46238 21935 -46210
rect 21615 -46542 21623 -46238
rect 21927 -46542 21935 -46238
rect 21615 -46550 21935 -46542
rect 22615 -46238 22935 -46210
rect 22615 -46542 22623 -46238
rect 22927 -46542 22935 -46238
rect 22615 -46550 22935 -46542
rect 23615 -46238 23935 -46210
rect 23615 -46542 23623 -46238
rect 23927 -46542 23935 -46238
rect 23615 -46550 23935 -46542
rect 24615 -46238 24935 -46210
rect 24615 -46542 24623 -46238
rect 24927 -46542 24935 -46238
rect 24615 -46550 24935 -46542
rect 25615 -46238 25935 -46210
rect 25615 -46542 25623 -46238
rect 25927 -46542 25935 -46238
rect 25615 -46550 25935 -46542
rect 26615 -46238 26935 -46210
rect 26615 -46542 26623 -46238
rect 26927 -46542 26935 -46238
rect 26615 -46550 26935 -46542
rect 27615 -46238 27935 -46210
rect 27615 -46542 27623 -46238
rect 27927 -46542 27935 -46238
rect 27615 -46550 27935 -46542
rect 28615 -46238 28935 -46210
rect 28615 -46542 28623 -46238
rect 28927 -46542 28935 -46238
rect 28615 -46550 28935 -46542
rect 29615 -46238 29935 -46210
rect 29615 -46542 29623 -46238
rect 29927 -46542 29935 -46238
rect 29615 -46550 29935 -46542
rect 30615 -46238 30935 -46210
rect 30615 -46542 30623 -46238
rect 30927 -46542 30935 -46238
rect 30615 -46550 30935 -46542
rect 31615 -46238 31935 -46210
rect 31615 -46542 31623 -46238
rect 31927 -46542 31935 -46238
rect 31615 -46550 31935 -46542
rect 32615 -46238 32935 -46210
rect 32615 -46542 32623 -46238
rect 32927 -46542 32935 -46238
rect 32615 -46550 32935 -46542
rect 33615 -46238 33935 -46210
rect 33615 -46542 33623 -46238
rect 33927 -46542 33935 -46238
rect 33615 -46550 33935 -46542
<< via3 >>
rect -74477 38538 -74173 38542
rect -74477 38242 -74473 38538
rect -74473 38242 -74177 38538
rect -74177 38242 -74173 38538
rect -74477 38238 -74173 38242
rect -73477 38538 -73173 38542
rect -73477 38242 -73473 38538
rect -73473 38242 -73177 38538
rect -73177 38242 -73173 38538
rect -73477 38238 -73173 38242
rect -72477 38538 -72173 38542
rect -72477 38242 -72473 38538
rect -72473 38242 -72177 38538
rect -72177 38242 -72173 38538
rect -72477 38238 -72173 38242
rect -71477 38538 -71173 38542
rect -71477 38242 -71473 38538
rect -71473 38242 -71177 38538
rect -71177 38242 -71173 38538
rect -71477 38238 -71173 38242
rect -70477 38538 -70173 38542
rect -70477 38242 -70473 38538
rect -70473 38242 -70177 38538
rect -70177 38242 -70173 38538
rect -70477 38238 -70173 38242
rect -69477 38538 -69173 38542
rect -69477 38242 -69473 38538
rect -69473 38242 -69177 38538
rect -69177 38242 -69173 38538
rect -69477 38238 -69173 38242
rect -68477 38538 -68173 38542
rect -68477 38242 -68473 38538
rect -68473 38242 -68177 38538
rect -68177 38242 -68173 38538
rect -68477 38238 -68173 38242
rect -67477 38538 -67173 38542
rect -67477 38242 -67473 38538
rect -67473 38242 -67177 38538
rect -67177 38242 -67173 38538
rect -67477 38238 -67173 38242
rect -66477 38538 -66173 38542
rect -66477 38242 -66473 38538
rect -66473 38242 -66177 38538
rect -66177 38242 -66173 38538
rect -66477 38238 -66173 38242
rect -65477 38538 -65173 38542
rect -65477 38242 -65473 38538
rect -65473 38242 -65177 38538
rect -65177 38242 -65173 38538
rect -65477 38238 -65173 38242
rect -64477 38538 -64173 38542
rect -64477 38242 -64473 38538
rect -64473 38242 -64177 38538
rect -64177 38242 -64173 38538
rect -64477 38238 -64173 38242
rect -63477 38538 -63173 38542
rect -63477 38242 -63473 38538
rect -63473 38242 -63177 38538
rect -63177 38242 -63173 38538
rect -63477 38238 -63173 38242
rect -62477 38538 -62173 38542
rect -62477 38242 -62473 38538
rect -62473 38242 -62177 38538
rect -62177 38242 -62173 38538
rect -62477 38238 -62173 38242
rect -61477 38538 -61173 38542
rect -61477 38242 -61473 38538
rect -61473 38242 -61177 38538
rect -61177 38242 -61173 38538
rect -61477 38238 -61173 38242
rect -60477 38538 -60173 38542
rect -60477 38242 -60473 38538
rect -60473 38242 -60177 38538
rect -60177 38242 -60173 38538
rect -60477 38238 -60173 38242
rect -59477 38538 -59173 38542
rect -59477 38242 -59473 38538
rect -59473 38242 -59177 38538
rect -59177 38242 -59173 38538
rect -59477 38238 -59173 38242
rect -74817 38198 -74513 38202
rect -74817 37902 -74813 38198
rect -74813 37902 -74517 38198
rect -74517 37902 -74513 38198
rect -74817 37898 -74513 37902
rect -74477 38198 -74173 38202
rect -74477 37902 -74473 38198
rect -74473 37902 -74177 38198
rect -74177 37902 -74173 38198
rect -74477 37898 -74173 37902
rect -74137 38198 -73513 38202
rect -74137 37902 -74133 38198
rect -74133 37902 -73517 38198
rect -73517 37902 -73513 38198
rect -74137 37898 -73513 37902
rect -73477 38198 -73173 38202
rect -73477 37902 -73473 38198
rect -73473 37902 -73177 38198
rect -73177 37902 -73173 38198
rect -73477 37898 -73173 37902
rect -73137 38198 -72513 38202
rect -73137 37902 -73133 38198
rect -73133 37902 -72517 38198
rect -72517 37902 -72513 38198
rect -73137 37898 -72513 37902
rect -72477 38198 -72173 38202
rect -72477 37902 -72473 38198
rect -72473 37902 -72177 38198
rect -72177 37902 -72173 38198
rect -72477 37898 -72173 37902
rect -72137 38198 -71513 38202
rect -72137 37902 -72133 38198
rect -72133 37902 -71517 38198
rect -71517 37902 -71513 38198
rect -72137 37898 -71513 37902
rect -71477 38198 -71173 38202
rect -71477 37902 -71473 38198
rect -71473 37902 -71177 38198
rect -71177 37902 -71173 38198
rect -71477 37898 -71173 37902
rect -71137 38198 -70513 38202
rect -71137 37902 -71133 38198
rect -71133 37902 -70517 38198
rect -70517 37902 -70513 38198
rect -71137 37898 -70513 37902
rect -70477 38198 -70173 38202
rect -70477 37902 -70473 38198
rect -70473 37902 -70177 38198
rect -70177 37902 -70173 38198
rect -70477 37898 -70173 37902
rect -70137 38198 -69513 38202
rect -70137 37902 -70133 38198
rect -70133 37902 -69517 38198
rect -69517 37902 -69513 38198
rect -70137 37898 -69513 37902
rect -69477 38198 -69173 38202
rect -69477 37902 -69473 38198
rect -69473 37902 -69177 38198
rect -69177 37902 -69173 38198
rect -69477 37898 -69173 37902
rect -69137 38198 -68513 38202
rect -69137 37902 -69133 38198
rect -69133 37902 -68517 38198
rect -68517 37902 -68513 38198
rect -69137 37898 -68513 37902
rect -68477 38198 -68173 38202
rect -68477 37902 -68473 38198
rect -68473 37902 -68177 38198
rect -68177 37902 -68173 38198
rect -68477 37898 -68173 37902
rect -68137 38198 -67513 38202
rect -68137 37902 -68133 38198
rect -68133 37902 -67517 38198
rect -67517 37902 -67513 38198
rect -68137 37898 -67513 37902
rect -67477 38198 -67173 38202
rect -67477 37902 -67473 38198
rect -67473 37902 -67177 38198
rect -67177 37902 -67173 38198
rect -67477 37898 -67173 37902
rect -67137 38198 -66513 38202
rect -67137 37902 -67133 38198
rect -67133 37902 -66517 38198
rect -66517 37902 -66513 38198
rect -67137 37898 -66513 37902
rect -66477 38198 -66173 38202
rect -66477 37902 -66473 38198
rect -66473 37902 -66177 38198
rect -66177 37902 -66173 38198
rect -66477 37898 -66173 37902
rect -66137 38198 -65513 38202
rect -66137 37902 -66133 38198
rect -66133 37902 -65517 38198
rect -65517 37902 -65513 38198
rect -66137 37898 -65513 37902
rect -65477 38198 -65173 38202
rect -65477 37902 -65473 38198
rect -65473 37902 -65177 38198
rect -65177 37902 -65173 38198
rect -65477 37898 -65173 37902
rect -65137 38198 -64513 38202
rect -65137 37902 -65133 38198
rect -65133 37902 -64517 38198
rect -64517 37902 -64513 38198
rect -65137 37898 -64513 37902
rect -64477 38198 -64173 38202
rect -64477 37902 -64473 38198
rect -64473 37902 -64177 38198
rect -64177 37902 -64173 38198
rect -64477 37898 -64173 37902
rect -64137 38198 -63513 38202
rect -64137 37902 -64133 38198
rect -64133 37902 -63517 38198
rect -63517 37902 -63513 38198
rect -64137 37898 -63513 37902
rect -63477 38198 -63173 38202
rect -63477 37902 -63473 38198
rect -63473 37902 -63177 38198
rect -63177 37902 -63173 38198
rect -63477 37898 -63173 37902
rect -63137 38198 -62513 38202
rect -63137 37902 -63133 38198
rect -63133 37902 -62517 38198
rect -62517 37902 -62513 38198
rect -63137 37898 -62513 37902
rect -62477 38198 -62173 38202
rect -62477 37902 -62473 38198
rect -62473 37902 -62177 38198
rect -62177 37902 -62173 38198
rect -62477 37898 -62173 37902
rect -62137 38198 -61513 38202
rect -62137 37902 -62133 38198
rect -62133 37902 -61517 38198
rect -61517 37902 -61513 38198
rect -62137 37898 -61513 37902
rect -61477 38198 -61173 38202
rect -61477 37902 -61473 38198
rect -61473 37902 -61177 38198
rect -61177 37902 -61173 38198
rect -61477 37898 -61173 37902
rect -61137 38198 -60513 38202
rect -61137 37902 -61133 38198
rect -61133 37902 -60517 38198
rect -60517 37902 -60513 38198
rect -61137 37898 -60513 37902
rect -60477 38198 -60173 38202
rect -60477 37902 -60473 38198
rect -60473 37902 -60177 38198
rect -60177 37902 -60173 38198
rect -60477 37898 -60173 37902
rect -60137 38198 -59513 38202
rect -60137 37902 -60133 38198
rect -60133 37902 -59517 38198
rect -59517 37902 -59513 38198
rect -60137 37898 -59513 37902
rect -59477 38198 -59173 38202
rect -59477 37902 -59473 38198
rect -59473 37902 -59177 38198
rect -59177 37902 -59173 38198
rect -59477 37898 -59173 37902
rect -59137 38198 -58833 38202
rect -59137 37902 -59133 38198
rect -59133 37902 -58837 38198
rect -58837 37902 -58833 38198
rect -59137 37898 -58833 37902
rect -74477 37858 -74173 37862
rect -74477 37242 -74473 37858
rect -74473 37242 -74177 37858
rect -74177 37242 -74173 37858
rect -74477 37238 -74173 37242
rect -73477 37858 -73173 37862
rect -73477 37242 -73473 37858
rect -73473 37242 -73177 37858
rect -73177 37242 -73173 37858
rect -73477 37238 -73173 37242
rect -72477 37858 -72173 37862
rect -72477 37242 -72473 37858
rect -72473 37242 -72177 37858
rect -72177 37242 -72173 37858
rect -72477 37238 -72173 37242
rect -71477 37858 -71173 37862
rect -71477 37242 -71473 37858
rect -71473 37242 -71177 37858
rect -71177 37242 -71173 37858
rect -71477 37238 -71173 37242
rect -70477 37858 -70173 37862
rect -70477 37242 -70473 37858
rect -70473 37242 -70177 37858
rect -70177 37242 -70173 37858
rect -70477 37238 -70173 37242
rect -69477 37858 -69173 37862
rect -69477 37242 -69473 37858
rect -69473 37242 -69177 37858
rect -69177 37242 -69173 37858
rect -69477 37238 -69173 37242
rect -68477 37858 -68173 37862
rect -68477 37242 -68473 37858
rect -68473 37242 -68177 37858
rect -68177 37242 -68173 37858
rect -68477 37238 -68173 37242
rect -67477 37858 -67173 37862
rect -67477 37242 -67473 37858
rect -67473 37242 -67177 37858
rect -67177 37242 -67173 37858
rect -67477 37238 -67173 37242
rect -66477 37858 -66173 37862
rect -66477 37242 -66473 37858
rect -66473 37242 -66177 37858
rect -66177 37242 -66173 37858
rect -66477 37238 -66173 37242
rect -65477 37858 -65173 37862
rect -65477 37242 -65473 37858
rect -65473 37242 -65177 37858
rect -65177 37242 -65173 37858
rect -65477 37238 -65173 37242
rect -64477 37858 -64173 37862
rect -64477 37242 -64473 37858
rect -64473 37242 -64177 37858
rect -64177 37242 -64173 37858
rect -64477 37238 -64173 37242
rect -63477 37858 -63173 37862
rect -63477 37242 -63473 37858
rect -63473 37242 -63177 37858
rect -63177 37242 -63173 37858
rect -63477 37238 -63173 37242
rect -62477 37858 -62173 37862
rect -62477 37242 -62473 37858
rect -62473 37242 -62177 37858
rect -62177 37242 -62173 37858
rect -62477 37238 -62173 37242
rect -61477 37858 -61173 37862
rect -61477 37242 -61473 37858
rect -61473 37242 -61177 37858
rect -61177 37242 -61173 37858
rect -61477 37238 -61173 37242
rect -60477 37858 -60173 37862
rect -60477 37242 -60473 37858
rect -60473 37242 -60177 37858
rect -60177 37242 -60173 37858
rect -60477 37238 -60173 37242
rect -59477 37858 -59173 37862
rect -59477 37242 -59473 37858
rect -59473 37242 -59177 37858
rect -59177 37242 -59173 37858
rect -59477 37238 -59173 37242
rect -74817 37198 -74513 37202
rect -74817 36902 -74813 37198
rect -74813 36902 -74517 37198
rect -74517 36902 -74513 37198
rect -74817 36898 -74513 36902
rect -74477 37198 -74173 37202
rect -74477 36902 -74473 37198
rect -74473 36902 -74177 37198
rect -74177 36902 -74173 37198
rect -74477 36898 -74173 36902
rect -74137 37198 -73513 37202
rect -74137 36902 -74133 37198
rect -74133 36902 -73517 37198
rect -73517 36902 -73513 37198
rect -74137 36898 -73513 36902
rect -73477 37198 -73173 37202
rect -73477 36902 -73473 37198
rect -73473 36902 -73177 37198
rect -73177 36902 -73173 37198
rect -73477 36898 -73173 36902
rect -73137 37198 -72513 37202
rect -73137 36902 -73133 37198
rect -73133 36902 -72517 37198
rect -72517 36902 -72513 37198
rect -73137 36898 -72513 36902
rect -72477 37198 -72173 37202
rect -72477 36902 -72473 37198
rect -72473 36902 -72177 37198
rect -72177 36902 -72173 37198
rect -72477 36898 -72173 36902
rect -72137 37198 -71513 37202
rect -72137 36902 -72133 37198
rect -72133 36902 -71517 37198
rect -71517 36902 -71513 37198
rect -72137 36898 -71513 36902
rect -71477 37198 -71173 37202
rect -71477 36902 -71473 37198
rect -71473 36902 -71177 37198
rect -71177 36902 -71173 37198
rect -71477 36898 -71173 36902
rect -71137 37198 -70513 37202
rect -71137 36902 -71133 37198
rect -71133 36902 -70517 37198
rect -70517 36902 -70513 37198
rect -71137 36898 -70513 36902
rect -70477 37198 -70173 37202
rect -70477 36902 -70473 37198
rect -70473 36902 -70177 37198
rect -70177 36902 -70173 37198
rect -70477 36898 -70173 36902
rect -70137 37198 -69513 37202
rect -70137 36902 -70133 37198
rect -70133 36902 -69517 37198
rect -69517 36902 -69513 37198
rect -70137 36898 -69513 36902
rect -69477 37198 -69173 37202
rect -69477 36902 -69473 37198
rect -69473 36902 -69177 37198
rect -69177 36902 -69173 37198
rect -69477 36898 -69173 36902
rect -69137 37198 -68513 37202
rect -69137 36902 -69133 37198
rect -69133 36902 -68517 37198
rect -68517 36902 -68513 37198
rect -69137 36898 -68513 36902
rect -68477 37198 -68173 37202
rect -68477 36902 -68473 37198
rect -68473 36902 -68177 37198
rect -68177 36902 -68173 37198
rect -68477 36898 -68173 36902
rect -68137 37198 -67513 37202
rect -68137 36902 -68133 37198
rect -68133 36902 -67517 37198
rect -67517 36902 -67513 37198
rect -68137 36898 -67513 36902
rect -67477 37198 -67173 37202
rect -67477 36902 -67473 37198
rect -67473 36902 -67177 37198
rect -67177 36902 -67173 37198
rect -67477 36898 -67173 36902
rect -67137 37198 -66513 37202
rect -67137 36902 -67133 37198
rect -67133 36902 -66517 37198
rect -66517 36902 -66513 37198
rect -67137 36898 -66513 36902
rect -66477 37198 -66173 37202
rect -66477 36902 -66473 37198
rect -66473 36902 -66177 37198
rect -66177 36902 -66173 37198
rect -66477 36898 -66173 36902
rect -66137 37198 -65513 37202
rect -66137 36902 -66133 37198
rect -66133 36902 -65517 37198
rect -65517 36902 -65513 37198
rect -66137 36898 -65513 36902
rect -65477 37198 -65173 37202
rect -65477 36902 -65473 37198
rect -65473 36902 -65177 37198
rect -65177 36902 -65173 37198
rect -65477 36898 -65173 36902
rect -65137 37198 -64513 37202
rect -65137 36902 -65133 37198
rect -65133 36902 -64517 37198
rect -64517 36902 -64513 37198
rect -65137 36898 -64513 36902
rect -64477 37198 -64173 37202
rect -64477 36902 -64473 37198
rect -64473 36902 -64177 37198
rect -64177 36902 -64173 37198
rect -64477 36898 -64173 36902
rect -64137 37198 -63513 37202
rect -64137 36902 -64133 37198
rect -64133 36902 -63517 37198
rect -63517 36902 -63513 37198
rect -64137 36898 -63513 36902
rect -63477 37198 -63173 37202
rect -63477 36902 -63473 37198
rect -63473 36902 -63177 37198
rect -63177 36902 -63173 37198
rect -63477 36898 -63173 36902
rect -63137 37198 -62513 37202
rect -63137 36902 -63133 37198
rect -63133 36902 -62517 37198
rect -62517 36902 -62513 37198
rect -63137 36898 -62513 36902
rect -62477 37198 -62173 37202
rect -62477 36902 -62473 37198
rect -62473 36902 -62177 37198
rect -62177 36902 -62173 37198
rect -62477 36898 -62173 36902
rect -62137 37198 -61513 37202
rect -62137 36902 -62133 37198
rect -62133 36902 -61517 37198
rect -61517 36902 -61513 37198
rect -62137 36898 -61513 36902
rect -61477 37198 -61173 37202
rect -61477 36902 -61473 37198
rect -61473 36902 -61177 37198
rect -61177 36902 -61173 37198
rect -61477 36898 -61173 36902
rect -61137 37198 -60513 37202
rect -61137 36902 -61133 37198
rect -61133 36902 -60517 37198
rect -60517 36902 -60513 37198
rect -61137 36898 -60513 36902
rect -60477 37198 -60173 37202
rect -60477 36902 -60473 37198
rect -60473 36902 -60177 37198
rect -60177 36902 -60173 37198
rect -60477 36898 -60173 36902
rect -60137 37198 -59513 37202
rect -60137 36902 -60133 37198
rect -60133 36902 -59517 37198
rect -59517 36902 -59513 37198
rect -60137 36898 -59513 36902
rect -59477 37198 -59173 37202
rect -59477 36902 -59473 37198
rect -59473 36902 -59177 37198
rect -59177 36902 -59173 37198
rect -59477 36898 -59173 36902
rect -59137 37198 -58833 37202
rect -59137 36902 -59133 37198
rect -59133 36902 -58837 37198
rect -58837 36902 -58833 37198
rect -59137 36898 -58833 36902
rect -74477 36858 -74173 36862
rect -74477 36242 -74473 36858
rect -74473 36242 -74177 36858
rect -74177 36242 -74173 36858
rect -74477 36238 -74173 36242
rect -73477 36858 -73173 36862
rect -73477 36242 -73473 36858
rect -73473 36242 -73177 36858
rect -73177 36242 -73173 36858
rect -73477 36238 -73173 36242
rect -72477 36858 -72173 36862
rect -72477 36242 -72473 36858
rect -72473 36242 -72177 36858
rect -72177 36242 -72173 36858
rect -72477 36238 -72173 36242
rect -71477 36858 -71173 36862
rect -71477 36242 -71473 36858
rect -71473 36242 -71177 36858
rect -71177 36242 -71173 36858
rect -71477 36238 -71173 36242
rect -70477 36858 -70173 36862
rect -70477 36242 -70473 36858
rect -70473 36242 -70177 36858
rect -70177 36242 -70173 36858
rect -70477 36238 -70173 36242
rect -69477 36858 -69173 36862
rect -69477 36242 -69473 36858
rect -69473 36242 -69177 36858
rect -69177 36242 -69173 36858
rect -69477 36238 -69173 36242
rect -68477 36858 -68173 36862
rect -68477 36242 -68473 36858
rect -68473 36242 -68177 36858
rect -68177 36242 -68173 36858
rect -68477 36238 -68173 36242
rect -67477 36858 -67173 36862
rect -67477 36242 -67473 36858
rect -67473 36242 -67177 36858
rect -67177 36242 -67173 36858
rect -67477 36238 -67173 36242
rect -66477 36858 -66173 36862
rect -66477 36242 -66473 36858
rect -66473 36242 -66177 36858
rect -66177 36242 -66173 36858
rect -66477 36238 -66173 36242
rect -65477 36858 -65173 36862
rect -65477 36242 -65473 36858
rect -65473 36242 -65177 36858
rect -65177 36242 -65173 36858
rect -65477 36238 -65173 36242
rect -64477 36858 -64173 36862
rect -64477 36242 -64473 36858
rect -64473 36242 -64177 36858
rect -64177 36242 -64173 36858
rect -64477 36238 -64173 36242
rect -63477 36858 -63173 36862
rect -63477 36242 -63473 36858
rect -63473 36242 -63177 36858
rect -63177 36242 -63173 36858
rect -63477 36238 -63173 36242
rect -62477 36858 -62173 36862
rect -62477 36242 -62473 36858
rect -62473 36242 -62177 36858
rect -62177 36242 -62173 36858
rect -62477 36238 -62173 36242
rect -61477 36858 -61173 36862
rect -61477 36242 -61473 36858
rect -61473 36242 -61177 36858
rect -61177 36242 -61173 36858
rect -61477 36238 -61173 36242
rect -60477 36858 -60173 36862
rect -60477 36242 -60473 36858
rect -60473 36242 -60177 36858
rect -60177 36242 -60173 36858
rect -60477 36238 -60173 36242
rect -59477 36858 -59173 36862
rect -59477 36242 -59473 36858
rect -59473 36242 -59177 36858
rect -59177 36242 -59173 36858
rect -59477 36238 -59173 36242
rect -74817 36198 -74513 36202
rect -74817 35902 -74813 36198
rect -74813 35902 -74517 36198
rect -74517 35902 -74513 36198
rect -74817 35898 -74513 35902
rect -74477 36198 -74173 36202
rect -74477 35902 -74473 36198
rect -74473 35902 -74177 36198
rect -74177 35902 -74173 36198
rect -74477 35898 -74173 35902
rect -74137 36198 -73513 36202
rect -74137 35902 -74133 36198
rect -74133 35902 -73517 36198
rect -73517 35902 -73513 36198
rect -74137 35898 -73513 35902
rect -73477 36198 -73173 36202
rect -73477 35902 -73473 36198
rect -73473 35902 -73177 36198
rect -73177 35902 -73173 36198
rect -73477 35898 -73173 35902
rect -73137 36198 -72513 36202
rect -73137 35902 -73133 36198
rect -73133 35902 -72517 36198
rect -72517 35902 -72513 36198
rect -73137 35898 -72513 35902
rect -72477 36198 -72173 36202
rect -72477 35902 -72473 36198
rect -72473 35902 -72177 36198
rect -72177 35902 -72173 36198
rect -72477 35898 -72173 35902
rect -72137 36198 -71513 36202
rect -72137 35902 -72133 36198
rect -72133 35902 -71517 36198
rect -71517 35902 -71513 36198
rect -72137 35898 -71513 35902
rect -71477 36198 -71173 36202
rect -71477 35902 -71473 36198
rect -71473 35902 -71177 36198
rect -71177 35902 -71173 36198
rect -71477 35898 -71173 35902
rect -71137 36198 -70513 36202
rect -71137 35902 -71133 36198
rect -71133 35902 -70517 36198
rect -70517 35902 -70513 36198
rect -71137 35898 -70513 35902
rect -70477 36198 -70173 36202
rect -70477 35902 -70473 36198
rect -70473 35902 -70177 36198
rect -70177 35902 -70173 36198
rect -70477 35898 -70173 35902
rect -70137 36198 -69513 36202
rect -70137 35902 -70133 36198
rect -70133 35902 -69517 36198
rect -69517 35902 -69513 36198
rect -70137 35898 -69513 35902
rect -69477 36198 -69173 36202
rect -69477 35902 -69473 36198
rect -69473 35902 -69177 36198
rect -69177 35902 -69173 36198
rect -69477 35898 -69173 35902
rect -69137 36198 -68513 36202
rect -69137 35902 -69133 36198
rect -69133 35902 -68517 36198
rect -68517 35902 -68513 36198
rect -69137 35898 -68513 35902
rect -68477 36198 -68173 36202
rect -68477 35902 -68473 36198
rect -68473 35902 -68177 36198
rect -68177 35902 -68173 36198
rect -68477 35898 -68173 35902
rect -68137 36198 -67513 36202
rect -68137 35902 -68133 36198
rect -68133 35902 -67517 36198
rect -67517 35902 -67513 36198
rect -68137 35898 -67513 35902
rect -67477 36198 -67173 36202
rect -67477 35902 -67473 36198
rect -67473 35902 -67177 36198
rect -67177 35902 -67173 36198
rect -67477 35898 -67173 35902
rect -67137 36198 -66513 36202
rect -67137 35902 -67133 36198
rect -67133 35902 -66517 36198
rect -66517 35902 -66513 36198
rect -67137 35898 -66513 35902
rect -66477 36198 -66173 36202
rect -66477 35902 -66473 36198
rect -66473 35902 -66177 36198
rect -66177 35902 -66173 36198
rect -66477 35898 -66173 35902
rect -66137 36198 -65513 36202
rect -66137 35902 -66133 36198
rect -66133 35902 -65517 36198
rect -65517 35902 -65513 36198
rect -66137 35898 -65513 35902
rect -65477 36198 -65173 36202
rect -65477 35902 -65473 36198
rect -65473 35902 -65177 36198
rect -65177 35902 -65173 36198
rect -65477 35898 -65173 35902
rect -65137 36198 -64513 36202
rect -65137 35902 -65133 36198
rect -65133 35902 -64517 36198
rect -64517 35902 -64513 36198
rect -65137 35898 -64513 35902
rect -64477 36198 -64173 36202
rect -64477 35902 -64473 36198
rect -64473 35902 -64177 36198
rect -64177 35902 -64173 36198
rect -64477 35898 -64173 35902
rect -64137 36198 -63513 36202
rect -64137 35902 -64133 36198
rect -64133 35902 -63517 36198
rect -63517 35902 -63513 36198
rect -64137 35898 -63513 35902
rect -63477 36198 -63173 36202
rect -63477 35902 -63473 36198
rect -63473 35902 -63177 36198
rect -63177 35902 -63173 36198
rect -63477 35898 -63173 35902
rect -63137 36198 -62513 36202
rect -63137 35902 -63133 36198
rect -63133 35902 -62517 36198
rect -62517 35902 -62513 36198
rect -63137 35898 -62513 35902
rect -62477 36198 -62173 36202
rect -62477 35902 -62473 36198
rect -62473 35902 -62177 36198
rect -62177 35902 -62173 36198
rect -62477 35898 -62173 35902
rect -62137 36198 -61513 36202
rect -62137 35902 -62133 36198
rect -62133 35902 -61517 36198
rect -61517 35902 -61513 36198
rect -62137 35898 -61513 35902
rect -61477 36198 -61173 36202
rect -61477 35902 -61473 36198
rect -61473 35902 -61177 36198
rect -61177 35902 -61173 36198
rect -61477 35898 -61173 35902
rect -61137 36198 -60513 36202
rect -61137 35902 -61133 36198
rect -61133 35902 -60517 36198
rect -60517 35902 -60513 36198
rect -61137 35898 -60513 35902
rect -60477 36198 -60173 36202
rect -60477 35902 -60473 36198
rect -60473 35902 -60177 36198
rect -60177 35902 -60173 36198
rect -60477 35898 -60173 35902
rect -60137 36198 -59513 36202
rect -60137 35902 -60133 36198
rect -60133 35902 -59517 36198
rect -59517 35902 -59513 36198
rect -60137 35898 -59513 35902
rect -59477 36198 -59173 36202
rect -59477 35902 -59473 36198
rect -59473 35902 -59177 36198
rect -59177 35902 -59173 36198
rect -59477 35898 -59173 35902
rect -59137 36198 -58833 36202
rect -59137 35902 -59133 36198
rect -59133 35902 -58837 36198
rect -58837 35902 -58833 36198
rect -59137 35898 -58833 35902
rect -74477 35858 -74173 35862
rect -74477 35242 -74473 35858
rect -74473 35242 -74177 35858
rect -74177 35242 -74173 35858
rect -74477 35238 -74173 35242
rect -73477 35858 -73173 35862
rect -73477 35242 -73473 35858
rect -73473 35242 -73177 35858
rect -73177 35242 -73173 35858
rect -73477 35238 -73173 35242
rect -72477 35858 -72173 35862
rect -72477 35242 -72473 35858
rect -72473 35242 -72177 35858
rect -72177 35242 -72173 35858
rect -72477 35238 -72173 35242
rect -71477 35858 -71173 35862
rect -71477 35242 -71473 35858
rect -71473 35242 -71177 35858
rect -71177 35242 -71173 35858
rect -71477 35238 -71173 35242
rect -70477 35858 -70173 35862
rect -70477 35242 -70473 35858
rect -70473 35242 -70177 35858
rect -70177 35242 -70173 35858
rect -70477 35238 -70173 35242
rect -69477 35858 -69173 35862
rect -69477 35242 -69473 35858
rect -69473 35242 -69177 35858
rect -69177 35242 -69173 35858
rect -69477 35238 -69173 35242
rect -68477 35858 -68173 35862
rect -68477 35242 -68473 35858
rect -68473 35242 -68177 35858
rect -68177 35242 -68173 35858
rect -68477 35238 -68173 35242
rect -67477 35858 -67173 35862
rect -67477 35242 -67473 35858
rect -67473 35242 -67177 35858
rect -67177 35242 -67173 35858
rect -67477 35238 -67173 35242
rect -66477 35858 -66173 35862
rect -66477 35242 -66473 35858
rect -66473 35242 -66177 35858
rect -66177 35242 -66173 35858
rect -66477 35238 -66173 35242
rect -65477 35858 -65173 35862
rect -65477 35242 -65473 35858
rect -65473 35242 -65177 35858
rect -65177 35242 -65173 35858
rect -65477 35238 -65173 35242
rect -64477 35858 -64173 35862
rect -64477 35242 -64473 35858
rect -64473 35242 -64177 35858
rect -64177 35242 -64173 35858
rect -64477 35238 -64173 35242
rect -63477 35858 -63173 35862
rect -63477 35242 -63473 35858
rect -63473 35242 -63177 35858
rect -63177 35242 -63173 35858
rect -63477 35238 -63173 35242
rect -62477 35858 -62173 35862
rect -62477 35242 -62473 35858
rect -62473 35242 -62177 35858
rect -62177 35242 -62173 35858
rect -62477 35238 -62173 35242
rect -61477 35858 -61173 35862
rect -61477 35242 -61473 35858
rect -61473 35242 -61177 35858
rect -61177 35242 -61173 35858
rect -61477 35238 -61173 35242
rect -60477 35858 -60173 35862
rect -60477 35242 -60473 35858
rect -60473 35242 -60177 35858
rect -60177 35242 -60173 35858
rect -60477 35238 -60173 35242
rect -59477 35858 -59173 35862
rect -59477 35242 -59473 35858
rect -59473 35242 -59177 35858
rect -59177 35242 -59173 35858
rect -59477 35238 -59173 35242
rect -74817 35198 -74513 35202
rect -74817 34902 -74813 35198
rect -74813 34902 -74517 35198
rect -74517 34902 -74513 35198
rect -74817 34898 -74513 34902
rect -74477 35198 -74173 35202
rect -74477 34902 -74473 35198
rect -74473 34902 -74177 35198
rect -74177 34902 -74173 35198
rect -74477 34898 -74173 34902
rect -74137 35198 -73513 35202
rect -74137 34902 -74133 35198
rect -74133 34902 -73517 35198
rect -73517 34902 -73513 35198
rect -74137 34898 -73513 34902
rect -73477 35198 -73173 35202
rect -73477 34902 -73473 35198
rect -73473 34902 -73177 35198
rect -73177 34902 -73173 35198
rect -73477 34898 -73173 34902
rect -73137 35198 -72513 35202
rect -73137 34902 -73133 35198
rect -73133 34902 -72517 35198
rect -72517 34902 -72513 35198
rect -73137 34898 -72513 34902
rect -72477 35198 -72173 35202
rect -72477 34902 -72473 35198
rect -72473 34902 -72177 35198
rect -72177 34902 -72173 35198
rect -72477 34898 -72173 34902
rect -72137 35198 -71513 35202
rect -72137 34902 -72133 35198
rect -72133 34902 -71517 35198
rect -71517 34902 -71513 35198
rect -72137 34898 -71513 34902
rect -71477 35198 -71173 35202
rect -71477 34902 -71473 35198
rect -71473 34902 -71177 35198
rect -71177 34902 -71173 35198
rect -71477 34898 -71173 34902
rect -71137 35198 -70513 35202
rect -71137 34902 -71133 35198
rect -71133 34902 -70517 35198
rect -70517 34902 -70513 35198
rect -71137 34898 -70513 34902
rect -70477 35198 -70173 35202
rect -70477 34902 -70473 35198
rect -70473 34902 -70177 35198
rect -70177 34902 -70173 35198
rect -70477 34898 -70173 34902
rect -70137 35198 -69513 35202
rect -70137 34902 -70133 35198
rect -70133 34902 -69517 35198
rect -69517 34902 -69513 35198
rect -70137 34898 -69513 34902
rect -69477 35198 -69173 35202
rect -69477 34902 -69473 35198
rect -69473 34902 -69177 35198
rect -69177 34902 -69173 35198
rect -69477 34898 -69173 34902
rect -69137 35198 -68513 35202
rect -69137 34902 -69133 35198
rect -69133 34902 -68517 35198
rect -68517 34902 -68513 35198
rect -69137 34898 -68513 34902
rect -68477 35198 -68173 35202
rect -68477 34902 -68473 35198
rect -68473 34902 -68177 35198
rect -68177 34902 -68173 35198
rect -68477 34898 -68173 34902
rect -68137 35198 -67513 35202
rect -68137 34902 -68133 35198
rect -68133 34902 -67517 35198
rect -67517 34902 -67513 35198
rect -68137 34898 -67513 34902
rect -67477 35198 -67173 35202
rect -67477 34902 -67473 35198
rect -67473 34902 -67177 35198
rect -67177 34902 -67173 35198
rect -67477 34898 -67173 34902
rect -67137 35198 -66513 35202
rect -67137 34902 -67133 35198
rect -67133 34902 -66517 35198
rect -66517 34902 -66513 35198
rect -67137 34898 -66513 34902
rect -66477 35198 -66173 35202
rect -66477 34902 -66473 35198
rect -66473 34902 -66177 35198
rect -66177 34902 -66173 35198
rect -66477 34898 -66173 34902
rect -66137 35198 -65513 35202
rect -66137 34902 -66133 35198
rect -66133 34902 -65517 35198
rect -65517 34902 -65513 35198
rect -66137 34898 -65513 34902
rect -65477 35198 -65173 35202
rect -65477 34902 -65473 35198
rect -65473 34902 -65177 35198
rect -65177 34902 -65173 35198
rect -65477 34898 -65173 34902
rect -65137 35198 -64513 35202
rect -65137 34902 -65133 35198
rect -65133 34902 -64517 35198
rect -64517 34902 -64513 35198
rect -65137 34898 -64513 34902
rect -64477 35198 -64173 35202
rect -64477 34902 -64473 35198
rect -64473 34902 -64177 35198
rect -64177 34902 -64173 35198
rect -64477 34898 -64173 34902
rect -64137 35198 -63513 35202
rect -64137 34902 -64133 35198
rect -64133 34902 -63517 35198
rect -63517 34902 -63513 35198
rect -64137 34898 -63513 34902
rect -63477 35198 -63173 35202
rect -63477 34902 -63473 35198
rect -63473 34902 -63177 35198
rect -63177 34902 -63173 35198
rect -63477 34898 -63173 34902
rect -63137 35198 -62513 35202
rect -63137 34902 -63133 35198
rect -63133 34902 -62517 35198
rect -62517 34902 -62513 35198
rect -63137 34898 -62513 34902
rect -62477 35198 -62173 35202
rect -62477 34902 -62473 35198
rect -62473 34902 -62177 35198
rect -62177 34902 -62173 35198
rect -62477 34898 -62173 34902
rect -62137 35198 -61513 35202
rect -62137 34902 -62133 35198
rect -62133 34902 -61517 35198
rect -61517 34902 -61513 35198
rect -62137 34898 -61513 34902
rect -61477 35198 -61173 35202
rect -61477 34902 -61473 35198
rect -61473 34902 -61177 35198
rect -61177 34902 -61173 35198
rect -61477 34898 -61173 34902
rect -61137 35198 -60513 35202
rect -61137 34902 -61133 35198
rect -61133 34902 -60517 35198
rect -60517 34902 -60513 35198
rect -61137 34898 -60513 34902
rect -60477 35198 -60173 35202
rect -60477 34902 -60473 35198
rect -60473 34902 -60177 35198
rect -60177 34902 -60173 35198
rect -60477 34898 -60173 34902
rect -60137 35198 -59513 35202
rect -60137 34902 -60133 35198
rect -60133 34902 -59517 35198
rect -59517 34902 -59513 35198
rect -60137 34898 -59513 34902
rect -59477 35198 -59173 35202
rect -59477 34902 -59473 35198
rect -59473 34902 -59177 35198
rect -59177 34902 -59173 35198
rect -59477 34898 -59173 34902
rect -59137 35198 -58833 35202
rect -59137 34902 -59133 35198
rect -59133 34902 -58837 35198
rect -58837 34902 -58833 35198
rect -59137 34898 -58833 34902
rect -74477 34858 -74173 34862
rect -74477 34242 -74473 34858
rect -74473 34242 -74177 34858
rect -74177 34242 -74173 34858
rect -74477 34238 -74173 34242
rect -73477 34858 -73173 34862
rect -73477 34242 -73473 34858
rect -73473 34242 -73177 34858
rect -73177 34242 -73173 34858
rect -73477 34238 -73173 34242
rect -72477 34858 -72173 34862
rect -72477 34242 -72473 34858
rect -72473 34242 -72177 34858
rect -72177 34242 -72173 34858
rect -72477 34238 -72173 34242
rect -71477 34858 -71173 34862
rect -71477 34242 -71473 34858
rect -71473 34242 -71177 34858
rect -71177 34242 -71173 34858
rect -71477 34238 -71173 34242
rect -70477 34858 -70173 34862
rect -70477 34242 -70473 34858
rect -70473 34242 -70177 34858
rect -70177 34242 -70173 34858
rect -70477 34238 -70173 34242
rect -69477 34858 -69173 34862
rect -69477 34242 -69473 34858
rect -69473 34242 -69177 34858
rect -69177 34242 -69173 34858
rect -69477 34238 -69173 34242
rect -68477 34858 -68173 34862
rect -68477 34242 -68473 34858
rect -68473 34242 -68177 34858
rect -68177 34242 -68173 34858
rect -68477 34238 -68173 34242
rect -67477 34858 -67173 34862
rect -67477 34242 -67473 34858
rect -67473 34242 -67177 34858
rect -67177 34242 -67173 34858
rect -67477 34238 -67173 34242
rect -66477 34858 -66173 34862
rect -66477 34242 -66473 34858
rect -66473 34242 -66177 34858
rect -66177 34242 -66173 34858
rect -66477 34238 -66173 34242
rect -65477 34858 -65173 34862
rect -65477 34242 -65473 34858
rect -65473 34242 -65177 34858
rect -65177 34242 -65173 34858
rect -65477 34238 -65173 34242
rect -64477 34858 -64173 34862
rect -64477 34242 -64473 34858
rect -64473 34242 -64177 34858
rect -64177 34242 -64173 34858
rect -64477 34238 -64173 34242
rect -63477 34858 -63173 34862
rect -63477 34242 -63473 34858
rect -63473 34242 -63177 34858
rect -63177 34242 -63173 34858
rect -63477 34238 -63173 34242
rect -62477 34858 -62173 34862
rect -62477 34242 -62473 34858
rect -62473 34242 -62177 34858
rect -62177 34242 -62173 34858
rect -62477 34238 -62173 34242
rect -61477 34858 -61173 34862
rect -61477 34242 -61473 34858
rect -61473 34242 -61177 34858
rect -61177 34242 -61173 34858
rect -61477 34238 -61173 34242
rect -60477 34858 -60173 34862
rect -60477 34242 -60473 34858
rect -60473 34242 -60177 34858
rect -60177 34242 -60173 34858
rect -60477 34238 -60173 34242
rect -59477 34858 -59173 34862
rect -59477 34242 -59473 34858
rect -59473 34242 -59177 34858
rect -59177 34242 -59173 34858
rect -59477 34238 -59173 34242
rect -74817 34198 -74513 34202
rect -74817 33902 -74813 34198
rect -74813 33902 -74517 34198
rect -74517 33902 -74513 34198
rect -74817 33898 -74513 33902
rect -74477 34198 -74173 34202
rect -74477 33902 -74473 34198
rect -74473 33902 -74177 34198
rect -74177 33902 -74173 34198
rect -74477 33898 -74173 33902
rect -74137 34198 -73513 34202
rect -74137 33902 -74133 34198
rect -74133 33902 -73517 34198
rect -73517 33902 -73513 34198
rect -74137 33898 -73513 33902
rect -73477 34198 -73173 34202
rect -73477 33902 -73473 34198
rect -73473 33902 -73177 34198
rect -73177 33902 -73173 34198
rect -73477 33898 -73173 33902
rect -73137 34198 -72513 34202
rect -73137 33902 -73133 34198
rect -73133 33902 -72517 34198
rect -72517 33902 -72513 34198
rect -73137 33898 -72513 33902
rect -72477 34198 -72173 34202
rect -72477 33902 -72473 34198
rect -72473 33902 -72177 34198
rect -72177 33902 -72173 34198
rect -72477 33898 -72173 33902
rect -72137 34198 -71513 34202
rect -72137 33902 -72133 34198
rect -72133 33902 -71517 34198
rect -71517 33902 -71513 34198
rect -72137 33898 -71513 33902
rect -71477 34198 -71173 34202
rect -71477 33902 -71473 34198
rect -71473 33902 -71177 34198
rect -71177 33902 -71173 34198
rect -71477 33898 -71173 33902
rect -71137 34198 -70513 34202
rect -71137 33902 -71133 34198
rect -71133 33902 -70517 34198
rect -70517 33902 -70513 34198
rect -71137 33898 -70513 33902
rect -70477 34198 -70173 34202
rect -70477 33902 -70473 34198
rect -70473 33902 -70177 34198
rect -70177 33902 -70173 34198
rect -70477 33898 -70173 33902
rect -70137 34198 -69513 34202
rect -70137 33902 -70133 34198
rect -70133 33902 -69517 34198
rect -69517 33902 -69513 34198
rect -70137 33898 -69513 33902
rect -69477 34198 -69173 34202
rect -69477 33902 -69473 34198
rect -69473 33902 -69177 34198
rect -69177 33902 -69173 34198
rect -69477 33898 -69173 33902
rect -69137 34198 -68513 34202
rect -69137 33902 -69133 34198
rect -69133 33902 -68517 34198
rect -68517 33902 -68513 34198
rect -69137 33898 -68513 33902
rect -68477 34198 -68173 34202
rect -68477 33902 -68473 34198
rect -68473 33902 -68177 34198
rect -68177 33902 -68173 34198
rect -68477 33898 -68173 33902
rect -68137 34198 -67513 34202
rect -68137 33902 -68133 34198
rect -68133 33902 -67517 34198
rect -67517 33902 -67513 34198
rect -68137 33898 -67513 33902
rect -67477 34198 -67173 34202
rect -67477 33902 -67473 34198
rect -67473 33902 -67177 34198
rect -67177 33902 -67173 34198
rect -67477 33898 -67173 33902
rect -67137 34198 -66513 34202
rect -67137 33902 -67133 34198
rect -67133 33902 -66517 34198
rect -66517 33902 -66513 34198
rect -67137 33898 -66513 33902
rect -66477 34198 -66173 34202
rect -66477 33902 -66473 34198
rect -66473 33902 -66177 34198
rect -66177 33902 -66173 34198
rect -66477 33898 -66173 33902
rect -66137 34198 -65513 34202
rect -66137 33902 -66133 34198
rect -66133 33902 -65517 34198
rect -65517 33902 -65513 34198
rect -66137 33898 -65513 33902
rect -65477 34198 -65173 34202
rect -65477 33902 -65473 34198
rect -65473 33902 -65177 34198
rect -65177 33902 -65173 34198
rect -65477 33898 -65173 33902
rect -65137 34198 -64513 34202
rect -65137 33902 -65133 34198
rect -65133 33902 -64517 34198
rect -64517 33902 -64513 34198
rect -65137 33898 -64513 33902
rect -64477 34198 -64173 34202
rect -64477 33902 -64473 34198
rect -64473 33902 -64177 34198
rect -64177 33902 -64173 34198
rect -64477 33898 -64173 33902
rect -64137 34198 -63513 34202
rect -64137 33902 -64133 34198
rect -64133 33902 -63517 34198
rect -63517 33902 -63513 34198
rect -64137 33898 -63513 33902
rect -63477 34198 -63173 34202
rect -63477 33902 -63473 34198
rect -63473 33902 -63177 34198
rect -63177 33902 -63173 34198
rect -63477 33898 -63173 33902
rect -63137 34198 -62513 34202
rect -63137 33902 -63133 34198
rect -63133 33902 -62517 34198
rect -62517 33902 -62513 34198
rect -63137 33898 -62513 33902
rect -62477 34198 -62173 34202
rect -62477 33902 -62473 34198
rect -62473 33902 -62177 34198
rect -62177 33902 -62173 34198
rect -62477 33898 -62173 33902
rect -62137 34198 -61513 34202
rect -62137 33902 -62133 34198
rect -62133 33902 -61517 34198
rect -61517 33902 -61513 34198
rect -62137 33898 -61513 33902
rect -61477 34198 -61173 34202
rect -61477 33902 -61473 34198
rect -61473 33902 -61177 34198
rect -61177 33902 -61173 34198
rect -61477 33898 -61173 33902
rect -61137 34198 -60513 34202
rect -61137 33902 -61133 34198
rect -61133 33902 -60517 34198
rect -60517 33902 -60513 34198
rect -61137 33898 -60513 33902
rect -60477 34198 -60173 34202
rect -60477 33902 -60473 34198
rect -60473 33902 -60177 34198
rect -60177 33902 -60173 34198
rect -60477 33898 -60173 33902
rect -60137 34198 -59513 34202
rect -60137 33902 -60133 34198
rect -60133 33902 -59517 34198
rect -59517 33902 -59513 34198
rect -60137 33898 -59513 33902
rect -59477 34198 -59173 34202
rect -59477 33902 -59473 34198
rect -59473 33902 -59177 34198
rect -59177 33902 -59173 34198
rect -59477 33898 -59173 33902
rect -59137 34198 -58833 34202
rect -59137 33902 -59133 34198
rect -59133 33902 -58837 34198
rect -58837 33902 -58833 34198
rect -59137 33898 -58833 33902
rect -74477 33858 -74173 33862
rect -74477 33242 -74473 33858
rect -74473 33242 -74177 33858
rect -74177 33242 -74173 33858
rect -74477 33238 -74173 33242
rect -73477 33858 -73173 33862
rect -73477 33242 -73473 33858
rect -73473 33242 -73177 33858
rect -73177 33242 -73173 33858
rect -73477 33238 -73173 33242
rect -72477 33858 -72173 33862
rect -72477 33242 -72473 33858
rect -72473 33242 -72177 33858
rect -72177 33242 -72173 33858
rect -72477 33238 -72173 33242
rect -71477 33858 -71173 33862
rect -71477 33242 -71473 33858
rect -71473 33242 -71177 33858
rect -71177 33242 -71173 33858
rect -71477 33238 -71173 33242
rect -70477 33858 -70173 33862
rect -70477 33242 -70473 33858
rect -70473 33242 -70177 33858
rect -70177 33242 -70173 33858
rect -70477 33238 -70173 33242
rect -69477 33858 -69173 33862
rect -69477 33242 -69473 33858
rect -69473 33242 -69177 33858
rect -69177 33242 -69173 33858
rect -69477 33238 -69173 33242
rect -68477 33858 -68173 33862
rect -68477 33242 -68473 33858
rect -68473 33242 -68177 33858
rect -68177 33242 -68173 33858
rect -68477 33238 -68173 33242
rect -67477 33858 -67173 33862
rect -67477 33242 -67473 33858
rect -67473 33242 -67177 33858
rect -67177 33242 -67173 33858
rect -67477 33238 -67173 33242
rect -66477 33858 -66173 33862
rect -66477 33242 -66473 33858
rect -66473 33242 -66177 33858
rect -66177 33242 -66173 33858
rect -66477 33238 -66173 33242
rect -65477 33858 -65173 33862
rect -65477 33242 -65473 33858
rect -65473 33242 -65177 33858
rect -65177 33242 -65173 33858
rect -65477 33238 -65173 33242
rect -64477 33858 -64173 33862
rect -64477 33242 -64473 33858
rect -64473 33242 -64177 33858
rect -64177 33242 -64173 33858
rect -64477 33238 -64173 33242
rect -63477 33858 -63173 33862
rect -63477 33242 -63473 33858
rect -63473 33242 -63177 33858
rect -63177 33242 -63173 33858
rect -63477 33238 -63173 33242
rect -62477 33858 -62173 33862
rect -62477 33242 -62473 33858
rect -62473 33242 -62177 33858
rect -62177 33242 -62173 33858
rect -62477 33238 -62173 33242
rect -61477 33858 -61173 33862
rect -61477 33242 -61473 33858
rect -61473 33242 -61177 33858
rect -61177 33242 -61173 33858
rect -61477 33238 -61173 33242
rect -60477 33858 -60173 33862
rect -60477 33242 -60473 33858
rect -60473 33242 -60177 33858
rect -60177 33242 -60173 33858
rect -60477 33238 -60173 33242
rect -59477 33858 -59173 33862
rect -59477 33242 -59473 33858
rect -59473 33242 -59177 33858
rect -59177 33242 -59173 33858
rect -59477 33238 -59173 33242
rect -74817 33198 -74513 33202
rect -74817 32902 -74813 33198
rect -74813 32902 -74517 33198
rect -74517 32902 -74513 33198
rect -74817 32898 -74513 32902
rect -74477 33198 -74173 33202
rect -74477 32902 -74473 33198
rect -74473 32902 -74177 33198
rect -74177 32902 -74173 33198
rect -74477 32898 -74173 32902
rect -74137 33198 -73513 33202
rect -74137 32902 -74133 33198
rect -74133 32902 -73517 33198
rect -73517 32902 -73513 33198
rect -74137 32898 -73513 32902
rect -73477 33198 -73173 33202
rect -73477 32902 -73473 33198
rect -73473 32902 -73177 33198
rect -73177 32902 -73173 33198
rect -73477 32898 -73173 32902
rect -73137 33198 -72513 33202
rect -73137 32902 -73133 33198
rect -73133 32902 -72517 33198
rect -72517 32902 -72513 33198
rect -73137 32898 -72513 32902
rect -72477 33198 -72173 33202
rect -72477 32902 -72473 33198
rect -72473 32902 -72177 33198
rect -72177 32902 -72173 33198
rect -72477 32898 -72173 32902
rect -72137 33198 -71513 33202
rect -72137 32902 -72133 33198
rect -72133 32902 -71517 33198
rect -71517 32902 -71513 33198
rect -72137 32898 -71513 32902
rect -71477 33198 -71173 33202
rect -71477 32902 -71473 33198
rect -71473 32902 -71177 33198
rect -71177 32902 -71173 33198
rect -71477 32898 -71173 32902
rect -71137 33198 -70513 33202
rect -71137 32902 -71133 33198
rect -71133 32902 -70517 33198
rect -70517 32902 -70513 33198
rect -71137 32898 -70513 32902
rect -70477 33198 -70173 33202
rect -70477 32902 -70473 33198
rect -70473 32902 -70177 33198
rect -70177 32902 -70173 33198
rect -70477 32898 -70173 32902
rect -70137 33198 -69513 33202
rect -70137 32902 -70133 33198
rect -70133 32902 -69517 33198
rect -69517 32902 -69513 33198
rect -70137 32898 -69513 32902
rect -69477 33198 -69173 33202
rect -69477 32902 -69473 33198
rect -69473 32902 -69177 33198
rect -69177 32902 -69173 33198
rect -69477 32898 -69173 32902
rect -69137 33198 -68513 33202
rect -69137 32902 -69133 33198
rect -69133 32902 -68517 33198
rect -68517 32902 -68513 33198
rect -69137 32898 -68513 32902
rect -68477 33198 -68173 33202
rect -68477 32902 -68473 33198
rect -68473 32902 -68177 33198
rect -68177 32902 -68173 33198
rect -68477 32898 -68173 32902
rect -68137 33198 -67513 33202
rect -68137 32902 -68133 33198
rect -68133 32902 -67517 33198
rect -67517 32902 -67513 33198
rect -68137 32898 -67513 32902
rect -67477 33198 -67173 33202
rect -67477 32902 -67473 33198
rect -67473 32902 -67177 33198
rect -67177 32902 -67173 33198
rect -67477 32898 -67173 32902
rect -67137 33198 -66513 33202
rect -67137 32902 -67133 33198
rect -67133 32902 -66517 33198
rect -66517 32902 -66513 33198
rect -67137 32898 -66513 32902
rect -66477 33198 -66173 33202
rect -66477 32902 -66473 33198
rect -66473 32902 -66177 33198
rect -66177 32902 -66173 33198
rect -66477 32898 -66173 32902
rect -66137 33198 -65513 33202
rect -66137 32902 -66133 33198
rect -66133 32902 -65517 33198
rect -65517 32902 -65513 33198
rect -66137 32898 -65513 32902
rect -65477 33198 -65173 33202
rect -65477 32902 -65473 33198
rect -65473 32902 -65177 33198
rect -65177 32902 -65173 33198
rect -65477 32898 -65173 32902
rect -65137 33198 -64513 33202
rect -65137 32902 -65133 33198
rect -65133 32902 -64517 33198
rect -64517 32902 -64513 33198
rect -65137 32898 -64513 32902
rect -64477 33198 -64173 33202
rect -64477 32902 -64473 33198
rect -64473 32902 -64177 33198
rect -64177 32902 -64173 33198
rect -64477 32898 -64173 32902
rect -64137 33198 -63513 33202
rect -64137 32902 -64133 33198
rect -64133 32902 -63517 33198
rect -63517 32902 -63513 33198
rect -64137 32898 -63513 32902
rect -63477 33198 -63173 33202
rect -63477 32902 -63473 33198
rect -63473 32902 -63177 33198
rect -63177 32902 -63173 33198
rect -63477 32898 -63173 32902
rect -63137 33198 -62513 33202
rect -63137 32902 -63133 33198
rect -63133 32902 -62517 33198
rect -62517 32902 -62513 33198
rect -63137 32898 -62513 32902
rect -62477 33198 -62173 33202
rect -62477 32902 -62473 33198
rect -62473 32902 -62177 33198
rect -62177 32902 -62173 33198
rect -62477 32898 -62173 32902
rect -62137 33198 -61513 33202
rect -62137 32902 -62133 33198
rect -62133 32902 -61517 33198
rect -61517 32902 -61513 33198
rect -62137 32898 -61513 32902
rect -61477 33198 -61173 33202
rect -61477 32902 -61473 33198
rect -61473 32902 -61177 33198
rect -61177 32902 -61173 33198
rect -61477 32898 -61173 32902
rect -61137 33198 -60513 33202
rect -61137 32902 -61133 33198
rect -61133 32902 -60517 33198
rect -60517 32902 -60513 33198
rect -61137 32898 -60513 32902
rect -60477 33198 -60173 33202
rect -60477 32902 -60473 33198
rect -60473 32902 -60177 33198
rect -60177 32902 -60173 33198
rect -60477 32898 -60173 32902
rect -60137 33198 -59513 33202
rect -60137 32902 -60133 33198
rect -60133 32902 -59517 33198
rect -59517 32902 -59513 33198
rect -60137 32898 -59513 32902
rect -59477 33198 -59173 33202
rect -59477 32902 -59473 33198
rect -59473 32902 -59177 33198
rect -59177 32902 -59173 33198
rect -59477 32898 -59173 32902
rect -59137 33198 -58833 33202
rect -59137 32902 -59133 33198
rect -59133 32902 -58837 33198
rect -58837 32902 -58833 33198
rect -59137 32898 -58833 32902
rect 10002 38538 10306 38542
rect 10002 38242 10006 38538
rect 10006 38242 10302 38538
rect 10302 38242 10306 38538
rect 10002 38238 10306 38242
rect 11002 38538 11306 38542
rect 11002 38242 11006 38538
rect 11006 38242 11302 38538
rect 11302 38242 11306 38538
rect 11002 38238 11306 38242
rect 12002 38538 12306 38542
rect 12002 38242 12006 38538
rect 12006 38242 12302 38538
rect 12302 38242 12306 38538
rect 12002 38238 12306 38242
rect 13002 38538 13306 38542
rect 13002 38242 13006 38538
rect 13006 38242 13302 38538
rect 13302 38242 13306 38538
rect 13002 38238 13306 38242
rect 14002 38538 14306 38542
rect 14002 38242 14006 38538
rect 14006 38242 14302 38538
rect 14302 38242 14306 38538
rect 14002 38238 14306 38242
rect 15002 38538 15306 38542
rect 15002 38242 15006 38538
rect 15006 38242 15302 38538
rect 15302 38242 15306 38538
rect 15002 38238 15306 38242
rect 16002 38538 16306 38542
rect 16002 38242 16006 38538
rect 16006 38242 16302 38538
rect 16302 38242 16306 38538
rect 16002 38238 16306 38242
rect 17002 38538 17306 38542
rect 17002 38242 17006 38538
rect 17006 38242 17302 38538
rect 17302 38242 17306 38538
rect 17002 38238 17306 38242
rect 18002 38538 18306 38542
rect 18002 38242 18006 38538
rect 18006 38242 18302 38538
rect 18302 38242 18306 38538
rect 18002 38238 18306 38242
rect 19002 38538 19306 38542
rect 19002 38242 19006 38538
rect 19006 38242 19302 38538
rect 19302 38242 19306 38538
rect 19002 38238 19306 38242
rect 20002 38538 20306 38542
rect 20002 38242 20006 38538
rect 20006 38242 20302 38538
rect 20302 38242 20306 38538
rect 20002 38238 20306 38242
rect 21002 38538 21306 38542
rect 21002 38242 21006 38538
rect 21006 38242 21302 38538
rect 21302 38242 21306 38538
rect 21002 38238 21306 38242
rect 22002 38538 22306 38542
rect 22002 38242 22006 38538
rect 22006 38242 22302 38538
rect 22302 38242 22306 38538
rect 22002 38238 22306 38242
rect 23002 38538 23306 38542
rect 23002 38242 23006 38538
rect 23006 38242 23302 38538
rect 23302 38242 23306 38538
rect 23002 38238 23306 38242
rect 24002 38538 24306 38542
rect 24002 38242 24006 38538
rect 24006 38242 24302 38538
rect 24302 38242 24306 38538
rect 24002 38238 24306 38242
rect 25002 38538 25306 38542
rect 25002 38242 25006 38538
rect 25006 38242 25302 38538
rect 25302 38242 25306 38538
rect 25002 38238 25306 38242
rect 26002 38538 26306 38542
rect 26002 38242 26006 38538
rect 26006 38242 26302 38538
rect 26302 38242 26306 38538
rect 26002 38238 26306 38242
rect 27002 38538 27306 38542
rect 27002 38242 27006 38538
rect 27006 38242 27302 38538
rect 27302 38242 27306 38538
rect 27002 38238 27306 38242
rect 28002 38538 28306 38542
rect 28002 38242 28006 38538
rect 28006 38242 28302 38538
rect 28302 38242 28306 38538
rect 28002 38238 28306 38242
rect 29002 38538 29306 38542
rect 29002 38242 29006 38538
rect 29006 38242 29302 38538
rect 29302 38242 29306 38538
rect 29002 38238 29306 38242
rect 30002 38538 30306 38542
rect 30002 38242 30006 38538
rect 30006 38242 30302 38538
rect 30302 38242 30306 38538
rect 30002 38238 30306 38242
rect 31002 38538 31306 38542
rect 31002 38242 31006 38538
rect 31006 38242 31302 38538
rect 31302 38242 31306 38538
rect 31002 38238 31306 38242
rect 32002 38538 32306 38542
rect 32002 38242 32006 38538
rect 32006 38242 32302 38538
rect 32302 38242 32306 38538
rect 32002 38238 32306 38242
rect 33002 38538 33306 38542
rect 33002 38242 33006 38538
rect 33006 38242 33302 38538
rect 33302 38242 33306 38538
rect 33002 38238 33306 38242
rect 34002 38538 34306 38542
rect 34002 38242 34006 38538
rect 34006 38242 34302 38538
rect 34302 38242 34306 38538
rect 34002 38238 34306 38242
rect 9662 38198 9966 38202
rect 9662 37902 9666 38198
rect 9666 37902 9962 38198
rect 9962 37902 9966 38198
rect 9662 37898 9966 37902
rect 10002 38198 10306 38202
rect 10002 37902 10006 38198
rect 10006 37902 10302 38198
rect 10302 37902 10306 38198
rect 10002 37898 10306 37902
rect 10342 38198 10966 38202
rect 10342 37902 10346 38198
rect 10346 37902 10962 38198
rect 10962 37902 10966 38198
rect 10342 37898 10966 37902
rect 11002 38198 11306 38202
rect 11002 37902 11006 38198
rect 11006 37902 11302 38198
rect 11302 37902 11306 38198
rect 11002 37898 11306 37902
rect 11342 38198 11966 38202
rect 11342 37902 11346 38198
rect 11346 37902 11962 38198
rect 11962 37902 11966 38198
rect 11342 37898 11966 37902
rect 12002 38198 12306 38202
rect 12002 37902 12006 38198
rect 12006 37902 12302 38198
rect 12302 37902 12306 38198
rect 12002 37898 12306 37902
rect 12342 38198 12966 38202
rect 12342 37902 12346 38198
rect 12346 37902 12962 38198
rect 12962 37902 12966 38198
rect 12342 37898 12966 37902
rect 13002 38198 13306 38202
rect 13002 37902 13006 38198
rect 13006 37902 13302 38198
rect 13302 37902 13306 38198
rect 13002 37898 13306 37902
rect 13342 38198 13966 38202
rect 13342 37902 13346 38198
rect 13346 37902 13962 38198
rect 13962 37902 13966 38198
rect 13342 37898 13966 37902
rect 14002 38198 14306 38202
rect 14002 37902 14006 38198
rect 14006 37902 14302 38198
rect 14302 37902 14306 38198
rect 14002 37898 14306 37902
rect 14342 38198 14966 38202
rect 14342 37902 14346 38198
rect 14346 37902 14962 38198
rect 14962 37902 14966 38198
rect 14342 37898 14966 37902
rect 15002 38198 15306 38202
rect 15002 37902 15006 38198
rect 15006 37902 15302 38198
rect 15302 37902 15306 38198
rect 15002 37898 15306 37902
rect 15342 38198 15966 38202
rect 15342 37902 15346 38198
rect 15346 37902 15962 38198
rect 15962 37902 15966 38198
rect 15342 37898 15966 37902
rect 16002 38198 16306 38202
rect 16002 37902 16006 38198
rect 16006 37902 16302 38198
rect 16302 37902 16306 38198
rect 16002 37898 16306 37902
rect 16342 38198 16966 38202
rect 16342 37902 16346 38198
rect 16346 37902 16962 38198
rect 16962 37902 16966 38198
rect 16342 37898 16966 37902
rect 17002 38198 17306 38202
rect 17002 37902 17006 38198
rect 17006 37902 17302 38198
rect 17302 37902 17306 38198
rect 17002 37898 17306 37902
rect 17342 38198 17966 38202
rect 17342 37902 17346 38198
rect 17346 37902 17962 38198
rect 17962 37902 17966 38198
rect 17342 37898 17966 37902
rect 18002 38198 18306 38202
rect 18002 37902 18006 38198
rect 18006 37902 18302 38198
rect 18302 37902 18306 38198
rect 18002 37898 18306 37902
rect 18342 38198 18966 38202
rect 18342 37902 18346 38198
rect 18346 37902 18962 38198
rect 18962 37902 18966 38198
rect 18342 37898 18966 37902
rect 19002 38198 19306 38202
rect 19002 37902 19006 38198
rect 19006 37902 19302 38198
rect 19302 37902 19306 38198
rect 19002 37898 19306 37902
rect 19342 38198 19966 38202
rect 19342 37902 19346 38198
rect 19346 37902 19962 38198
rect 19962 37902 19966 38198
rect 19342 37898 19966 37902
rect 20002 38198 20306 38202
rect 20002 37902 20006 38198
rect 20006 37902 20302 38198
rect 20302 37902 20306 38198
rect 20002 37898 20306 37902
rect 20342 38198 20966 38202
rect 20342 37902 20346 38198
rect 20346 37902 20962 38198
rect 20962 37902 20966 38198
rect 20342 37898 20966 37902
rect 21002 38198 21306 38202
rect 21002 37902 21006 38198
rect 21006 37902 21302 38198
rect 21302 37902 21306 38198
rect 21002 37898 21306 37902
rect 21342 38198 21966 38202
rect 21342 37902 21346 38198
rect 21346 37902 21962 38198
rect 21962 37902 21966 38198
rect 21342 37898 21966 37902
rect 22002 38198 22306 38202
rect 22002 37902 22006 38198
rect 22006 37902 22302 38198
rect 22302 37902 22306 38198
rect 22002 37898 22306 37902
rect 22342 38198 22966 38202
rect 22342 37902 22346 38198
rect 22346 37902 22962 38198
rect 22962 37902 22966 38198
rect 22342 37898 22966 37902
rect 23002 38198 23306 38202
rect 23002 37902 23006 38198
rect 23006 37902 23302 38198
rect 23302 37902 23306 38198
rect 23002 37898 23306 37902
rect 23342 38198 23966 38202
rect 23342 37902 23346 38198
rect 23346 37902 23962 38198
rect 23962 37902 23966 38198
rect 23342 37898 23966 37902
rect 24002 38198 24306 38202
rect 24002 37902 24006 38198
rect 24006 37902 24302 38198
rect 24302 37902 24306 38198
rect 24002 37898 24306 37902
rect 24342 38198 24966 38202
rect 24342 37902 24346 38198
rect 24346 37902 24962 38198
rect 24962 37902 24966 38198
rect 24342 37898 24966 37902
rect 25002 38198 25306 38202
rect 25002 37902 25006 38198
rect 25006 37902 25302 38198
rect 25302 37902 25306 38198
rect 25002 37898 25306 37902
rect 25342 38198 25966 38202
rect 25342 37902 25346 38198
rect 25346 37902 25962 38198
rect 25962 37902 25966 38198
rect 25342 37898 25966 37902
rect 26002 38198 26306 38202
rect 26002 37902 26006 38198
rect 26006 37902 26302 38198
rect 26302 37902 26306 38198
rect 26002 37898 26306 37902
rect 26342 38198 26966 38202
rect 26342 37902 26346 38198
rect 26346 37902 26962 38198
rect 26962 37902 26966 38198
rect 26342 37898 26966 37902
rect 27002 38198 27306 38202
rect 27002 37902 27006 38198
rect 27006 37902 27302 38198
rect 27302 37902 27306 38198
rect 27002 37898 27306 37902
rect 27342 38198 27966 38202
rect 27342 37902 27346 38198
rect 27346 37902 27962 38198
rect 27962 37902 27966 38198
rect 27342 37898 27966 37902
rect 28002 38198 28306 38202
rect 28002 37902 28006 38198
rect 28006 37902 28302 38198
rect 28302 37902 28306 38198
rect 28002 37898 28306 37902
rect 28342 38198 28966 38202
rect 28342 37902 28346 38198
rect 28346 37902 28962 38198
rect 28962 37902 28966 38198
rect 28342 37898 28966 37902
rect 29002 38198 29306 38202
rect 29002 37902 29006 38198
rect 29006 37902 29302 38198
rect 29302 37902 29306 38198
rect 29002 37898 29306 37902
rect 29342 38198 29966 38202
rect 29342 37902 29346 38198
rect 29346 37902 29962 38198
rect 29962 37902 29966 38198
rect 29342 37898 29966 37902
rect 30002 38198 30306 38202
rect 30002 37902 30006 38198
rect 30006 37902 30302 38198
rect 30302 37902 30306 38198
rect 30002 37898 30306 37902
rect 30342 38198 30966 38202
rect 30342 37902 30346 38198
rect 30346 37902 30962 38198
rect 30962 37902 30966 38198
rect 30342 37898 30966 37902
rect 31002 38198 31306 38202
rect 31002 37902 31006 38198
rect 31006 37902 31302 38198
rect 31302 37902 31306 38198
rect 31002 37898 31306 37902
rect 31342 38198 31966 38202
rect 31342 37902 31346 38198
rect 31346 37902 31962 38198
rect 31962 37902 31966 38198
rect 31342 37898 31966 37902
rect 32002 38198 32306 38202
rect 32002 37902 32006 38198
rect 32006 37902 32302 38198
rect 32302 37902 32306 38198
rect 32002 37898 32306 37902
rect 32342 38198 32966 38202
rect 32342 37902 32346 38198
rect 32346 37902 32962 38198
rect 32962 37902 32966 38198
rect 32342 37898 32966 37902
rect 33002 38198 33306 38202
rect 33002 37902 33006 38198
rect 33006 37902 33302 38198
rect 33302 37902 33306 38198
rect 33002 37898 33306 37902
rect 33342 38198 33966 38202
rect 33342 37902 33346 38198
rect 33346 37902 33962 38198
rect 33962 37902 33966 38198
rect 33342 37898 33966 37902
rect 34002 38198 34306 38202
rect 34002 37902 34006 38198
rect 34006 37902 34302 38198
rect 34302 37902 34306 38198
rect 34002 37898 34306 37902
rect 34342 38198 34646 38202
rect 34342 37902 34346 38198
rect 34346 37902 34642 38198
rect 34642 37902 34646 38198
rect 34342 37898 34646 37902
rect 10002 37858 10306 37862
rect 10002 37242 10006 37858
rect 10006 37242 10302 37858
rect 10302 37242 10306 37858
rect 10002 37238 10306 37242
rect 11002 37858 11306 37862
rect 11002 37242 11006 37858
rect 11006 37242 11302 37858
rect 11302 37242 11306 37858
rect 11002 37238 11306 37242
rect 12002 37858 12306 37862
rect 12002 37242 12006 37858
rect 12006 37242 12302 37858
rect 12302 37242 12306 37858
rect 12002 37238 12306 37242
rect 13002 37858 13306 37862
rect 13002 37242 13006 37858
rect 13006 37242 13302 37858
rect 13302 37242 13306 37858
rect 13002 37238 13306 37242
rect 14002 37858 14306 37862
rect 14002 37242 14006 37858
rect 14006 37242 14302 37858
rect 14302 37242 14306 37858
rect 14002 37238 14306 37242
rect 15002 37858 15306 37862
rect 15002 37242 15006 37858
rect 15006 37242 15302 37858
rect 15302 37242 15306 37858
rect 15002 37238 15306 37242
rect 16002 37858 16306 37862
rect 16002 37242 16006 37858
rect 16006 37242 16302 37858
rect 16302 37242 16306 37858
rect 16002 37238 16306 37242
rect 17002 37858 17306 37862
rect 17002 37242 17006 37858
rect 17006 37242 17302 37858
rect 17302 37242 17306 37858
rect 17002 37238 17306 37242
rect 18002 37858 18306 37862
rect 18002 37242 18006 37858
rect 18006 37242 18302 37858
rect 18302 37242 18306 37858
rect 18002 37238 18306 37242
rect 19002 37858 19306 37862
rect 19002 37242 19006 37858
rect 19006 37242 19302 37858
rect 19302 37242 19306 37858
rect 19002 37238 19306 37242
rect 20002 37858 20306 37862
rect 20002 37242 20006 37858
rect 20006 37242 20302 37858
rect 20302 37242 20306 37858
rect 20002 37238 20306 37242
rect 21002 37858 21306 37862
rect 21002 37242 21006 37858
rect 21006 37242 21302 37858
rect 21302 37242 21306 37858
rect 21002 37238 21306 37242
rect 22002 37858 22306 37862
rect 22002 37242 22006 37858
rect 22006 37242 22302 37858
rect 22302 37242 22306 37858
rect 22002 37238 22306 37242
rect 23002 37858 23306 37862
rect 23002 37242 23006 37858
rect 23006 37242 23302 37858
rect 23302 37242 23306 37858
rect 23002 37238 23306 37242
rect 24002 37858 24306 37862
rect 24002 37242 24006 37858
rect 24006 37242 24302 37858
rect 24302 37242 24306 37858
rect 24002 37238 24306 37242
rect 25002 37858 25306 37862
rect 25002 37242 25006 37858
rect 25006 37242 25302 37858
rect 25302 37242 25306 37858
rect 25002 37238 25306 37242
rect 26002 37858 26306 37862
rect 26002 37242 26006 37858
rect 26006 37242 26302 37858
rect 26302 37242 26306 37858
rect 26002 37238 26306 37242
rect 27002 37858 27306 37862
rect 27002 37242 27006 37858
rect 27006 37242 27302 37858
rect 27302 37242 27306 37858
rect 27002 37238 27306 37242
rect 28002 37858 28306 37862
rect 28002 37242 28006 37858
rect 28006 37242 28302 37858
rect 28302 37242 28306 37858
rect 28002 37238 28306 37242
rect 29002 37858 29306 37862
rect 29002 37242 29006 37858
rect 29006 37242 29302 37858
rect 29302 37242 29306 37858
rect 29002 37238 29306 37242
rect 30002 37858 30306 37862
rect 30002 37242 30006 37858
rect 30006 37242 30302 37858
rect 30302 37242 30306 37858
rect 30002 37238 30306 37242
rect 31002 37858 31306 37862
rect 31002 37242 31006 37858
rect 31006 37242 31302 37858
rect 31302 37242 31306 37858
rect 31002 37238 31306 37242
rect 32002 37858 32306 37862
rect 32002 37242 32006 37858
rect 32006 37242 32302 37858
rect 32302 37242 32306 37858
rect 32002 37238 32306 37242
rect 33002 37858 33306 37862
rect 33002 37242 33006 37858
rect 33006 37242 33302 37858
rect 33302 37242 33306 37858
rect 33002 37238 33306 37242
rect 34002 37858 34306 37862
rect 34002 37242 34006 37858
rect 34006 37242 34302 37858
rect 34302 37242 34306 37858
rect 34002 37238 34306 37242
rect 9662 37198 9966 37202
rect 9662 36902 9666 37198
rect 9666 36902 9962 37198
rect 9962 36902 9966 37198
rect 9662 36898 9966 36902
rect 10002 37198 10306 37202
rect 10002 36902 10006 37198
rect 10006 36902 10302 37198
rect 10302 36902 10306 37198
rect 10002 36898 10306 36902
rect 10342 37198 10966 37202
rect 10342 36902 10346 37198
rect 10346 36902 10962 37198
rect 10962 36902 10966 37198
rect 10342 36898 10966 36902
rect 11002 37198 11306 37202
rect 11002 36902 11006 37198
rect 11006 36902 11302 37198
rect 11302 36902 11306 37198
rect 11002 36898 11306 36902
rect 11342 37198 11966 37202
rect 11342 36902 11346 37198
rect 11346 36902 11962 37198
rect 11962 36902 11966 37198
rect 11342 36898 11966 36902
rect 12002 37198 12306 37202
rect 12002 36902 12006 37198
rect 12006 36902 12302 37198
rect 12302 36902 12306 37198
rect 12002 36898 12306 36902
rect 12342 37198 12966 37202
rect 12342 36902 12346 37198
rect 12346 36902 12962 37198
rect 12962 36902 12966 37198
rect 12342 36898 12966 36902
rect 13002 37198 13306 37202
rect 13002 36902 13006 37198
rect 13006 36902 13302 37198
rect 13302 36902 13306 37198
rect 13002 36898 13306 36902
rect 13342 37198 13966 37202
rect 13342 36902 13346 37198
rect 13346 36902 13962 37198
rect 13962 36902 13966 37198
rect 13342 36898 13966 36902
rect 14002 37198 14306 37202
rect 14002 36902 14006 37198
rect 14006 36902 14302 37198
rect 14302 36902 14306 37198
rect 14002 36898 14306 36902
rect 14342 37198 14966 37202
rect 14342 36902 14346 37198
rect 14346 36902 14962 37198
rect 14962 36902 14966 37198
rect 14342 36898 14966 36902
rect 15002 37198 15306 37202
rect 15002 36902 15006 37198
rect 15006 36902 15302 37198
rect 15302 36902 15306 37198
rect 15002 36898 15306 36902
rect 15342 37198 15966 37202
rect 15342 36902 15346 37198
rect 15346 36902 15962 37198
rect 15962 36902 15966 37198
rect 15342 36898 15966 36902
rect 16002 37198 16306 37202
rect 16002 36902 16006 37198
rect 16006 36902 16302 37198
rect 16302 36902 16306 37198
rect 16002 36898 16306 36902
rect 16342 37198 16966 37202
rect 16342 36902 16346 37198
rect 16346 36902 16962 37198
rect 16962 36902 16966 37198
rect 16342 36898 16966 36902
rect 17002 37198 17306 37202
rect 17002 36902 17006 37198
rect 17006 36902 17302 37198
rect 17302 36902 17306 37198
rect 17002 36898 17306 36902
rect 17342 37198 17966 37202
rect 17342 36902 17346 37198
rect 17346 36902 17962 37198
rect 17962 36902 17966 37198
rect 17342 36898 17966 36902
rect 18002 37198 18306 37202
rect 18002 36902 18006 37198
rect 18006 36902 18302 37198
rect 18302 36902 18306 37198
rect 18002 36898 18306 36902
rect 18342 37198 18966 37202
rect 18342 36902 18346 37198
rect 18346 36902 18962 37198
rect 18962 36902 18966 37198
rect 18342 36898 18966 36902
rect 19002 37198 19306 37202
rect 19002 36902 19006 37198
rect 19006 36902 19302 37198
rect 19302 36902 19306 37198
rect 19002 36898 19306 36902
rect 19342 37198 19966 37202
rect 19342 36902 19346 37198
rect 19346 36902 19962 37198
rect 19962 36902 19966 37198
rect 19342 36898 19966 36902
rect 20002 37198 20306 37202
rect 20002 36902 20006 37198
rect 20006 36902 20302 37198
rect 20302 36902 20306 37198
rect 20002 36898 20306 36902
rect 20342 37198 20966 37202
rect 20342 36902 20346 37198
rect 20346 36902 20962 37198
rect 20962 36902 20966 37198
rect 20342 36898 20966 36902
rect 21002 37198 21306 37202
rect 21002 36902 21006 37198
rect 21006 36902 21302 37198
rect 21302 36902 21306 37198
rect 21002 36898 21306 36902
rect 21342 37198 21966 37202
rect 21342 36902 21346 37198
rect 21346 36902 21962 37198
rect 21962 36902 21966 37198
rect 21342 36898 21966 36902
rect 22002 37198 22306 37202
rect 22002 36902 22006 37198
rect 22006 36902 22302 37198
rect 22302 36902 22306 37198
rect 22002 36898 22306 36902
rect 22342 37198 22966 37202
rect 22342 36902 22346 37198
rect 22346 36902 22962 37198
rect 22962 36902 22966 37198
rect 22342 36898 22966 36902
rect 23002 37198 23306 37202
rect 23002 36902 23006 37198
rect 23006 36902 23302 37198
rect 23302 36902 23306 37198
rect 23002 36898 23306 36902
rect 23342 37198 23966 37202
rect 23342 36902 23346 37198
rect 23346 36902 23962 37198
rect 23962 36902 23966 37198
rect 23342 36898 23966 36902
rect 24002 37198 24306 37202
rect 24002 36902 24006 37198
rect 24006 36902 24302 37198
rect 24302 36902 24306 37198
rect 24002 36898 24306 36902
rect 24342 37198 24966 37202
rect 24342 36902 24346 37198
rect 24346 36902 24962 37198
rect 24962 36902 24966 37198
rect 24342 36898 24966 36902
rect 25002 37198 25306 37202
rect 25002 36902 25006 37198
rect 25006 36902 25302 37198
rect 25302 36902 25306 37198
rect 25002 36898 25306 36902
rect 25342 37198 25966 37202
rect 25342 36902 25346 37198
rect 25346 36902 25962 37198
rect 25962 36902 25966 37198
rect 25342 36898 25966 36902
rect 26002 37198 26306 37202
rect 26002 36902 26006 37198
rect 26006 36902 26302 37198
rect 26302 36902 26306 37198
rect 26002 36898 26306 36902
rect 26342 37198 26966 37202
rect 26342 36902 26346 37198
rect 26346 36902 26962 37198
rect 26962 36902 26966 37198
rect 26342 36898 26966 36902
rect 27002 37198 27306 37202
rect 27002 36902 27006 37198
rect 27006 36902 27302 37198
rect 27302 36902 27306 37198
rect 27002 36898 27306 36902
rect 27342 37198 27966 37202
rect 27342 36902 27346 37198
rect 27346 36902 27962 37198
rect 27962 36902 27966 37198
rect 27342 36898 27966 36902
rect 28002 37198 28306 37202
rect 28002 36902 28006 37198
rect 28006 36902 28302 37198
rect 28302 36902 28306 37198
rect 28002 36898 28306 36902
rect 28342 37198 28966 37202
rect 28342 36902 28346 37198
rect 28346 36902 28962 37198
rect 28962 36902 28966 37198
rect 28342 36898 28966 36902
rect 29002 37198 29306 37202
rect 29002 36902 29006 37198
rect 29006 36902 29302 37198
rect 29302 36902 29306 37198
rect 29002 36898 29306 36902
rect 29342 37198 29966 37202
rect 29342 36902 29346 37198
rect 29346 36902 29962 37198
rect 29962 36902 29966 37198
rect 29342 36898 29966 36902
rect 30002 37198 30306 37202
rect 30002 36902 30006 37198
rect 30006 36902 30302 37198
rect 30302 36902 30306 37198
rect 30002 36898 30306 36902
rect 30342 37198 30966 37202
rect 30342 36902 30346 37198
rect 30346 36902 30962 37198
rect 30962 36902 30966 37198
rect 30342 36898 30966 36902
rect 31002 37198 31306 37202
rect 31002 36902 31006 37198
rect 31006 36902 31302 37198
rect 31302 36902 31306 37198
rect 31002 36898 31306 36902
rect 31342 37198 31966 37202
rect 31342 36902 31346 37198
rect 31346 36902 31962 37198
rect 31962 36902 31966 37198
rect 31342 36898 31966 36902
rect 32002 37198 32306 37202
rect 32002 36902 32006 37198
rect 32006 36902 32302 37198
rect 32302 36902 32306 37198
rect 32002 36898 32306 36902
rect 32342 37198 32966 37202
rect 32342 36902 32346 37198
rect 32346 36902 32962 37198
rect 32962 36902 32966 37198
rect 32342 36898 32966 36902
rect 33002 37198 33306 37202
rect 33002 36902 33006 37198
rect 33006 36902 33302 37198
rect 33302 36902 33306 37198
rect 33002 36898 33306 36902
rect 33342 37198 33966 37202
rect 33342 36902 33346 37198
rect 33346 36902 33962 37198
rect 33962 36902 33966 37198
rect 33342 36898 33966 36902
rect 34002 37198 34306 37202
rect 34002 36902 34006 37198
rect 34006 36902 34302 37198
rect 34302 36902 34306 37198
rect 34002 36898 34306 36902
rect 34342 37198 34646 37202
rect 34342 36902 34346 37198
rect 34346 36902 34642 37198
rect 34642 36902 34646 37198
rect 34342 36898 34646 36902
rect 10002 36858 10306 36862
rect 10002 36242 10006 36858
rect 10006 36242 10302 36858
rect 10302 36242 10306 36858
rect 10002 36238 10306 36242
rect 11002 36858 11306 36862
rect 11002 36242 11006 36858
rect 11006 36242 11302 36858
rect 11302 36242 11306 36858
rect 11002 36238 11306 36242
rect 12002 36858 12306 36862
rect 12002 36242 12006 36858
rect 12006 36242 12302 36858
rect 12302 36242 12306 36858
rect 12002 36238 12306 36242
rect 13002 36858 13306 36862
rect 13002 36242 13006 36858
rect 13006 36242 13302 36858
rect 13302 36242 13306 36858
rect 13002 36238 13306 36242
rect 14002 36858 14306 36862
rect 14002 36242 14006 36858
rect 14006 36242 14302 36858
rect 14302 36242 14306 36858
rect 14002 36238 14306 36242
rect 15002 36858 15306 36862
rect 15002 36242 15006 36858
rect 15006 36242 15302 36858
rect 15302 36242 15306 36858
rect 15002 36238 15306 36242
rect 16002 36858 16306 36862
rect 16002 36242 16006 36858
rect 16006 36242 16302 36858
rect 16302 36242 16306 36858
rect 16002 36238 16306 36242
rect 17002 36858 17306 36862
rect 17002 36242 17006 36858
rect 17006 36242 17302 36858
rect 17302 36242 17306 36858
rect 17002 36238 17306 36242
rect 18002 36858 18306 36862
rect 18002 36242 18006 36858
rect 18006 36242 18302 36858
rect 18302 36242 18306 36858
rect 18002 36238 18306 36242
rect 19002 36858 19306 36862
rect 19002 36242 19006 36858
rect 19006 36242 19302 36858
rect 19302 36242 19306 36858
rect 19002 36238 19306 36242
rect 20002 36858 20306 36862
rect 20002 36242 20006 36858
rect 20006 36242 20302 36858
rect 20302 36242 20306 36858
rect 20002 36238 20306 36242
rect 21002 36858 21306 36862
rect 21002 36242 21006 36858
rect 21006 36242 21302 36858
rect 21302 36242 21306 36858
rect 21002 36238 21306 36242
rect 22002 36858 22306 36862
rect 22002 36242 22006 36858
rect 22006 36242 22302 36858
rect 22302 36242 22306 36858
rect 22002 36238 22306 36242
rect 23002 36858 23306 36862
rect 23002 36242 23006 36858
rect 23006 36242 23302 36858
rect 23302 36242 23306 36858
rect 23002 36238 23306 36242
rect 24002 36858 24306 36862
rect 24002 36242 24006 36858
rect 24006 36242 24302 36858
rect 24302 36242 24306 36858
rect 24002 36238 24306 36242
rect 25002 36858 25306 36862
rect 25002 36242 25006 36858
rect 25006 36242 25302 36858
rect 25302 36242 25306 36858
rect 25002 36238 25306 36242
rect 26002 36858 26306 36862
rect 26002 36242 26006 36858
rect 26006 36242 26302 36858
rect 26302 36242 26306 36858
rect 26002 36238 26306 36242
rect 27002 36858 27306 36862
rect 27002 36242 27006 36858
rect 27006 36242 27302 36858
rect 27302 36242 27306 36858
rect 27002 36238 27306 36242
rect 28002 36858 28306 36862
rect 28002 36242 28006 36858
rect 28006 36242 28302 36858
rect 28302 36242 28306 36858
rect 28002 36238 28306 36242
rect 29002 36858 29306 36862
rect 29002 36242 29006 36858
rect 29006 36242 29302 36858
rect 29302 36242 29306 36858
rect 29002 36238 29306 36242
rect 30002 36858 30306 36862
rect 30002 36242 30006 36858
rect 30006 36242 30302 36858
rect 30302 36242 30306 36858
rect 30002 36238 30306 36242
rect 31002 36858 31306 36862
rect 31002 36242 31006 36858
rect 31006 36242 31302 36858
rect 31302 36242 31306 36858
rect 31002 36238 31306 36242
rect 32002 36858 32306 36862
rect 32002 36242 32006 36858
rect 32006 36242 32302 36858
rect 32302 36242 32306 36858
rect 32002 36238 32306 36242
rect 33002 36858 33306 36862
rect 33002 36242 33006 36858
rect 33006 36242 33302 36858
rect 33302 36242 33306 36858
rect 33002 36238 33306 36242
rect 34002 36858 34306 36862
rect 34002 36242 34006 36858
rect 34006 36242 34302 36858
rect 34302 36242 34306 36858
rect 34002 36238 34306 36242
rect 9662 36198 9966 36202
rect 9662 35902 9666 36198
rect 9666 35902 9962 36198
rect 9962 35902 9966 36198
rect 9662 35898 9966 35902
rect 10002 36198 10306 36202
rect 10002 35902 10006 36198
rect 10006 35902 10302 36198
rect 10302 35902 10306 36198
rect 10002 35898 10306 35902
rect 10342 36198 10966 36202
rect 10342 35902 10346 36198
rect 10346 35902 10962 36198
rect 10962 35902 10966 36198
rect 10342 35898 10966 35902
rect 11002 36198 11306 36202
rect 11002 35902 11006 36198
rect 11006 35902 11302 36198
rect 11302 35902 11306 36198
rect 11002 35898 11306 35902
rect 11342 36198 11966 36202
rect 11342 35902 11346 36198
rect 11346 35902 11962 36198
rect 11962 35902 11966 36198
rect 11342 35898 11966 35902
rect 12002 36198 12306 36202
rect 12002 35902 12006 36198
rect 12006 35902 12302 36198
rect 12302 35902 12306 36198
rect 12002 35898 12306 35902
rect 12342 36198 12966 36202
rect 12342 35902 12346 36198
rect 12346 35902 12962 36198
rect 12962 35902 12966 36198
rect 12342 35898 12966 35902
rect 13002 36198 13306 36202
rect 13002 35902 13006 36198
rect 13006 35902 13302 36198
rect 13302 35902 13306 36198
rect 13002 35898 13306 35902
rect 13342 36198 13966 36202
rect 13342 35902 13346 36198
rect 13346 35902 13962 36198
rect 13962 35902 13966 36198
rect 13342 35898 13966 35902
rect 14002 36198 14306 36202
rect 14002 35902 14006 36198
rect 14006 35902 14302 36198
rect 14302 35902 14306 36198
rect 14002 35898 14306 35902
rect 14342 36198 14966 36202
rect 14342 35902 14346 36198
rect 14346 35902 14962 36198
rect 14962 35902 14966 36198
rect 14342 35898 14966 35902
rect 15002 36198 15306 36202
rect 15002 35902 15006 36198
rect 15006 35902 15302 36198
rect 15302 35902 15306 36198
rect 15002 35898 15306 35902
rect 15342 36198 15966 36202
rect 15342 35902 15346 36198
rect 15346 35902 15962 36198
rect 15962 35902 15966 36198
rect 15342 35898 15966 35902
rect 16002 36198 16306 36202
rect 16002 35902 16006 36198
rect 16006 35902 16302 36198
rect 16302 35902 16306 36198
rect 16002 35898 16306 35902
rect 16342 36198 16966 36202
rect 16342 35902 16346 36198
rect 16346 35902 16962 36198
rect 16962 35902 16966 36198
rect 16342 35898 16966 35902
rect 17002 36198 17306 36202
rect 17002 35902 17006 36198
rect 17006 35902 17302 36198
rect 17302 35902 17306 36198
rect 17002 35898 17306 35902
rect 17342 36198 17966 36202
rect 17342 35902 17346 36198
rect 17346 35902 17962 36198
rect 17962 35902 17966 36198
rect 17342 35898 17966 35902
rect 18002 36198 18306 36202
rect 18002 35902 18006 36198
rect 18006 35902 18302 36198
rect 18302 35902 18306 36198
rect 18002 35898 18306 35902
rect 18342 36198 18966 36202
rect 18342 35902 18346 36198
rect 18346 35902 18962 36198
rect 18962 35902 18966 36198
rect 18342 35898 18966 35902
rect 19002 36198 19306 36202
rect 19002 35902 19006 36198
rect 19006 35902 19302 36198
rect 19302 35902 19306 36198
rect 19002 35898 19306 35902
rect 19342 36198 19966 36202
rect 19342 35902 19346 36198
rect 19346 35902 19962 36198
rect 19962 35902 19966 36198
rect 19342 35898 19966 35902
rect 20002 36198 20306 36202
rect 20002 35902 20006 36198
rect 20006 35902 20302 36198
rect 20302 35902 20306 36198
rect 20002 35898 20306 35902
rect 20342 36198 20966 36202
rect 20342 35902 20346 36198
rect 20346 35902 20962 36198
rect 20962 35902 20966 36198
rect 20342 35898 20966 35902
rect 21002 36198 21306 36202
rect 21002 35902 21006 36198
rect 21006 35902 21302 36198
rect 21302 35902 21306 36198
rect 21002 35898 21306 35902
rect 21342 36198 21966 36202
rect 21342 35902 21346 36198
rect 21346 35902 21962 36198
rect 21962 35902 21966 36198
rect 21342 35898 21966 35902
rect 22002 36198 22306 36202
rect 22002 35902 22006 36198
rect 22006 35902 22302 36198
rect 22302 35902 22306 36198
rect 22002 35898 22306 35902
rect 22342 36198 22966 36202
rect 22342 35902 22346 36198
rect 22346 35902 22962 36198
rect 22962 35902 22966 36198
rect 22342 35898 22966 35902
rect 23002 36198 23306 36202
rect 23002 35902 23006 36198
rect 23006 35902 23302 36198
rect 23302 35902 23306 36198
rect 23002 35898 23306 35902
rect 23342 36198 23966 36202
rect 23342 35902 23346 36198
rect 23346 35902 23962 36198
rect 23962 35902 23966 36198
rect 23342 35898 23966 35902
rect 24002 36198 24306 36202
rect 24002 35902 24006 36198
rect 24006 35902 24302 36198
rect 24302 35902 24306 36198
rect 24002 35898 24306 35902
rect 24342 36198 24966 36202
rect 24342 35902 24346 36198
rect 24346 35902 24962 36198
rect 24962 35902 24966 36198
rect 24342 35898 24966 35902
rect 25002 36198 25306 36202
rect 25002 35902 25006 36198
rect 25006 35902 25302 36198
rect 25302 35902 25306 36198
rect 25002 35898 25306 35902
rect 25342 36198 25966 36202
rect 25342 35902 25346 36198
rect 25346 35902 25962 36198
rect 25962 35902 25966 36198
rect 25342 35898 25966 35902
rect 26002 36198 26306 36202
rect 26002 35902 26006 36198
rect 26006 35902 26302 36198
rect 26302 35902 26306 36198
rect 26002 35898 26306 35902
rect 26342 36198 26966 36202
rect 26342 35902 26346 36198
rect 26346 35902 26962 36198
rect 26962 35902 26966 36198
rect 26342 35898 26966 35902
rect 27002 36198 27306 36202
rect 27002 35902 27006 36198
rect 27006 35902 27302 36198
rect 27302 35902 27306 36198
rect 27002 35898 27306 35902
rect 27342 36198 27966 36202
rect 27342 35902 27346 36198
rect 27346 35902 27962 36198
rect 27962 35902 27966 36198
rect 27342 35898 27966 35902
rect 28002 36198 28306 36202
rect 28002 35902 28006 36198
rect 28006 35902 28302 36198
rect 28302 35902 28306 36198
rect 28002 35898 28306 35902
rect 28342 36198 28966 36202
rect 28342 35902 28346 36198
rect 28346 35902 28962 36198
rect 28962 35902 28966 36198
rect 28342 35898 28966 35902
rect 29002 36198 29306 36202
rect 29002 35902 29006 36198
rect 29006 35902 29302 36198
rect 29302 35902 29306 36198
rect 29002 35898 29306 35902
rect 29342 36198 29966 36202
rect 29342 35902 29346 36198
rect 29346 35902 29962 36198
rect 29962 35902 29966 36198
rect 29342 35898 29966 35902
rect 30002 36198 30306 36202
rect 30002 35902 30006 36198
rect 30006 35902 30302 36198
rect 30302 35902 30306 36198
rect 30002 35898 30306 35902
rect 30342 36198 30966 36202
rect 30342 35902 30346 36198
rect 30346 35902 30962 36198
rect 30962 35902 30966 36198
rect 30342 35898 30966 35902
rect 31002 36198 31306 36202
rect 31002 35902 31006 36198
rect 31006 35902 31302 36198
rect 31302 35902 31306 36198
rect 31002 35898 31306 35902
rect 31342 36198 31966 36202
rect 31342 35902 31346 36198
rect 31346 35902 31962 36198
rect 31962 35902 31966 36198
rect 31342 35898 31966 35902
rect 32002 36198 32306 36202
rect 32002 35902 32006 36198
rect 32006 35902 32302 36198
rect 32302 35902 32306 36198
rect 32002 35898 32306 35902
rect 32342 36198 32966 36202
rect 32342 35902 32346 36198
rect 32346 35902 32962 36198
rect 32962 35902 32966 36198
rect 32342 35898 32966 35902
rect 33002 36198 33306 36202
rect 33002 35902 33006 36198
rect 33006 35902 33302 36198
rect 33302 35902 33306 36198
rect 33002 35898 33306 35902
rect 33342 36198 33966 36202
rect 33342 35902 33346 36198
rect 33346 35902 33962 36198
rect 33962 35902 33966 36198
rect 33342 35898 33966 35902
rect 34002 36198 34306 36202
rect 34002 35902 34006 36198
rect 34006 35902 34302 36198
rect 34302 35902 34306 36198
rect 34002 35898 34306 35902
rect 34342 36198 34646 36202
rect 34342 35902 34346 36198
rect 34346 35902 34642 36198
rect 34642 35902 34646 36198
rect 34342 35898 34646 35902
rect 10002 35858 10306 35862
rect 10002 35242 10006 35858
rect 10006 35242 10302 35858
rect 10302 35242 10306 35858
rect 10002 35238 10306 35242
rect 11002 35858 11306 35862
rect 11002 35242 11006 35858
rect 11006 35242 11302 35858
rect 11302 35242 11306 35858
rect 11002 35238 11306 35242
rect 12002 35858 12306 35862
rect 12002 35242 12006 35858
rect 12006 35242 12302 35858
rect 12302 35242 12306 35858
rect 12002 35238 12306 35242
rect 13002 35858 13306 35862
rect 13002 35242 13006 35858
rect 13006 35242 13302 35858
rect 13302 35242 13306 35858
rect 13002 35238 13306 35242
rect 14002 35858 14306 35862
rect 14002 35242 14006 35858
rect 14006 35242 14302 35858
rect 14302 35242 14306 35858
rect 14002 35238 14306 35242
rect 15002 35858 15306 35862
rect 15002 35242 15006 35858
rect 15006 35242 15302 35858
rect 15302 35242 15306 35858
rect 15002 35238 15306 35242
rect 16002 35858 16306 35862
rect 16002 35242 16006 35858
rect 16006 35242 16302 35858
rect 16302 35242 16306 35858
rect 16002 35238 16306 35242
rect 17002 35858 17306 35862
rect 17002 35242 17006 35858
rect 17006 35242 17302 35858
rect 17302 35242 17306 35858
rect 17002 35238 17306 35242
rect 18002 35858 18306 35862
rect 18002 35242 18006 35858
rect 18006 35242 18302 35858
rect 18302 35242 18306 35858
rect 18002 35238 18306 35242
rect 19002 35858 19306 35862
rect 19002 35242 19006 35858
rect 19006 35242 19302 35858
rect 19302 35242 19306 35858
rect 19002 35238 19306 35242
rect 20002 35858 20306 35862
rect 20002 35242 20006 35858
rect 20006 35242 20302 35858
rect 20302 35242 20306 35858
rect 20002 35238 20306 35242
rect 21002 35858 21306 35862
rect 21002 35242 21006 35858
rect 21006 35242 21302 35858
rect 21302 35242 21306 35858
rect 21002 35238 21306 35242
rect 22002 35858 22306 35862
rect 22002 35242 22006 35858
rect 22006 35242 22302 35858
rect 22302 35242 22306 35858
rect 22002 35238 22306 35242
rect 23002 35858 23306 35862
rect 23002 35242 23006 35858
rect 23006 35242 23302 35858
rect 23302 35242 23306 35858
rect 23002 35238 23306 35242
rect 24002 35858 24306 35862
rect 24002 35242 24006 35858
rect 24006 35242 24302 35858
rect 24302 35242 24306 35858
rect 24002 35238 24306 35242
rect 25002 35858 25306 35862
rect 25002 35242 25006 35858
rect 25006 35242 25302 35858
rect 25302 35242 25306 35858
rect 25002 35238 25306 35242
rect 26002 35858 26306 35862
rect 26002 35242 26006 35858
rect 26006 35242 26302 35858
rect 26302 35242 26306 35858
rect 26002 35238 26306 35242
rect 27002 35858 27306 35862
rect 27002 35242 27006 35858
rect 27006 35242 27302 35858
rect 27302 35242 27306 35858
rect 27002 35238 27306 35242
rect 28002 35858 28306 35862
rect 28002 35242 28006 35858
rect 28006 35242 28302 35858
rect 28302 35242 28306 35858
rect 28002 35238 28306 35242
rect 29002 35858 29306 35862
rect 29002 35242 29006 35858
rect 29006 35242 29302 35858
rect 29302 35242 29306 35858
rect 29002 35238 29306 35242
rect 30002 35858 30306 35862
rect 30002 35242 30006 35858
rect 30006 35242 30302 35858
rect 30302 35242 30306 35858
rect 30002 35238 30306 35242
rect 31002 35858 31306 35862
rect 31002 35242 31006 35858
rect 31006 35242 31302 35858
rect 31302 35242 31306 35858
rect 31002 35238 31306 35242
rect 32002 35858 32306 35862
rect 32002 35242 32006 35858
rect 32006 35242 32302 35858
rect 32302 35242 32306 35858
rect 32002 35238 32306 35242
rect 33002 35858 33306 35862
rect 33002 35242 33006 35858
rect 33006 35242 33302 35858
rect 33302 35242 33306 35858
rect 33002 35238 33306 35242
rect 34002 35858 34306 35862
rect 34002 35242 34006 35858
rect 34006 35242 34302 35858
rect 34302 35242 34306 35858
rect 34002 35238 34306 35242
rect 9662 35198 9966 35202
rect 9662 34902 9666 35198
rect 9666 34902 9962 35198
rect 9962 34902 9966 35198
rect 9662 34898 9966 34902
rect 10002 35198 10306 35202
rect 10002 34902 10006 35198
rect 10006 34902 10302 35198
rect 10302 34902 10306 35198
rect 10002 34898 10306 34902
rect 10342 35198 10966 35202
rect 10342 34902 10346 35198
rect 10346 34902 10962 35198
rect 10962 34902 10966 35198
rect 10342 34898 10966 34902
rect 11002 35198 11306 35202
rect 11002 34902 11006 35198
rect 11006 34902 11302 35198
rect 11302 34902 11306 35198
rect 11002 34898 11306 34902
rect 11342 35198 11966 35202
rect 11342 34902 11346 35198
rect 11346 34902 11962 35198
rect 11962 34902 11966 35198
rect 11342 34898 11966 34902
rect 12002 35198 12306 35202
rect 12002 34902 12006 35198
rect 12006 34902 12302 35198
rect 12302 34902 12306 35198
rect 12002 34898 12306 34902
rect 12342 35198 12966 35202
rect 12342 34902 12346 35198
rect 12346 34902 12962 35198
rect 12962 34902 12966 35198
rect 12342 34898 12966 34902
rect 13002 35198 13306 35202
rect 13002 34902 13006 35198
rect 13006 34902 13302 35198
rect 13302 34902 13306 35198
rect 13002 34898 13306 34902
rect 13342 35198 13966 35202
rect 13342 34902 13346 35198
rect 13346 34902 13962 35198
rect 13962 34902 13966 35198
rect 13342 34898 13966 34902
rect 14002 35198 14306 35202
rect 14002 34902 14006 35198
rect 14006 34902 14302 35198
rect 14302 34902 14306 35198
rect 14002 34898 14306 34902
rect 14342 35198 14966 35202
rect 14342 34902 14346 35198
rect 14346 34902 14962 35198
rect 14962 34902 14966 35198
rect 14342 34898 14966 34902
rect 15002 35198 15306 35202
rect 15002 34902 15006 35198
rect 15006 34902 15302 35198
rect 15302 34902 15306 35198
rect 15002 34898 15306 34902
rect 15342 35198 15966 35202
rect 15342 34902 15346 35198
rect 15346 34902 15962 35198
rect 15962 34902 15966 35198
rect 15342 34898 15966 34902
rect 16002 35198 16306 35202
rect 16002 34902 16006 35198
rect 16006 34902 16302 35198
rect 16302 34902 16306 35198
rect 16002 34898 16306 34902
rect 16342 35198 16966 35202
rect 16342 34902 16346 35198
rect 16346 34902 16962 35198
rect 16962 34902 16966 35198
rect 16342 34898 16966 34902
rect 17002 35198 17306 35202
rect 17002 34902 17006 35198
rect 17006 34902 17302 35198
rect 17302 34902 17306 35198
rect 17002 34898 17306 34902
rect 17342 35198 17966 35202
rect 17342 34902 17346 35198
rect 17346 34902 17962 35198
rect 17962 34902 17966 35198
rect 17342 34898 17966 34902
rect 18002 35198 18306 35202
rect 18002 34902 18006 35198
rect 18006 34902 18302 35198
rect 18302 34902 18306 35198
rect 18002 34898 18306 34902
rect 18342 35198 18966 35202
rect 18342 34902 18346 35198
rect 18346 34902 18962 35198
rect 18962 34902 18966 35198
rect 18342 34898 18966 34902
rect 19002 35198 19306 35202
rect 19002 34902 19006 35198
rect 19006 34902 19302 35198
rect 19302 34902 19306 35198
rect 19002 34898 19306 34902
rect 19342 35198 19966 35202
rect 19342 34902 19346 35198
rect 19346 34902 19962 35198
rect 19962 34902 19966 35198
rect 19342 34898 19966 34902
rect 20002 35198 20306 35202
rect 20002 34902 20006 35198
rect 20006 34902 20302 35198
rect 20302 34902 20306 35198
rect 20002 34898 20306 34902
rect 20342 35198 20966 35202
rect 20342 34902 20346 35198
rect 20346 34902 20962 35198
rect 20962 34902 20966 35198
rect 20342 34898 20966 34902
rect 21002 35198 21306 35202
rect 21002 34902 21006 35198
rect 21006 34902 21302 35198
rect 21302 34902 21306 35198
rect 21002 34898 21306 34902
rect 21342 35198 21966 35202
rect 21342 34902 21346 35198
rect 21346 34902 21962 35198
rect 21962 34902 21966 35198
rect 21342 34898 21966 34902
rect 22002 35198 22306 35202
rect 22002 34902 22006 35198
rect 22006 34902 22302 35198
rect 22302 34902 22306 35198
rect 22002 34898 22306 34902
rect 22342 35198 22966 35202
rect 22342 34902 22346 35198
rect 22346 34902 22962 35198
rect 22962 34902 22966 35198
rect 22342 34898 22966 34902
rect 23002 35198 23306 35202
rect 23002 34902 23006 35198
rect 23006 34902 23302 35198
rect 23302 34902 23306 35198
rect 23002 34898 23306 34902
rect 23342 35198 23966 35202
rect 23342 34902 23346 35198
rect 23346 34902 23962 35198
rect 23962 34902 23966 35198
rect 23342 34898 23966 34902
rect 24002 35198 24306 35202
rect 24002 34902 24006 35198
rect 24006 34902 24302 35198
rect 24302 34902 24306 35198
rect 24002 34898 24306 34902
rect 24342 35198 24966 35202
rect 24342 34902 24346 35198
rect 24346 34902 24962 35198
rect 24962 34902 24966 35198
rect 24342 34898 24966 34902
rect 25002 35198 25306 35202
rect 25002 34902 25006 35198
rect 25006 34902 25302 35198
rect 25302 34902 25306 35198
rect 25002 34898 25306 34902
rect 25342 35198 25966 35202
rect 25342 34902 25346 35198
rect 25346 34902 25962 35198
rect 25962 34902 25966 35198
rect 25342 34898 25966 34902
rect 26002 35198 26306 35202
rect 26002 34902 26006 35198
rect 26006 34902 26302 35198
rect 26302 34902 26306 35198
rect 26002 34898 26306 34902
rect 26342 35198 26966 35202
rect 26342 34902 26346 35198
rect 26346 34902 26962 35198
rect 26962 34902 26966 35198
rect 26342 34898 26966 34902
rect 27002 35198 27306 35202
rect 27002 34902 27006 35198
rect 27006 34902 27302 35198
rect 27302 34902 27306 35198
rect 27002 34898 27306 34902
rect 27342 35198 27966 35202
rect 27342 34902 27346 35198
rect 27346 34902 27962 35198
rect 27962 34902 27966 35198
rect 27342 34898 27966 34902
rect 28002 35198 28306 35202
rect 28002 34902 28006 35198
rect 28006 34902 28302 35198
rect 28302 34902 28306 35198
rect 28002 34898 28306 34902
rect 28342 35198 28966 35202
rect 28342 34902 28346 35198
rect 28346 34902 28962 35198
rect 28962 34902 28966 35198
rect 28342 34898 28966 34902
rect 29002 35198 29306 35202
rect 29002 34902 29006 35198
rect 29006 34902 29302 35198
rect 29302 34902 29306 35198
rect 29002 34898 29306 34902
rect 29342 35198 29966 35202
rect 29342 34902 29346 35198
rect 29346 34902 29962 35198
rect 29962 34902 29966 35198
rect 29342 34898 29966 34902
rect 30002 35198 30306 35202
rect 30002 34902 30006 35198
rect 30006 34902 30302 35198
rect 30302 34902 30306 35198
rect 30002 34898 30306 34902
rect 30342 35198 30966 35202
rect 30342 34902 30346 35198
rect 30346 34902 30962 35198
rect 30962 34902 30966 35198
rect 30342 34898 30966 34902
rect 31002 35198 31306 35202
rect 31002 34902 31006 35198
rect 31006 34902 31302 35198
rect 31302 34902 31306 35198
rect 31002 34898 31306 34902
rect 31342 35198 31966 35202
rect 31342 34902 31346 35198
rect 31346 34902 31962 35198
rect 31962 34902 31966 35198
rect 31342 34898 31966 34902
rect 32002 35198 32306 35202
rect 32002 34902 32006 35198
rect 32006 34902 32302 35198
rect 32302 34902 32306 35198
rect 32002 34898 32306 34902
rect 32342 35198 32966 35202
rect 32342 34902 32346 35198
rect 32346 34902 32962 35198
rect 32962 34902 32966 35198
rect 32342 34898 32966 34902
rect 33002 35198 33306 35202
rect 33002 34902 33006 35198
rect 33006 34902 33302 35198
rect 33302 34902 33306 35198
rect 33002 34898 33306 34902
rect 33342 35198 33966 35202
rect 33342 34902 33346 35198
rect 33346 34902 33962 35198
rect 33962 34902 33966 35198
rect 33342 34898 33966 34902
rect 34002 35198 34306 35202
rect 34002 34902 34006 35198
rect 34006 34902 34302 35198
rect 34302 34902 34306 35198
rect 34002 34898 34306 34902
rect 34342 35198 34646 35202
rect 34342 34902 34346 35198
rect 34346 34902 34642 35198
rect 34642 34902 34646 35198
rect 34342 34898 34646 34902
rect 10002 34858 10306 34862
rect 10002 34242 10006 34858
rect 10006 34242 10302 34858
rect 10302 34242 10306 34858
rect 10002 34238 10306 34242
rect 11002 34858 11306 34862
rect 11002 34242 11006 34858
rect 11006 34242 11302 34858
rect 11302 34242 11306 34858
rect 11002 34238 11306 34242
rect 12002 34858 12306 34862
rect 12002 34242 12006 34858
rect 12006 34242 12302 34858
rect 12302 34242 12306 34858
rect 12002 34238 12306 34242
rect 13002 34858 13306 34862
rect 13002 34242 13006 34858
rect 13006 34242 13302 34858
rect 13302 34242 13306 34858
rect 13002 34238 13306 34242
rect 14002 34858 14306 34862
rect 14002 34242 14006 34858
rect 14006 34242 14302 34858
rect 14302 34242 14306 34858
rect 14002 34238 14306 34242
rect 15002 34858 15306 34862
rect 15002 34242 15006 34858
rect 15006 34242 15302 34858
rect 15302 34242 15306 34858
rect 15002 34238 15306 34242
rect 16002 34858 16306 34862
rect 16002 34242 16006 34858
rect 16006 34242 16302 34858
rect 16302 34242 16306 34858
rect 16002 34238 16306 34242
rect 17002 34858 17306 34862
rect 17002 34242 17006 34858
rect 17006 34242 17302 34858
rect 17302 34242 17306 34858
rect 17002 34238 17306 34242
rect 18002 34858 18306 34862
rect 18002 34242 18006 34858
rect 18006 34242 18302 34858
rect 18302 34242 18306 34858
rect 18002 34238 18306 34242
rect 19002 34858 19306 34862
rect 19002 34242 19006 34858
rect 19006 34242 19302 34858
rect 19302 34242 19306 34858
rect 19002 34238 19306 34242
rect 20002 34858 20306 34862
rect 20002 34242 20006 34858
rect 20006 34242 20302 34858
rect 20302 34242 20306 34858
rect 20002 34238 20306 34242
rect 21002 34858 21306 34862
rect 21002 34242 21006 34858
rect 21006 34242 21302 34858
rect 21302 34242 21306 34858
rect 21002 34238 21306 34242
rect 22002 34858 22306 34862
rect 22002 34242 22006 34858
rect 22006 34242 22302 34858
rect 22302 34242 22306 34858
rect 22002 34238 22306 34242
rect 23002 34858 23306 34862
rect 23002 34242 23006 34858
rect 23006 34242 23302 34858
rect 23302 34242 23306 34858
rect 23002 34238 23306 34242
rect 24002 34858 24306 34862
rect 24002 34242 24006 34858
rect 24006 34242 24302 34858
rect 24302 34242 24306 34858
rect 24002 34238 24306 34242
rect 25002 34858 25306 34862
rect 25002 34242 25006 34858
rect 25006 34242 25302 34858
rect 25302 34242 25306 34858
rect 25002 34238 25306 34242
rect 26002 34858 26306 34862
rect 26002 34242 26006 34858
rect 26006 34242 26302 34858
rect 26302 34242 26306 34858
rect 26002 34238 26306 34242
rect 27002 34858 27306 34862
rect 27002 34242 27006 34858
rect 27006 34242 27302 34858
rect 27302 34242 27306 34858
rect 27002 34238 27306 34242
rect 28002 34858 28306 34862
rect 28002 34242 28006 34858
rect 28006 34242 28302 34858
rect 28302 34242 28306 34858
rect 28002 34238 28306 34242
rect 29002 34858 29306 34862
rect 29002 34242 29006 34858
rect 29006 34242 29302 34858
rect 29302 34242 29306 34858
rect 29002 34238 29306 34242
rect 30002 34858 30306 34862
rect 30002 34242 30006 34858
rect 30006 34242 30302 34858
rect 30302 34242 30306 34858
rect 30002 34238 30306 34242
rect 31002 34858 31306 34862
rect 31002 34242 31006 34858
rect 31006 34242 31302 34858
rect 31302 34242 31306 34858
rect 31002 34238 31306 34242
rect 32002 34858 32306 34862
rect 32002 34242 32006 34858
rect 32006 34242 32302 34858
rect 32302 34242 32306 34858
rect 32002 34238 32306 34242
rect 33002 34858 33306 34862
rect 33002 34242 33006 34858
rect 33006 34242 33302 34858
rect 33302 34242 33306 34858
rect 33002 34238 33306 34242
rect 34002 34858 34306 34862
rect 34002 34242 34006 34858
rect 34006 34242 34302 34858
rect 34302 34242 34306 34858
rect 34002 34238 34306 34242
rect 9662 34198 9966 34202
rect 9662 33902 9666 34198
rect 9666 33902 9962 34198
rect 9962 33902 9966 34198
rect 9662 33898 9966 33902
rect 10002 34198 10306 34202
rect 10002 33902 10006 34198
rect 10006 33902 10302 34198
rect 10302 33902 10306 34198
rect 10002 33898 10306 33902
rect 10342 34198 10966 34202
rect 10342 33902 10346 34198
rect 10346 33902 10962 34198
rect 10962 33902 10966 34198
rect 10342 33898 10966 33902
rect 11002 34198 11306 34202
rect 11002 33902 11006 34198
rect 11006 33902 11302 34198
rect 11302 33902 11306 34198
rect 11002 33898 11306 33902
rect 11342 34198 11966 34202
rect 11342 33902 11346 34198
rect 11346 33902 11962 34198
rect 11962 33902 11966 34198
rect 11342 33898 11966 33902
rect 12002 34198 12306 34202
rect 12002 33902 12006 34198
rect 12006 33902 12302 34198
rect 12302 33902 12306 34198
rect 12002 33898 12306 33902
rect 12342 34198 12966 34202
rect 12342 33902 12346 34198
rect 12346 33902 12962 34198
rect 12962 33902 12966 34198
rect 12342 33898 12966 33902
rect 13002 34198 13306 34202
rect 13002 33902 13006 34198
rect 13006 33902 13302 34198
rect 13302 33902 13306 34198
rect 13002 33898 13306 33902
rect 13342 34198 13966 34202
rect 13342 33902 13346 34198
rect 13346 33902 13962 34198
rect 13962 33902 13966 34198
rect 13342 33898 13966 33902
rect 14002 34198 14306 34202
rect 14002 33902 14006 34198
rect 14006 33902 14302 34198
rect 14302 33902 14306 34198
rect 14002 33898 14306 33902
rect 14342 34198 14966 34202
rect 14342 33902 14346 34198
rect 14346 33902 14962 34198
rect 14962 33902 14966 34198
rect 14342 33898 14966 33902
rect 15002 34198 15306 34202
rect 15002 33902 15006 34198
rect 15006 33902 15302 34198
rect 15302 33902 15306 34198
rect 15002 33898 15306 33902
rect 15342 34198 15966 34202
rect 15342 33902 15346 34198
rect 15346 33902 15962 34198
rect 15962 33902 15966 34198
rect 15342 33898 15966 33902
rect 16002 34198 16306 34202
rect 16002 33902 16006 34198
rect 16006 33902 16302 34198
rect 16302 33902 16306 34198
rect 16002 33898 16306 33902
rect 16342 34198 16966 34202
rect 16342 33902 16346 34198
rect 16346 33902 16962 34198
rect 16962 33902 16966 34198
rect 16342 33898 16966 33902
rect 17002 34198 17306 34202
rect 17002 33902 17006 34198
rect 17006 33902 17302 34198
rect 17302 33902 17306 34198
rect 17002 33898 17306 33902
rect 17342 34198 17966 34202
rect 17342 33902 17346 34198
rect 17346 33902 17962 34198
rect 17962 33902 17966 34198
rect 17342 33898 17966 33902
rect 18002 34198 18306 34202
rect 18002 33902 18006 34198
rect 18006 33902 18302 34198
rect 18302 33902 18306 34198
rect 18002 33898 18306 33902
rect 18342 34198 18966 34202
rect 18342 33902 18346 34198
rect 18346 33902 18962 34198
rect 18962 33902 18966 34198
rect 18342 33898 18966 33902
rect 19002 34198 19306 34202
rect 19002 33902 19006 34198
rect 19006 33902 19302 34198
rect 19302 33902 19306 34198
rect 19002 33898 19306 33902
rect 19342 34198 19966 34202
rect 19342 33902 19346 34198
rect 19346 33902 19962 34198
rect 19962 33902 19966 34198
rect 19342 33898 19966 33902
rect 20002 34198 20306 34202
rect 20002 33902 20006 34198
rect 20006 33902 20302 34198
rect 20302 33902 20306 34198
rect 20002 33898 20306 33902
rect 20342 34198 20966 34202
rect 20342 33902 20346 34198
rect 20346 33902 20962 34198
rect 20962 33902 20966 34198
rect 20342 33898 20966 33902
rect 21002 34198 21306 34202
rect 21002 33902 21006 34198
rect 21006 33902 21302 34198
rect 21302 33902 21306 34198
rect 21002 33898 21306 33902
rect 21342 34198 21966 34202
rect 21342 33902 21346 34198
rect 21346 33902 21962 34198
rect 21962 33902 21966 34198
rect 21342 33898 21966 33902
rect 22002 34198 22306 34202
rect 22002 33902 22006 34198
rect 22006 33902 22302 34198
rect 22302 33902 22306 34198
rect 22002 33898 22306 33902
rect 22342 34198 22966 34202
rect 22342 33902 22346 34198
rect 22346 33902 22962 34198
rect 22962 33902 22966 34198
rect 22342 33898 22966 33902
rect 23002 34198 23306 34202
rect 23002 33902 23006 34198
rect 23006 33902 23302 34198
rect 23302 33902 23306 34198
rect 23002 33898 23306 33902
rect 23342 34198 23966 34202
rect 23342 33902 23346 34198
rect 23346 33902 23962 34198
rect 23962 33902 23966 34198
rect 23342 33898 23966 33902
rect 24002 34198 24306 34202
rect 24002 33902 24006 34198
rect 24006 33902 24302 34198
rect 24302 33902 24306 34198
rect 24002 33898 24306 33902
rect 24342 34198 24966 34202
rect 24342 33902 24346 34198
rect 24346 33902 24962 34198
rect 24962 33902 24966 34198
rect 24342 33898 24966 33902
rect 25002 34198 25306 34202
rect 25002 33902 25006 34198
rect 25006 33902 25302 34198
rect 25302 33902 25306 34198
rect 25002 33898 25306 33902
rect 25342 34198 25966 34202
rect 25342 33902 25346 34198
rect 25346 33902 25962 34198
rect 25962 33902 25966 34198
rect 25342 33898 25966 33902
rect 26002 34198 26306 34202
rect 26002 33902 26006 34198
rect 26006 33902 26302 34198
rect 26302 33902 26306 34198
rect 26002 33898 26306 33902
rect 26342 34198 26966 34202
rect 26342 33902 26346 34198
rect 26346 33902 26962 34198
rect 26962 33902 26966 34198
rect 26342 33898 26966 33902
rect 27002 34198 27306 34202
rect 27002 33902 27006 34198
rect 27006 33902 27302 34198
rect 27302 33902 27306 34198
rect 27002 33898 27306 33902
rect 27342 34198 27966 34202
rect 27342 33902 27346 34198
rect 27346 33902 27962 34198
rect 27962 33902 27966 34198
rect 27342 33898 27966 33902
rect 28002 34198 28306 34202
rect 28002 33902 28006 34198
rect 28006 33902 28302 34198
rect 28302 33902 28306 34198
rect 28002 33898 28306 33902
rect 28342 34198 28966 34202
rect 28342 33902 28346 34198
rect 28346 33902 28962 34198
rect 28962 33902 28966 34198
rect 28342 33898 28966 33902
rect 29002 34198 29306 34202
rect 29002 33902 29006 34198
rect 29006 33902 29302 34198
rect 29302 33902 29306 34198
rect 29002 33898 29306 33902
rect 29342 34198 29966 34202
rect 29342 33902 29346 34198
rect 29346 33902 29962 34198
rect 29962 33902 29966 34198
rect 29342 33898 29966 33902
rect 30002 34198 30306 34202
rect 30002 33902 30006 34198
rect 30006 33902 30302 34198
rect 30302 33902 30306 34198
rect 30002 33898 30306 33902
rect 30342 34198 30966 34202
rect 30342 33902 30346 34198
rect 30346 33902 30962 34198
rect 30962 33902 30966 34198
rect 30342 33898 30966 33902
rect 31002 34198 31306 34202
rect 31002 33902 31006 34198
rect 31006 33902 31302 34198
rect 31302 33902 31306 34198
rect 31002 33898 31306 33902
rect 31342 34198 31966 34202
rect 31342 33902 31346 34198
rect 31346 33902 31962 34198
rect 31962 33902 31966 34198
rect 31342 33898 31966 33902
rect 32002 34198 32306 34202
rect 32002 33902 32006 34198
rect 32006 33902 32302 34198
rect 32302 33902 32306 34198
rect 32002 33898 32306 33902
rect 32342 34198 32966 34202
rect 32342 33902 32346 34198
rect 32346 33902 32962 34198
rect 32962 33902 32966 34198
rect 32342 33898 32966 33902
rect 33002 34198 33306 34202
rect 33002 33902 33006 34198
rect 33006 33902 33302 34198
rect 33302 33902 33306 34198
rect 33002 33898 33306 33902
rect 33342 34198 33966 34202
rect 33342 33902 33346 34198
rect 33346 33902 33962 34198
rect 33962 33902 33966 34198
rect 33342 33898 33966 33902
rect 34002 34198 34306 34202
rect 34002 33902 34006 34198
rect 34006 33902 34302 34198
rect 34302 33902 34306 34198
rect 34002 33898 34306 33902
rect 34342 34198 34646 34202
rect 34342 33902 34346 34198
rect 34346 33902 34642 34198
rect 34642 33902 34646 34198
rect 34342 33898 34646 33902
rect 10002 33858 10306 33862
rect 10002 33242 10006 33858
rect 10006 33242 10302 33858
rect 10302 33242 10306 33858
rect 10002 33238 10306 33242
rect 11002 33858 11306 33862
rect 11002 33242 11006 33858
rect 11006 33242 11302 33858
rect 11302 33242 11306 33858
rect 11002 33238 11306 33242
rect 12002 33858 12306 33862
rect 12002 33242 12006 33858
rect 12006 33242 12302 33858
rect 12302 33242 12306 33858
rect 12002 33238 12306 33242
rect 13002 33858 13306 33862
rect 13002 33242 13006 33858
rect 13006 33242 13302 33858
rect 13302 33242 13306 33858
rect 13002 33238 13306 33242
rect 14002 33858 14306 33862
rect 14002 33242 14006 33858
rect 14006 33242 14302 33858
rect 14302 33242 14306 33858
rect 14002 33238 14306 33242
rect 15002 33858 15306 33862
rect 15002 33242 15006 33858
rect 15006 33242 15302 33858
rect 15302 33242 15306 33858
rect 15002 33238 15306 33242
rect 16002 33858 16306 33862
rect 16002 33242 16006 33858
rect 16006 33242 16302 33858
rect 16302 33242 16306 33858
rect 16002 33238 16306 33242
rect 17002 33858 17306 33862
rect 17002 33242 17006 33858
rect 17006 33242 17302 33858
rect 17302 33242 17306 33858
rect 17002 33238 17306 33242
rect 18002 33858 18306 33862
rect 18002 33242 18006 33858
rect 18006 33242 18302 33858
rect 18302 33242 18306 33858
rect 18002 33238 18306 33242
rect 19002 33858 19306 33862
rect 19002 33242 19006 33858
rect 19006 33242 19302 33858
rect 19302 33242 19306 33858
rect 19002 33238 19306 33242
rect 20002 33858 20306 33862
rect 20002 33242 20006 33858
rect 20006 33242 20302 33858
rect 20302 33242 20306 33858
rect 20002 33238 20306 33242
rect 21002 33858 21306 33862
rect 21002 33242 21006 33858
rect 21006 33242 21302 33858
rect 21302 33242 21306 33858
rect 21002 33238 21306 33242
rect 22002 33858 22306 33862
rect 22002 33242 22006 33858
rect 22006 33242 22302 33858
rect 22302 33242 22306 33858
rect 22002 33238 22306 33242
rect 23002 33858 23306 33862
rect 23002 33242 23006 33858
rect 23006 33242 23302 33858
rect 23302 33242 23306 33858
rect 23002 33238 23306 33242
rect 24002 33858 24306 33862
rect 24002 33242 24006 33858
rect 24006 33242 24302 33858
rect 24302 33242 24306 33858
rect 24002 33238 24306 33242
rect 25002 33858 25306 33862
rect 25002 33242 25006 33858
rect 25006 33242 25302 33858
rect 25302 33242 25306 33858
rect 25002 33238 25306 33242
rect 26002 33858 26306 33862
rect 26002 33242 26006 33858
rect 26006 33242 26302 33858
rect 26302 33242 26306 33858
rect 26002 33238 26306 33242
rect 27002 33858 27306 33862
rect 27002 33242 27006 33858
rect 27006 33242 27302 33858
rect 27302 33242 27306 33858
rect 27002 33238 27306 33242
rect 28002 33858 28306 33862
rect 28002 33242 28006 33858
rect 28006 33242 28302 33858
rect 28302 33242 28306 33858
rect 28002 33238 28306 33242
rect 29002 33858 29306 33862
rect 29002 33242 29006 33858
rect 29006 33242 29302 33858
rect 29302 33242 29306 33858
rect 29002 33238 29306 33242
rect 30002 33858 30306 33862
rect 30002 33242 30006 33858
rect 30006 33242 30302 33858
rect 30302 33242 30306 33858
rect 30002 33238 30306 33242
rect 31002 33858 31306 33862
rect 31002 33242 31006 33858
rect 31006 33242 31302 33858
rect 31302 33242 31306 33858
rect 31002 33238 31306 33242
rect 32002 33858 32306 33862
rect 32002 33242 32006 33858
rect 32006 33242 32302 33858
rect 32302 33242 32306 33858
rect 32002 33238 32306 33242
rect 33002 33858 33306 33862
rect 33002 33242 33006 33858
rect 33006 33242 33302 33858
rect 33302 33242 33306 33858
rect 33002 33238 33306 33242
rect 34002 33858 34306 33862
rect 34002 33242 34006 33858
rect 34006 33242 34302 33858
rect 34302 33242 34306 33858
rect 34002 33238 34306 33242
rect -74477 32858 -74173 32862
rect -74477 32242 -74473 32858
rect -74473 32242 -74177 32858
rect -74177 32242 -74173 32858
rect -74477 32238 -74173 32242
rect -73477 32858 -73173 32862
rect -73477 32242 -73473 32858
rect -73473 32242 -73177 32858
rect -73177 32242 -73173 32858
rect -73477 32238 -73173 32242
rect -72477 32858 -72173 32862
rect -72477 32242 -72473 32858
rect -72473 32242 -72177 32858
rect -72177 32242 -72173 32858
rect -72477 32238 -72173 32242
rect -71477 32858 -71173 32862
rect -71477 32242 -71473 32858
rect -71473 32242 -71177 32858
rect -71177 32242 -71173 32858
rect -71477 32238 -71173 32242
rect -70477 32858 -70173 32862
rect -70477 32242 -70473 32858
rect -70473 32242 -70177 32858
rect -70177 32242 -70173 32858
rect -70477 32238 -70173 32242
rect -69477 32858 -69173 32862
rect -69477 32242 -69473 32858
rect -69473 32242 -69177 32858
rect -69177 32242 -69173 32858
rect -69477 32238 -69173 32242
rect -68477 32858 -68173 32862
rect -68477 32242 -68473 32858
rect -68473 32242 -68177 32858
rect -68177 32242 -68173 32858
rect -68477 32238 -68173 32242
rect -67477 32858 -67173 32862
rect -67477 32242 -67473 32858
rect -67473 32242 -67177 32858
rect -67177 32242 -67173 32858
rect -67477 32238 -67173 32242
rect -66477 32858 -66173 32862
rect -66477 32242 -66473 32858
rect -66473 32242 -66177 32858
rect -66177 32242 -66173 32858
rect -66477 32238 -66173 32242
rect -65477 32858 -65173 32862
rect -65477 32242 -65473 32858
rect -65473 32242 -65177 32858
rect -65177 32242 -65173 32858
rect -65477 32238 -65173 32242
rect -64477 32858 -64173 32862
rect -64477 32242 -64473 32858
rect -64473 32242 -64177 32858
rect -64177 32242 -64173 32858
rect -64477 32238 -64173 32242
rect -63477 32858 -63173 32862
rect -63477 32242 -63473 32858
rect -63473 32242 -63177 32858
rect -63177 32242 -63173 32858
rect -63477 32238 -63173 32242
rect -62477 32858 -62173 32862
rect -62477 32242 -62473 32858
rect -62473 32242 -62177 32858
rect -62177 32242 -62173 32858
rect -62477 32238 -62173 32242
rect -61477 32858 -61173 32862
rect -61477 32242 -61473 32858
rect -61473 32242 -61177 32858
rect -61177 32242 -61173 32858
rect -61477 32238 -61173 32242
rect -60477 32858 -60173 32862
rect -60477 32242 -60473 32858
rect -60473 32242 -60177 32858
rect -60177 32242 -60173 32858
rect -60477 32238 -60173 32242
rect -59477 32858 -59173 32862
rect -59477 32242 -59473 32858
rect -59473 32242 -59177 32858
rect -59177 32242 -59173 32858
rect -59477 32238 -59173 32242
rect 9662 33198 9966 33202
rect 9662 32902 9666 33198
rect 9666 32902 9962 33198
rect 9962 32902 9966 33198
rect 9662 32898 9966 32902
rect 10002 33198 10306 33202
rect 10002 32902 10006 33198
rect 10006 32902 10302 33198
rect 10302 32902 10306 33198
rect 10002 32898 10306 32902
rect 10342 33198 10966 33202
rect 10342 32902 10346 33198
rect 10346 32902 10962 33198
rect 10962 32902 10966 33198
rect 10342 32898 10966 32902
rect 11002 33198 11306 33202
rect 11002 32902 11006 33198
rect 11006 32902 11302 33198
rect 11302 32902 11306 33198
rect 11002 32898 11306 32902
rect 11342 33198 11966 33202
rect 11342 32902 11346 33198
rect 11346 32902 11962 33198
rect 11962 32902 11966 33198
rect 11342 32898 11966 32902
rect 12002 33198 12306 33202
rect 12002 32902 12006 33198
rect 12006 32902 12302 33198
rect 12302 32902 12306 33198
rect 12002 32898 12306 32902
rect 12342 33198 12966 33202
rect 12342 32902 12346 33198
rect 12346 32902 12962 33198
rect 12962 32902 12966 33198
rect 12342 32898 12966 32902
rect 13002 33198 13306 33202
rect 13002 32902 13006 33198
rect 13006 32902 13302 33198
rect 13302 32902 13306 33198
rect 13002 32898 13306 32902
rect 13342 33198 13966 33202
rect 13342 32902 13346 33198
rect 13346 32902 13962 33198
rect 13962 32902 13966 33198
rect 13342 32898 13966 32902
rect 14002 33198 14306 33202
rect 14002 32902 14006 33198
rect 14006 32902 14302 33198
rect 14302 32902 14306 33198
rect 14002 32898 14306 32902
rect 14342 33198 14966 33202
rect 14342 32902 14346 33198
rect 14346 32902 14962 33198
rect 14962 32902 14966 33198
rect 14342 32898 14966 32902
rect 15002 33198 15306 33202
rect 15002 32902 15006 33198
rect 15006 32902 15302 33198
rect 15302 32902 15306 33198
rect 15002 32898 15306 32902
rect 15342 33198 15966 33202
rect 15342 32902 15346 33198
rect 15346 32902 15962 33198
rect 15962 32902 15966 33198
rect 15342 32898 15966 32902
rect 16002 33198 16306 33202
rect 16002 32902 16006 33198
rect 16006 32902 16302 33198
rect 16302 32902 16306 33198
rect 16002 32898 16306 32902
rect 16342 33198 16966 33202
rect 16342 32902 16346 33198
rect 16346 32902 16962 33198
rect 16962 32902 16966 33198
rect 16342 32898 16966 32902
rect 17002 33198 17306 33202
rect 17002 32902 17006 33198
rect 17006 32902 17302 33198
rect 17302 32902 17306 33198
rect 17002 32898 17306 32902
rect 17342 33198 17966 33202
rect 17342 32902 17346 33198
rect 17346 32902 17962 33198
rect 17962 32902 17966 33198
rect 17342 32898 17966 32902
rect 18002 33198 18306 33202
rect 18002 32902 18006 33198
rect 18006 32902 18302 33198
rect 18302 32902 18306 33198
rect 18002 32898 18306 32902
rect 18342 33198 18966 33202
rect 18342 32902 18346 33198
rect 18346 32902 18962 33198
rect 18962 32902 18966 33198
rect 18342 32898 18966 32902
rect 19002 33198 19306 33202
rect 19002 32902 19006 33198
rect 19006 32902 19302 33198
rect 19302 32902 19306 33198
rect 19002 32898 19306 32902
rect 19342 33198 19966 33202
rect 19342 32902 19346 33198
rect 19346 32902 19962 33198
rect 19962 32902 19966 33198
rect 19342 32898 19966 32902
rect 20002 33198 20306 33202
rect 20002 32902 20006 33198
rect 20006 32902 20302 33198
rect 20302 32902 20306 33198
rect 20002 32898 20306 32902
rect 20342 33198 20966 33202
rect 20342 32902 20346 33198
rect 20346 32902 20962 33198
rect 20962 32902 20966 33198
rect 20342 32898 20966 32902
rect 21002 33198 21306 33202
rect 21002 32902 21006 33198
rect 21006 32902 21302 33198
rect 21302 32902 21306 33198
rect 21002 32898 21306 32902
rect 21342 33198 21966 33202
rect 21342 32902 21346 33198
rect 21346 32902 21962 33198
rect 21962 32902 21966 33198
rect 21342 32898 21966 32902
rect 22002 33198 22306 33202
rect 22002 32902 22006 33198
rect 22006 32902 22302 33198
rect 22302 32902 22306 33198
rect 22002 32898 22306 32902
rect 22342 33198 22966 33202
rect 22342 32902 22346 33198
rect 22346 32902 22962 33198
rect 22962 32902 22966 33198
rect 22342 32898 22966 32902
rect 23002 33198 23306 33202
rect 23002 32902 23006 33198
rect 23006 32902 23302 33198
rect 23302 32902 23306 33198
rect 23002 32898 23306 32902
rect 23342 33198 23966 33202
rect 23342 32902 23346 33198
rect 23346 32902 23962 33198
rect 23962 32902 23966 33198
rect 23342 32898 23966 32902
rect 24002 33198 24306 33202
rect 24002 32902 24006 33198
rect 24006 32902 24302 33198
rect 24302 32902 24306 33198
rect 24002 32898 24306 32902
rect 24342 33198 24966 33202
rect 24342 32902 24346 33198
rect 24346 32902 24962 33198
rect 24962 32902 24966 33198
rect 24342 32898 24966 32902
rect 25002 33198 25306 33202
rect 25002 32902 25006 33198
rect 25006 32902 25302 33198
rect 25302 32902 25306 33198
rect 25002 32898 25306 32902
rect 25342 33198 25966 33202
rect 25342 32902 25346 33198
rect 25346 32902 25962 33198
rect 25962 32902 25966 33198
rect 25342 32898 25966 32902
rect 26002 33198 26306 33202
rect 26002 32902 26006 33198
rect 26006 32902 26302 33198
rect 26302 32902 26306 33198
rect 26002 32898 26306 32902
rect 26342 33198 26966 33202
rect 26342 32902 26346 33198
rect 26346 32902 26962 33198
rect 26962 32902 26966 33198
rect 26342 32898 26966 32902
rect 27002 33198 27306 33202
rect 27002 32902 27006 33198
rect 27006 32902 27302 33198
rect 27302 32902 27306 33198
rect 27002 32898 27306 32902
rect 27342 33198 27966 33202
rect 27342 32902 27346 33198
rect 27346 32902 27962 33198
rect 27962 32902 27966 33198
rect 27342 32898 27966 32902
rect 28002 33198 28306 33202
rect 28002 32902 28006 33198
rect 28006 32902 28302 33198
rect 28302 32902 28306 33198
rect 28002 32898 28306 32902
rect 28342 33198 28966 33202
rect 28342 32902 28346 33198
rect 28346 32902 28962 33198
rect 28962 32902 28966 33198
rect 28342 32898 28966 32902
rect 29002 33198 29306 33202
rect 29002 32902 29006 33198
rect 29006 32902 29302 33198
rect 29302 32902 29306 33198
rect 29002 32898 29306 32902
rect 29342 33198 29966 33202
rect 29342 32902 29346 33198
rect 29346 32902 29962 33198
rect 29962 32902 29966 33198
rect 29342 32898 29966 32902
rect 30002 33198 30306 33202
rect 30002 32902 30006 33198
rect 30006 32902 30302 33198
rect 30302 32902 30306 33198
rect 30002 32898 30306 32902
rect 30342 33198 30966 33202
rect 30342 32902 30346 33198
rect 30346 32902 30962 33198
rect 30962 32902 30966 33198
rect 30342 32898 30966 32902
rect 31002 33198 31306 33202
rect 31002 32902 31006 33198
rect 31006 32902 31302 33198
rect 31302 32902 31306 33198
rect 31002 32898 31306 32902
rect 31342 33198 31966 33202
rect 31342 32902 31346 33198
rect 31346 32902 31962 33198
rect 31962 32902 31966 33198
rect 31342 32898 31966 32902
rect 32002 33198 32306 33202
rect 32002 32902 32006 33198
rect 32006 32902 32302 33198
rect 32302 32902 32306 33198
rect 32002 32898 32306 32902
rect 32342 33198 32966 33202
rect 32342 32902 32346 33198
rect 32346 32902 32962 33198
rect 32962 32902 32966 33198
rect 32342 32898 32966 32902
rect 33002 33198 33306 33202
rect 33002 32902 33006 33198
rect 33006 32902 33302 33198
rect 33302 32902 33306 33198
rect 33002 32898 33306 32902
rect 33342 33198 33966 33202
rect 33342 32902 33346 33198
rect 33346 32902 33962 33198
rect 33962 32902 33966 33198
rect 33342 32898 33966 32902
rect 34002 33198 34306 33202
rect 34002 32902 34006 33198
rect 34006 32902 34302 33198
rect 34302 32902 34306 33198
rect 34002 32898 34306 32902
rect 34342 33198 34646 33202
rect 34342 32902 34346 33198
rect 34346 32902 34642 33198
rect 34642 32902 34646 33198
rect 34342 32898 34646 32902
rect 10002 32858 10306 32862
rect 10002 32242 10006 32858
rect 10006 32242 10302 32858
rect 10302 32242 10306 32858
rect 10002 32238 10306 32242
rect 11002 32858 11306 32862
rect 11002 32242 11006 32858
rect 11006 32242 11302 32858
rect 11302 32242 11306 32858
rect 11002 32238 11306 32242
rect 12002 32858 12306 32862
rect 12002 32242 12006 32858
rect 12006 32242 12302 32858
rect 12302 32242 12306 32858
rect 12002 32238 12306 32242
rect 13002 32858 13306 32862
rect 13002 32242 13006 32858
rect 13006 32242 13302 32858
rect 13302 32242 13306 32858
rect 13002 32238 13306 32242
rect 14002 32858 14306 32862
rect 14002 32242 14006 32858
rect 14006 32242 14302 32858
rect 14302 32242 14306 32858
rect 14002 32238 14306 32242
rect 15002 32858 15306 32862
rect 15002 32242 15006 32858
rect 15006 32242 15302 32858
rect 15302 32242 15306 32858
rect 15002 32238 15306 32242
rect 16002 32858 16306 32862
rect 16002 32242 16006 32858
rect 16006 32242 16302 32858
rect 16302 32242 16306 32858
rect 16002 32238 16306 32242
rect 17002 32858 17306 32862
rect 17002 32242 17006 32858
rect 17006 32242 17302 32858
rect 17302 32242 17306 32858
rect 17002 32238 17306 32242
rect 18002 32858 18306 32862
rect 18002 32242 18006 32858
rect 18006 32242 18302 32858
rect 18302 32242 18306 32858
rect 18002 32238 18306 32242
rect 19002 32858 19306 32862
rect 19002 32242 19006 32858
rect 19006 32242 19302 32858
rect 19302 32242 19306 32858
rect 19002 32238 19306 32242
rect 20002 32858 20306 32862
rect 20002 32242 20006 32858
rect 20006 32242 20302 32858
rect 20302 32242 20306 32858
rect 20002 32238 20306 32242
rect 21002 32858 21306 32862
rect 21002 32242 21006 32858
rect 21006 32242 21302 32858
rect 21302 32242 21306 32858
rect 21002 32238 21306 32242
rect 22002 32858 22306 32862
rect 22002 32242 22006 32858
rect 22006 32242 22302 32858
rect 22302 32242 22306 32858
rect 22002 32238 22306 32242
rect 23002 32858 23306 32862
rect 23002 32242 23006 32858
rect 23006 32242 23302 32858
rect 23302 32242 23306 32858
rect 23002 32238 23306 32242
rect 24002 32858 24306 32862
rect 24002 32242 24006 32858
rect 24006 32242 24302 32858
rect 24302 32242 24306 32858
rect 24002 32238 24306 32242
rect 25002 32858 25306 32862
rect 25002 32242 25006 32858
rect 25006 32242 25302 32858
rect 25302 32242 25306 32858
rect 25002 32238 25306 32242
rect 26002 32858 26306 32862
rect 26002 32242 26006 32858
rect 26006 32242 26302 32858
rect 26302 32242 26306 32858
rect 26002 32238 26306 32242
rect 27002 32858 27306 32862
rect 27002 32242 27006 32858
rect 27006 32242 27302 32858
rect 27302 32242 27306 32858
rect 27002 32238 27306 32242
rect 28002 32858 28306 32862
rect 28002 32242 28006 32858
rect 28006 32242 28302 32858
rect 28302 32242 28306 32858
rect 28002 32238 28306 32242
rect 29002 32858 29306 32862
rect 29002 32242 29006 32858
rect 29006 32242 29302 32858
rect 29302 32242 29306 32858
rect 29002 32238 29306 32242
rect 30002 32858 30306 32862
rect 30002 32242 30006 32858
rect 30006 32242 30302 32858
rect 30302 32242 30306 32858
rect 30002 32238 30306 32242
rect 31002 32858 31306 32862
rect 31002 32242 31006 32858
rect 31006 32242 31302 32858
rect 31302 32242 31306 32858
rect 31002 32238 31306 32242
rect 32002 32858 32306 32862
rect 32002 32242 32006 32858
rect 32006 32242 32302 32858
rect 32302 32242 32306 32858
rect 32002 32238 32306 32242
rect 33002 32858 33306 32862
rect 33002 32242 33006 32858
rect 33006 32242 33302 32858
rect 33302 32242 33306 32858
rect 33002 32238 33306 32242
rect 34002 32858 34306 32862
rect 34002 32242 34006 32858
rect 34006 32242 34302 32858
rect 34302 32242 34306 32858
rect 34002 32238 34306 32242
rect -74817 32198 -74513 32202
rect -74817 31902 -74813 32198
rect -74813 31902 -74517 32198
rect -74517 31902 -74513 32198
rect -74817 31898 -74513 31902
rect -74477 32198 -74173 32202
rect -74477 31902 -74473 32198
rect -74473 31902 -74177 32198
rect -74177 31902 -74173 32198
rect -74477 31898 -74173 31902
rect -74137 32198 -73513 32202
rect -74137 31902 -74133 32198
rect -74133 31902 -73517 32198
rect -73517 31902 -73513 32198
rect -74137 31898 -73513 31902
rect -73477 32198 -73173 32202
rect -73477 31902 -73473 32198
rect -73473 31902 -73177 32198
rect -73177 31902 -73173 32198
rect -73477 31898 -73173 31902
rect -73137 32198 -72513 32202
rect -73137 31902 -73133 32198
rect -73133 31902 -72517 32198
rect -72517 31902 -72513 32198
rect -73137 31898 -72513 31902
rect -72477 32198 -72173 32202
rect -72477 31902 -72473 32198
rect -72473 31902 -72177 32198
rect -72177 31902 -72173 32198
rect -72477 31898 -72173 31902
rect -72137 32198 -71513 32202
rect -72137 31902 -72133 32198
rect -72133 31902 -71517 32198
rect -71517 31902 -71513 32198
rect -72137 31898 -71513 31902
rect -71477 32198 -71173 32202
rect -71477 31902 -71473 32198
rect -71473 31902 -71177 32198
rect -71177 31902 -71173 32198
rect -71477 31898 -71173 31902
rect -71137 32198 -70513 32202
rect -71137 31902 -71133 32198
rect -71133 31902 -70517 32198
rect -70517 31902 -70513 32198
rect -71137 31898 -70513 31902
rect -70477 32198 -70173 32202
rect -70477 31902 -70473 32198
rect -70473 31902 -70177 32198
rect -70177 31902 -70173 32198
rect -70477 31898 -70173 31902
rect -70137 32198 -69513 32202
rect -70137 31902 -70133 32198
rect -70133 31902 -69517 32198
rect -69517 31902 -69513 32198
rect -70137 31898 -69513 31902
rect -69477 32198 -69173 32202
rect -69477 31902 -69473 32198
rect -69473 31902 -69177 32198
rect -69177 31902 -69173 32198
rect -69477 31898 -69173 31902
rect -69137 32198 -68513 32202
rect -69137 31902 -69133 32198
rect -69133 31902 -68517 32198
rect -68517 31902 -68513 32198
rect -69137 31898 -68513 31902
rect -68477 32198 -68173 32202
rect -68477 31902 -68473 32198
rect -68473 31902 -68177 32198
rect -68177 31902 -68173 32198
rect -68477 31898 -68173 31902
rect -68137 32198 -67513 32202
rect -68137 31902 -68133 32198
rect -68133 31902 -67517 32198
rect -67517 31902 -67513 32198
rect -68137 31898 -67513 31902
rect -67477 32198 -67173 32202
rect -67477 31902 -67473 32198
rect -67473 31902 -67177 32198
rect -67177 31902 -67173 32198
rect -67477 31898 -67173 31902
rect -67137 32198 -66513 32202
rect -67137 31902 -67133 32198
rect -67133 31902 -66517 32198
rect -66517 31902 -66513 32198
rect -67137 31898 -66513 31902
rect -66477 32198 -66173 32202
rect -66477 31902 -66473 32198
rect -66473 31902 -66177 32198
rect -66177 31902 -66173 32198
rect -66477 31898 -66173 31902
rect -66137 32198 -65513 32202
rect -66137 31902 -66133 32198
rect -66133 31902 -65517 32198
rect -65517 31902 -65513 32198
rect -66137 31898 -65513 31902
rect -65477 32198 -65173 32202
rect -65477 31902 -65473 32198
rect -65473 31902 -65177 32198
rect -65177 31902 -65173 32198
rect -65477 31898 -65173 31902
rect -65137 32198 -64513 32202
rect -65137 31902 -65133 32198
rect -65133 31902 -64517 32198
rect -64517 31902 -64513 32198
rect -65137 31898 -64513 31902
rect -64477 32198 -64173 32202
rect -64477 31902 -64473 32198
rect -64473 31902 -64177 32198
rect -64177 31902 -64173 32198
rect -64477 31898 -64173 31902
rect -64137 32198 -63513 32202
rect -64137 31902 -64133 32198
rect -64133 31902 -63517 32198
rect -63517 31902 -63513 32198
rect -64137 31898 -63513 31902
rect -63477 32198 -63173 32202
rect -63477 31902 -63473 32198
rect -63473 31902 -63177 32198
rect -63177 31902 -63173 32198
rect -63477 31898 -63173 31902
rect -63137 32198 -62513 32202
rect -63137 31902 -63133 32198
rect -63133 31902 -62517 32198
rect -62517 31902 -62513 32198
rect -63137 31898 -62513 31902
rect -62477 32198 -62173 32202
rect -62477 31902 -62473 32198
rect -62473 31902 -62177 32198
rect -62177 31902 -62173 32198
rect -62477 31898 -62173 31902
rect -62137 32198 -61513 32202
rect -62137 31902 -62133 32198
rect -62133 31902 -61517 32198
rect -61517 31902 -61513 32198
rect -62137 31898 -61513 31902
rect -61477 32198 -61173 32202
rect -61477 31902 -61473 32198
rect -61473 31902 -61177 32198
rect -61177 31902 -61173 32198
rect -61477 31898 -61173 31902
rect -61137 32198 -60513 32202
rect -61137 31902 -61133 32198
rect -61133 31902 -60517 32198
rect -60517 31902 -60513 32198
rect -61137 31898 -60513 31902
rect -60477 32198 -60173 32202
rect -60477 31902 -60473 32198
rect -60473 31902 -60177 32198
rect -60177 31902 -60173 32198
rect -60477 31898 -60173 31902
rect -60137 32198 -59513 32202
rect -60137 31902 -60133 32198
rect -60133 31902 -59517 32198
rect -59517 31902 -59513 32198
rect -60137 31898 -59513 31902
rect -59477 32198 -59173 32202
rect -59477 31902 -59473 32198
rect -59473 31902 -59177 32198
rect -59177 31902 -59173 32198
rect -59477 31898 -59173 31902
rect -59137 32198 -58833 32202
rect -59137 31902 -59133 32198
rect -59133 31902 -58837 32198
rect -58837 31902 -58833 32198
rect -59137 31898 -58833 31902
rect 9662 32198 9966 32202
rect 9662 31902 9666 32198
rect 9666 31902 9962 32198
rect 9962 31902 9966 32198
rect 9662 31898 9966 31902
rect 10002 32198 10306 32202
rect 10002 31902 10006 32198
rect 10006 31902 10302 32198
rect 10302 31902 10306 32198
rect 10002 31898 10306 31902
rect 10342 32198 10966 32202
rect 10342 31902 10346 32198
rect 10346 31902 10962 32198
rect 10962 31902 10966 32198
rect 10342 31898 10966 31902
rect 11002 32198 11306 32202
rect 11002 31902 11006 32198
rect 11006 31902 11302 32198
rect 11302 31902 11306 32198
rect 11002 31898 11306 31902
rect 11342 32198 11966 32202
rect 11342 31902 11346 32198
rect 11346 31902 11962 32198
rect 11962 31902 11966 32198
rect 11342 31898 11966 31902
rect 12002 32198 12306 32202
rect 12002 31902 12006 32198
rect 12006 31902 12302 32198
rect 12302 31902 12306 32198
rect 12002 31898 12306 31902
rect 12342 32198 12966 32202
rect 12342 31902 12346 32198
rect 12346 31902 12962 32198
rect 12962 31902 12966 32198
rect 12342 31898 12966 31902
rect 13002 32198 13306 32202
rect 13002 31902 13006 32198
rect 13006 31902 13302 32198
rect 13302 31902 13306 32198
rect 13002 31898 13306 31902
rect 13342 32198 13966 32202
rect 13342 31902 13346 32198
rect 13346 31902 13962 32198
rect 13962 31902 13966 32198
rect 13342 31898 13966 31902
rect 14002 32198 14306 32202
rect 14002 31902 14006 32198
rect 14006 31902 14302 32198
rect 14302 31902 14306 32198
rect 14002 31898 14306 31902
rect 14342 32198 14966 32202
rect 14342 31902 14346 32198
rect 14346 31902 14962 32198
rect 14962 31902 14966 32198
rect 14342 31898 14966 31902
rect 15002 32198 15306 32202
rect 15002 31902 15006 32198
rect 15006 31902 15302 32198
rect 15302 31902 15306 32198
rect 15002 31898 15306 31902
rect 15342 32198 15966 32202
rect 15342 31902 15346 32198
rect 15346 31902 15962 32198
rect 15962 31902 15966 32198
rect 15342 31898 15966 31902
rect 16002 32198 16306 32202
rect 16002 31902 16006 32198
rect 16006 31902 16302 32198
rect 16302 31902 16306 32198
rect 16002 31898 16306 31902
rect 16342 32198 16966 32202
rect 16342 31902 16346 32198
rect 16346 31902 16962 32198
rect 16962 31902 16966 32198
rect 16342 31898 16966 31902
rect 17002 32198 17306 32202
rect 17002 31902 17006 32198
rect 17006 31902 17302 32198
rect 17302 31902 17306 32198
rect 17002 31898 17306 31902
rect 17342 32198 17966 32202
rect 17342 31902 17346 32198
rect 17346 31902 17962 32198
rect 17962 31902 17966 32198
rect 17342 31898 17966 31902
rect 18002 32198 18306 32202
rect 18002 31902 18006 32198
rect 18006 31902 18302 32198
rect 18302 31902 18306 32198
rect 18002 31898 18306 31902
rect 18342 32198 18966 32202
rect 18342 31902 18346 32198
rect 18346 31902 18962 32198
rect 18962 31902 18966 32198
rect 18342 31898 18966 31902
rect 19002 32198 19306 32202
rect 19002 31902 19006 32198
rect 19006 31902 19302 32198
rect 19302 31902 19306 32198
rect 19002 31898 19306 31902
rect 19342 32198 19966 32202
rect 19342 31902 19346 32198
rect 19346 31902 19962 32198
rect 19962 31902 19966 32198
rect 19342 31898 19966 31902
rect 20002 32198 20306 32202
rect 20002 31902 20006 32198
rect 20006 31902 20302 32198
rect 20302 31902 20306 32198
rect 20002 31898 20306 31902
rect 20342 32198 20966 32202
rect 20342 31902 20346 32198
rect 20346 31902 20962 32198
rect 20962 31902 20966 32198
rect 20342 31898 20966 31902
rect 21002 32198 21306 32202
rect 21002 31902 21006 32198
rect 21006 31902 21302 32198
rect 21302 31902 21306 32198
rect 21002 31898 21306 31902
rect 21342 32198 21966 32202
rect 21342 31902 21346 32198
rect 21346 31902 21962 32198
rect 21962 31902 21966 32198
rect 21342 31898 21966 31902
rect 22002 32198 22306 32202
rect 22002 31902 22006 32198
rect 22006 31902 22302 32198
rect 22302 31902 22306 32198
rect 22002 31898 22306 31902
rect 22342 32198 22966 32202
rect 22342 31902 22346 32198
rect 22346 31902 22962 32198
rect 22962 31902 22966 32198
rect 22342 31898 22966 31902
rect 23002 32198 23306 32202
rect 23002 31902 23006 32198
rect 23006 31902 23302 32198
rect 23302 31902 23306 32198
rect 23002 31898 23306 31902
rect 23342 32198 23966 32202
rect 23342 31902 23346 32198
rect 23346 31902 23962 32198
rect 23962 31902 23966 32198
rect 23342 31898 23966 31902
rect 24002 32198 24306 32202
rect 24002 31902 24006 32198
rect 24006 31902 24302 32198
rect 24302 31902 24306 32198
rect 24002 31898 24306 31902
rect 24342 32198 24966 32202
rect 24342 31902 24346 32198
rect 24346 31902 24962 32198
rect 24962 31902 24966 32198
rect 24342 31898 24966 31902
rect 25002 32198 25306 32202
rect 25002 31902 25006 32198
rect 25006 31902 25302 32198
rect 25302 31902 25306 32198
rect 25002 31898 25306 31902
rect 25342 32198 25966 32202
rect 25342 31902 25346 32198
rect 25346 31902 25962 32198
rect 25962 31902 25966 32198
rect 25342 31898 25966 31902
rect 26002 32198 26306 32202
rect 26002 31902 26006 32198
rect 26006 31902 26302 32198
rect 26302 31902 26306 32198
rect 26002 31898 26306 31902
rect 26342 32198 26966 32202
rect 26342 31902 26346 32198
rect 26346 31902 26962 32198
rect 26962 31902 26966 32198
rect 26342 31898 26966 31902
rect 27002 32198 27306 32202
rect 27002 31902 27006 32198
rect 27006 31902 27302 32198
rect 27302 31902 27306 32198
rect 27002 31898 27306 31902
rect 27342 32198 27966 32202
rect 27342 31902 27346 32198
rect 27346 31902 27962 32198
rect 27962 31902 27966 32198
rect 27342 31898 27966 31902
rect 28002 32198 28306 32202
rect 28002 31902 28006 32198
rect 28006 31902 28302 32198
rect 28302 31902 28306 32198
rect 28002 31898 28306 31902
rect 28342 32198 28966 32202
rect 28342 31902 28346 32198
rect 28346 31902 28962 32198
rect 28962 31902 28966 32198
rect 28342 31898 28966 31902
rect 29002 32198 29306 32202
rect 29002 31902 29006 32198
rect 29006 31902 29302 32198
rect 29302 31902 29306 32198
rect 29002 31898 29306 31902
rect 29342 32198 29966 32202
rect 29342 31902 29346 32198
rect 29346 31902 29962 32198
rect 29962 31902 29966 32198
rect 29342 31898 29966 31902
rect 30002 32198 30306 32202
rect 30002 31902 30006 32198
rect 30006 31902 30302 32198
rect 30302 31902 30306 32198
rect 30002 31898 30306 31902
rect 30342 32198 30966 32202
rect 30342 31902 30346 32198
rect 30346 31902 30962 32198
rect 30962 31902 30966 32198
rect 30342 31898 30966 31902
rect 31002 32198 31306 32202
rect 31002 31902 31006 32198
rect 31006 31902 31302 32198
rect 31302 31902 31306 32198
rect 31002 31898 31306 31902
rect 31342 32198 31966 32202
rect 31342 31902 31346 32198
rect 31346 31902 31962 32198
rect 31962 31902 31966 32198
rect 31342 31898 31966 31902
rect 32002 32198 32306 32202
rect 32002 31902 32006 32198
rect 32006 31902 32302 32198
rect 32302 31902 32306 32198
rect 32002 31898 32306 31902
rect 32342 32198 32966 32202
rect 32342 31902 32346 32198
rect 32346 31902 32962 32198
rect 32962 31902 32966 32198
rect 32342 31898 32966 31902
rect 33002 32198 33306 32202
rect 33002 31902 33006 32198
rect 33006 31902 33302 32198
rect 33302 31902 33306 32198
rect 33002 31898 33306 31902
rect 33342 32198 33966 32202
rect 33342 31902 33346 32198
rect 33346 31902 33962 32198
rect 33962 31902 33966 32198
rect 33342 31898 33966 31902
rect 34002 32198 34306 32202
rect 34002 31902 34006 32198
rect 34006 31902 34302 32198
rect 34302 31902 34306 32198
rect 34002 31898 34306 31902
rect 34342 32198 34646 32202
rect 34342 31902 34346 32198
rect 34346 31902 34642 32198
rect 34642 31902 34646 32198
rect 34342 31898 34646 31902
rect -74477 31858 -74173 31862
rect -74477 31242 -74473 31858
rect -74473 31242 -74177 31858
rect -74177 31242 -74173 31858
rect -74477 31238 -74173 31242
rect -73477 31858 -73173 31862
rect -73477 31242 -73473 31858
rect -73473 31242 -73177 31858
rect -73177 31242 -73173 31858
rect -73477 31238 -73173 31242
rect -72477 31858 -72173 31862
rect -72477 31242 -72473 31858
rect -72473 31242 -72177 31858
rect -72177 31242 -72173 31858
rect -72477 31238 -72173 31242
rect -71477 31858 -71173 31862
rect -71477 31242 -71473 31858
rect -71473 31242 -71177 31858
rect -71177 31242 -71173 31858
rect -71477 31238 -71173 31242
rect -70477 31858 -70173 31862
rect -70477 31242 -70473 31858
rect -70473 31242 -70177 31858
rect -70177 31242 -70173 31858
rect -70477 31238 -70173 31242
rect -69477 31858 -69173 31862
rect -69477 31242 -69473 31858
rect -69473 31242 -69177 31858
rect -69177 31242 -69173 31858
rect -69477 31238 -69173 31242
rect -68477 31858 -68173 31862
rect -68477 31242 -68473 31858
rect -68473 31242 -68177 31858
rect -68177 31242 -68173 31858
rect -68477 31238 -68173 31242
rect -67477 31858 -67173 31862
rect -67477 31242 -67473 31858
rect -67473 31242 -67177 31858
rect -67177 31242 -67173 31858
rect -67477 31238 -67173 31242
rect -66477 31858 -66173 31862
rect -66477 31242 -66473 31858
rect -66473 31242 -66177 31858
rect -66177 31242 -66173 31858
rect -66477 31238 -66173 31242
rect -65477 31858 -65173 31862
rect -65477 31242 -65473 31858
rect -65473 31242 -65177 31858
rect -65177 31242 -65173 31858
rect -65477 31238 -65173 31242
rect -64477 31858 -64173 31862
rect -64477 31242 -64473 31858
rect -64473 31242 -64177 31858
rect -64177 31242 -64173 31858
rect -64477 31238 -64173 31242
rect -63477 31858 -63173 31862
rect -63477 31242 -63473 31858
rect -63473 31242 -63177 31858
rect -63177 31242 -63173 31858
rect -63477 31238 -63173 31242
rect -62477 31858 -62173 31862
rect -62477 31242 -62473 31858
rect -62473 31242 -62177 31858
rect -62177 31242 -62173 31858
rect -62477 31238 -62173 31242
rect -61477 31858 -61173 31862
rect -61477 31242 -61473 31858
rect -61473 31242 -61177 31858
rect -61177 31242 -61173 31858
rect -61477 31238 -61173 31242
rect -60477 31858 -60173 31862
rect -60477 31242 -60473 31858
rect -60473 31242 -60177 31858
rect -60177 31242 -60173 31858
rect -60477 31238 -60173 31242
rect -59477 31858 -59173 31862
rect -59477 31242 -59473 31858
rect -59473 31242 -59177 31858
rect -59177 31242 -59173 31858
rect -59477 31238 -59173 31242
rect 10002 31858 10306 31862
rect 10002 31242 10006 31858
rect 10006 31242 10302 31858
rect 10302 31242 10306 31858
rect 10002 31238 10306 31242
rect 11002 31858 11306 31862
rect 11002 31242 11006 31858
rect 11006 31242 11302 31858
rect 11302 31242 11306 31858
rect 11002 31238 11306 31242
rect 12002 31858 12306 31862
rect 12002 31242 12006 31858
rect 12006 31242 12302 31858
rect 12302 31242 12306 31858
rect 12002 31238 12306 31242
rect 13002 31858 13306 31862
rect 13002 31242 13006 31858
rect 13006 31242 13302 31858
rect 13302 31242 13306 31858
rect 13002 31238 13306 31242
rect 14002 31858 14306 31862
rect 14002 31242 14006 31858
rect 14006 31242 14302 31858
rect 14302 31242 14306 31858
rect 14002 31238 14306 31242
rect 15002 31858 15306 31862
rect 15002 31242 15006 31858
rect 15006 31242 15302 31858
rect 15302 31242 15306 31858
rect 15002 31238 15306 31242
rect 16002 31858 16306 31862
rect 16002 31242 16006 31858
rect 16006 31242 16302 31858
rect 16302 31242 16306 31858
rect 16002 31238 16306 31242
rect 17002 31858 17306 31862
rect 17002 31242 17006 31858
rect 17006 31242 17302 31858
rect 17302 31242 17306 31858
rect 17002 31238 17306 31242
rect 18002 31858 18306 31862
rect 18002 31242 18006 31858
rect 18006 31242 18302 31858
rect 18302 31242 18306 31858
rect 18002 31238 18306 31242
rect 19002 31858 19306 31862
rect 19002 31242 19006 31858
rect 19006 31242 19302 31858
rect 19302 31242 19306 31858
rect 19002 31238 19306 31242
rect 20002 31858 20306 31862
rect 20002 31242 20006 31858
rect 20006 31242 20302 31858
rect 20302 31242 20306 31858
rect 20002 31238 20306 31242
rect 21002 31858 21306 31862
rect 21002 31242 21006 31858
rect 21006 31242 21302 31858
rect 21302 31242 21306 31858
rect 21002 31238 21306 31242
rect 22002 31858 22306 31862
rect 22002 31242 22006 31858
rect 22006 31242 22302 31858
rect 22302 31242 22306 31858
rect 22002 31238 22306 31242
rect 23002 31858 23306 31862
rect 23002 31242 23006 31858
rect 23006 31242 23302 31858
rect 23302 31242 23306 31858
rect 23002 31238 23306 31242
rect 24002 31858 24306 31862
rect 24002 31242 24006 31858
rect 24006 31242 24302 31858
rect 24302 31242 24306 31858
rect 24002 31238 24306 31242
rect 25002 31858 25306 31862
rect 25002 31242 25006 31858
rect 25006 31242 25302 31858
rect 25302 31242 25306 31858
rect 25002 31238 25306 31242
rect 26002 31858 26306 31862
rect 26002 31242 26006 31858
rect 26006 31242 26302 31858
rect 26302 31242 26306 31858
rect 26002 31238 26306 31242
rect 27002 31858 27306 31862
rect 27002 31242 27006 31858
rect 27006 31242 27302 31858
rect 27302 31242 27306 31858
rect 27002 31238 27306 31242
rect 28002 31858 28306 31862
rect 28002 31242 28006 31858
rect 28006 31242 28302 31858
rect 28302 31242 28306 31858
rect 28002 31238 28306 31242
rect 29002 31858 29306 31862
rect 29002 31242 29006 31858
rect 29006 31242 29302 31858
rect 29302 31242 29306 31858
rect 29002 31238 29306 31242
rect 30002 31858 30306 31862
rect 30002 31242 30006 31858
rect 30006 31242 30302 31858
rect 30302 31242 30306 31858
rect 30002 31238 30306 31242
rect 31002 31858 31306 31862
rect 31002 31242 31006 31858
rect 31006 31242 31302 31858
rect 31302 31242 31306 31858
rect 31002 31238 31306 31242
rect 32002 31858 32306 31862
rect 32002 31242 32006 31858
rect 32006 31242 32302 31858
rect 32302 31242 32306 31858
rect 32002 31238 32306 31242
rect 33002 31858 33306 31862
rect 33002 31242 33006 31858
rect 33006 31242 33302 31858
rect 33302 31242 33306 31858
rect 33002 31238 33306 31242
rect 34002 31858 34306 31862
rect 34002 31242 34006 31858
rect 34006 31242 34302 31858
rect 34302 31242 34306 31858
rect 34002 31238 34306 31242
rect -74817 31198 -74513 31202
rect -74817 30902 -74813 31198
rect -74813 30902 -74517 31198
rect -74517 30902 -74513 31198
rect -74817 30898 -74513 30902
rect -74477 31198 -74173 31202
rect -74477 30902 -74473 31198
rect -74473 30902 -74177 31198
rect -74177 30902 -74173 31198
rect -74477 30898 -74173 30902
rect -74137 31198 -73513 31202
rect -74137 30902 -74133 31198
rect -74133 30902 -73517 31198
rect -73517 30902 -73513 31198
rect -74137 30898 -73513 30902
rect -73477 31198 -73173 31202
rect -73477 30902 -73473 31198
rect -73473 30902 -73177 31198
rect -73177 30902 -73173 31198
rect -73477 30898 -73173 30902
rect -73137 31198 -72513 31202
rect -73137 30902 -73133 31198
rect -73133 30902 -72517 31198
rect -72517 30902 -72513 31198
rect -73137 30898 -72513 30902
rect -72477 31198 -72173 31202
rect -72477 30902 -72473 31198
rect -72473 30902 -72177 31198
rect -72177 30902 -72173 31198
rect -72477 30898 -72173 30902
rect -72137 31198 -71513 31202
rect -72137 30902 -72133 31198
rect -72133 30902 -71517 31198
rect -71517 30902 -71513 31198
rect -72137 30898 -71513 30902
rect -71477 31198 -71173 31202
rect -71477 30902 -71473 31198
rect -71473 30902 -71177 31198
rect -71177 30902 -71173 31198
rect -71477 30898 -71173 30902
rect -71137 31198 -70513 31202
rect -71137 30902 -71133 31198
rect -71133 30902 -70517 31198
rect -70517 30902 -70513 31198
rect -71137 30898 -70513 30902
rect -70477 31198 -70173 31202
rect -70477 30902 -70473 31198
rect -70473 30902 -70177 31198
rect -70177 30902 -70173 31198
rect -70477 30898 -70173 30902
rect -70137 31198 -69513 31202
rect -70137 30902 -70133 31198
rect -70133 30902 -69517 31198
rect -69517 30902 -69513 31198
rect -70137 30898 -69513 30902
rect -69477 31198 -69173 31202
rect -69477 30902 -69473 31198
rect -69473 30902 -69177 31198
rect -69177 30902 -69173 31198
rect -69477 30898 -69173 30902
rect -69137 31198 -68513 31202
rect -69137 30902 -69133 31198
rect -69133 30902 -68517 31198
rect -68517 30902 -68513 31198
rect -69137 30898 -68513 30902
rect -68477 31198 -68173 31202
rect -68477 30902 -68473 31198
rect -68473 30902 -68177 31198
rect -68177 30902 -68173 31198
rect -68477 30898 -68173 30902
rect -68137 31198 -67513 31202
rect -68137 30902 -68133 31198
rect -68133 30902 -67517 31198
rect -67517 30902 -67513 31198
rect -68137 30898 -67513 30902
rect -67477 31198 -67173 31202
rect -67477 30902 -67473 31198
rect -67473 30902 -67177 31198
rect -67177 30902 -67173 31198
rect -67477 30898 -67173 30902
rect -67137 31198 -66513 31202
rect -67137 30902 -67133 31198
rect -67133 30902 -66517 31198
rect -66517 30902 -66513 31198
rect -67137 30898 -66513 30902
rect -66477 31198 -66173 31202
rect -66477 30902 -66473 31198
rect -66473 30902 -66177 31198
rect -66177 30902 -66173 31198
rect -66477 30898 -66173 30902
rect -66137 31198 -65513 31202
rect -66137 30902 -66133 31198
rect -66133 30902 -65517 31198
rect -65517 30902 -65513 31198
rect -66137 30898 -65513 30902
rect -65477 31198 -65173 31202
rect -65477 30902 -65473 31198
rect -65473 30902 -65177 31198
rect -65177 30902 -65173 31198
rect -65477 30898 -65173 30902
rect -65137 31198 -64513 31202
rect -65137 30902 -65133 31198
rect -65133 30902 -64517 31198
rect -64517 30902 -64513 31198
rect -65137 30898 -64513 30902
rect -64477 31198 -64173 31202
rect -64477 30902 -64473 31198
rect -64473 30902 -64177 31198
rect -64177 30902 -64173 31198
rect -64477 30898 -64173 30902
rect -64137 31198 -63513 31202
rect -64137 30902 -64133 31198
rect -64133 30902 -63517 31198
rect -63517 30902 -63513 31198
rect -64137 30898 -63513 30902
rect -63477 31198 -63173 31202
rect -63477 30902 -63473 31198
rect -63473 30902 -63177 31198
rect -63177 30902 -63173 31198
rect -63477 30898 -63173 30902
rect -63137 31198 -62513 31202
rect -63137 30902 -63133 31198
rect -63133 30902 -62517 31198
rect -62517 30902 -62513 31198
rect -63137 30898 -62513 30902
rect -62477 31198 -62173 31202
rect -62477 30902 -62473 31198
rect -62473 30902 -62177 31198
rect -62177 30902 -62173 31198
rect -62477 30898 -62173 30902
rect -62137 31198 -61513 31202
rect -62137 30902 -62133 31198
rect -62133 30902 -61517 31198
rect -61517 30902 -61513 31198
rect -62137 30898 -61513 30902
rect -61477 31198 -61173 31202
rect -61477 30902 -61473 31198
rect -61473 30902 -61177 31198
rect -61177 30902 -61173 31198
rect -61477 30898 -61173 30902
rect -61137 31198 -60513 31202
rect -61137 30902 -61133 31198
rect -61133 30902 -60517 31198
rect -60517 30902 -60513 31198
rect -61137 30898 -60513 30902
rect -60477 31198 -60173 31202
rect -60477 30902 -60473 31198
rect -60473 30902 -60177 31198
rect -60177 30902 -60173 31198
rect -60477 30898 -60173 30902
rect -60137 31198 -59513 31202
rect -60137 30902 -60133 31198
rect -60133 30902 -59517 31198
rect -59517 30902 -59513 31198
rect -60137 30898 -59513 30902
rect -59477 31198 -59173 31202
rect -59477 30902 -59473 31198
rect -59473 30902 -59177 31198
rect -59177 30902 -59173 31198
rect -59477 30898 -59173 30902
rect -59137 31198 -58833 31202
rect -59137 30902 -59133 31198
rect -59133 30902 -58837 31198
rect -58837 30902 -58833 31198
rect -59137 30898 -58833 30902
rect 9662 31198 9966 31202
rect 9662 30902 9666 31198
rect 9666 30902 9962 31198
rect 9962 30902 9966 31198
rect 9662 30898 9966 30902
rect 10002 31198 10306 31202
rect 10002 30902 10006 31198
rect 10006 30902 10302 31198
rect 10302 30902 10306 31198
rect 10002 30898 10306 30902
rect 10342 31198 10966 31202
rect 10342 30902 10346 31198
rect 10346 30902 10962 31198
rect 10962 30902 10966 31198
rect 10342 30898 10966 30902
rect 11002 31198 11306 31202
rect 11002 30902 11006 31198
rect 11006 30902 11302 31198
rect 11302 30902 11306 31198
rect 11002 30898 11306 30902
rect 11342 31198 11966 31202
rect 11342 30902 11346 31198
rect 11346 30902 11962 31198
rect 11962 30902 11966 31198
rect 11342 30898 11966 30902
rect 12002 31198 12306 31202
rect 12002 30902 12006 31198
rect 12006 30902 12302 31198
rect 12302 30902 12306 31198
rect 12002 30898 12306 30902
rect 12342 31198 12966 31202
rect 12342 30902 12346 31198
rect 12346 30902 12962 31198
rect 12962 30902 12966 31198
rect 12342 30898 12966 30902
rect 13002 31198 13306 31202
rect 13002 30902 13006 31198
rect 13006 30902 13302 31198
rect 13302 30902 13306 31198
rect 13002 30898 13306 30902
rect 13342 31198 13966 31202
rect 13342 30902 13346 31198
rect 13346 30902 13962 31198
rect 13962 30902 13966 31198
rect 13342 30898 13966 30902
rect 14002 31198 14306 31202
rect 14002 30902 14006 31198
rect 14006 30902 14302 31198
rect 14302 30902 14306 31198
rect 14002 30898 14306 30902
rect 14342 31198 14966 31202
rect 14342 30902 14346 31198
rect 14346 30902 14962 31198
rect 14962 30902 14966 31198
rect 14342 30898 14966 30902
rect 15002 31198 15306 31202
rect 15002 30902 15006 31198
rect 15006 30902 15302 31198
rect 15302 30902 15306 31198
rect 15002 30898 15306 30902
rect 15342 31198 15966 31202
rect 15342 30902 15346 31198
rect 15346 30902 15962 31198
rect 15962 30902 15966 31198
rect 15342 30898 15966 30902
rect 16002 31198 16306 31202
rect 16002 30902 16006 31198
rect 16006 30902 16302 31198
rect 16302 30902 16306 31198
rect 16002 30898 16306 30902
rect 16342 31198 16966 31202
rect 16342 30902 16346 31198
rect 16346 30902 16962 31198
rect 16962 30902 16966 31198
rect 16342 30898 16966 30902
rect 17002 31198 17306 31202
rect 17002 30902 17006 31198
rect 17006 30902 17302 31198
rect 17302 30902 17306 31198
rect 17002 30898 17306 30902
rect 17342 31198 17966 31202
rect 17342 30902 17346 31198
rect 17346 30902 17962 31198
rect 17962 30902 17966 31198
rect 17342 30898 17966 30902
rect 18002 31198 18306 31202
rect 18002 30902 18006 31198
rect 18006 30902 18302 31198
rect 18302 30902 18306 31198
rect 18002 30898 18306 30902
rect 18342 31198 18966 31202
rect 18342 30902 18346 31198
rect 18346 30902 18962 31198
rect 18962 30902 18966 31198
rect 18342 30898 18966 30902
rect 19002 31198 19306 31202
rect 19002 30902 19006 31198
rect 19006 30902 19302 31198
rect 19302 30902 19306 31198
rect 19002 30898 19306 30902
rect 19342 31198 19966 31202
rect 19342 30902 19346 31198
rect 19346 30902 19962 31198
rect 19962 30902 19966 31198
rect 19342 30898 19966 30902
rect 20002 31198 20306 31202
rect 20002 30902 20006 31198
rect 20006 30902 20302 31198
rect 20302 30902 20306 31198
rect 20002 30898 20306 30902
rect 20342 31198 20966 31202
rect 20342 30902 20346 31198
rect 20346 30902 20962 31198
rect 20962 30902 20966 31198
rect 20342 30898 20966 30902
rect 21002 31198 21306 31202
rect 21002 30902 21006 31198
rect 21006 30902 21302 31198
rect 21302 30902 21306 31198
rect 21002 30898 21306 30902
rect 21342 31198 21966 31202
rect 21342 30902 21346 31198
rect 21346 30902 21962 31198
rect 21962 30902 21966 31198
rect 21342 30898 21966 30902
rect 22002 31198 22306 31202
rect 22002 30902 22006 31198
rect 22006 30902 22302 31198
rect 22302 30902 22306 31198
rect 22002 30898 22306 30902
rect 22342 31198 22966 31202
rect 22342 30902 22346 31198
rect 22346 30902 22962 31198
rect 22962 30902 22966 31198
rect 22342 30898 22966 30902
rect 23002 31198 23306 31202
rect 23002 30902 23006 31198
rect 23006 30902 23302 31198
rect 23302 30902 23306 31198
rect 23002 30898 23306 30902
rect 23342 31198 23966 31202
rect 23342 30902 23346 31198
rect 23346 30902 23962 31198
rect 23962 30902 23966 31198
rect 23342 30898 23966 30902
rect 24002 31198 24306 31202
rect 24002 30902 24006 31198
rect 24006 30902 24302 31198
rect 24302 30902 24306 31198
rect 24002 30898 24306 30902
rect 24342 31198 24966 31202
rect 24342 30902 24346 31198
rect 24346 30902 24962 31198
rect 24962 30902 24966 31198
rect 24342 30898 24966 30902
rect 25002 31198 25306 31202
rect 25002 30902 25006 31198
rect 25006 30902 25302 31198
rect 25302 30902 25306 31198
rect 25002 30898 25306 30902
rect 25342 31198 25966 31202
rect 25342 30902 25346 31198
rect 25346 30902 25962 31198
rect 25962 30902 25966 31198
rect 25342 30898 25966 30902
rect 26002 31198 26306 31202
rect 26002 30902 26006 31198
rect 26006 30902 26302 31198
rect 26302 30902 26306 31198
rect 26002 30898 26306 30902
rect 26342 31198 26966 31202
rect 26342 30902 26346 31198
rect 26346 30902 26962 31198
rect 26962 30902 26966 31198
rect 26342 30898 26966 30902
rect 27002 31198 27306 31202
rect 27002 30902 27006 31198
rect 27006 30902 27302 31198
rect 27302 30902 27306 31198
rect 27002 30898 27306 30902
rect 27342 31198 27966 31202
rect 27342 30902 27346 31198
rect 27346 30902 27962 31198
rect 27962 30902 27966 31198
rect 27342 30898 27966 30902
rect 28002 31198 28306 31202
rect 28002 30902 28006 31198
rect 28006 30902 28302 31198
rect 28302 30902 28306 31198
rect 28002 30898 28306 30902
rect 28342 31198 28966 31202
rect 28342 30902 28346 31198
rect 28346 30902 28962 31198
rect 28962 30902 28966 31198
rect 28342 30898 28966 30902
rect 29002 31198 29306 31202
rect 29002 30902 29006 31198
rect 29006 30902 29302 31198
rect 29302 30902 29306 31198
rect 29002 30898 29306 30902
rect 29342 31198 29966 31202
rect 29342 30902 29346 31198
rect 29346 30902 29962 31198
rect 29962 30902 29966 31198
rect 29342 30898 29966 30902
rect 30002 31198 30306 31202
rect 30002 30902 30006 31198
rect 30006 30902 30302 31198
rect 30302 30902 30306 31198
rect 30002 30898 30306 30902
rect 30342 31198 30966 31202
rect 30342 30902 30346 31198
rect 30346 30902 30962 31198
rect 30962 30902 30966 31198
rect 30342 30898 30966 30902
rect 31002 31198 31306 31202
rect 31002 30902 31006 31198
rect 31006 30902 31302 31198
rect 31302 30902 31306 31198
rect 31002 30898 31306 30902
rect 31342 31198 31966 31202
rect 31342 30902 31346 31198
rect 31346 30902 31962 31198
rect 31962 30902 31966 31198
rect 31342 30898 31966 30902
rect 32002 31198 32306 31202
rect 32002 30902 32006 31198
rect 32006 30902 32302 31198
rect 32302 30902 32306 31198
rect 32002 30898 32306 30902
rect 32342 31198 32966 31202
rect 32342 30902 32346 31198
rect 32346 30902 32962 31198
rect 32962 30902 32966 31198
rect 32342 30898 32966 30902
rect 33002 31198 33306 31202
rect 33002 30902 33006 31198
rect 33006 30902 33302 31198
rect 33302 30902 33306 31198
rect 33002 30898 33306 30902
rect 33342 31198 33966 31202
rect 33342 30902 33346 31198
rect 33346 30902 33962 31198
rect 33962 30902 33966 31198
rect 33342 30898 33966 30902
rect 34002 31198 34306 31202
rect 34002 30902 34006 31198
rect 34006 30902 34302 31198
rect 34302 30902 34306 31198
rect 34002 30898 34306 30902
rect 34342 31198 34646 31202
rect 34342 30902 34346 31198
rect 34346 30902 34642 31198
rect 34642 30902 34646 31198
rect 34342 30898 34646 30902
rect -74477 30858 -74173 30862
rect -74477 30242 -74473 30858
rect -74473 30242 -74177 30858
rect -74177 30242 -74173 30858
rect -74477 30238 -74173 30242
rect -73477 30858 -73173 30862
rect -73477 30242 -73473 30858
rect -73473 30242 -73177 30858
rect -73177 30242 -73173 30858
rect -73477 30238 -73173 30242
rect -72477 30858 -72173 30862
rect -72477 30242 -72473 30858
rect -72473 30242 -72177 30858
rect -72177 30242 -72173 30858
rect -72477 30238 -72173 30242
rect -71477 30858 -71173 30862
rect -71477 30242 -71473 30858
rect -71473 30242 -71177 30858
rect -71177 30242 -71173 30858
rect -71477 30238 -71173 30242
rect -70477 30858 -70173 30862
rect -70477 30242 -70473 30858
rect -70473 30242 -70177 30858
rect -70177 30242 -70173 30858
rect -70477 30238 -70173 30242
rect -69477 30858 -69173 30862
rect -69477 30242 -69473 30858
rect -69473 30242 -69177 30858
rect -69177 30242 -69173 30858
rect -69477 30238 -69173 30242
rect -68477 30858 -68173 30862
rect -68477 30242 -68473 30858
rect -68473 30242 -68177 30858
rect -68177 30242 -68173 30858
rect -68477 30238 -68173 30242
rect -67477 30858 -67173 30862
rect -67477 30242 -67473 30858
rect -67473 30242 -67177 30858
rect -67177 30242 -67173 30858
rect -67477 30238 -67173 30242
rect -66477 30858 -66173 30862
rect -66477 30242 -66473 30858
rect -66473 30242 -66177 30858
rect -66177 30242 -66173 30858
rect -66477 30238 -66173 30242
rect -65477 30858 -65173 30862
rect -65477 30242 -65473 30858
rect -65473 30242 -65177 30858
rect -65177 30242 -65173 30858
rect -65477 30238 -65173 30242
rect -64477 30858 -64173 30862
rect -64477 30242 -64473 30858
rect -64473 30242 -64177 30858
rect -64177 30242 -64173 30858
rect -64477 30238 -64173 30242
rect -63477 30858 -63173 30862
rect -63477 30242 -63473 30858
rect -63473 30242 -63177 30858
rect -63177 30242 -63173 30858
rect -63477 30238 -63173 30242
rect -62477 30858 -62173 30862
rect -62477 30242 -62473 30858
rect -62473 30242 -62177 30858
rect -62177 30242 -62173 30858
rect -62477 30238 -62173 30242
rect -61477 30858 -61173 30862
rect -61477 30242 -61473 30858
rect -61473 30242 -61177 30858
rect -61177 30242 -61173 30858
rect -61477 30238 -61173 30242
rect -60477 30858 -60173 30862
rect -60477 30242 -60473 30858
rect -60473 30242 -60177 30858
rect -60177 30242 -60173 30858
rect -60477 30238 -60173 30242
rect -59477 30858 -59173 30862
rect -59477 30242 -59473 30858
rect -59473 30242 -59177 30858
rect -59177 30242 -59173 30858
rect -59477 30238 -59173 30242
rect 10002 30858 10306 30862
rect 10002 30242 10006 30858
rect 10006 30242 10302 30858
rect 10302 30242 10306 30858
rect 10002 30238 10306 30242
rect 11002 30858 11306 30862
rect 11002 30242 11006 30858
rect 11006 30242 11302 30858
rect 11302 30242 11306 30858
rect 11002 30238 11306 30242
rect 12002 30858 12306 30862
rect 12002 30242 12006 30858
rect 12006 30242 12302 30858
rect 12302 30242 12306 30858
rect 12002 30238 12306 30242
rect 13002 30858 13306 30862
rect 13002 30242 13006 30858
rect 13006 30242 13302 30858
rect 13302 30242 13306 30858
rect 13002 30238 13306 30242
rect 14002 30858 14306 30862
rect 14002 30242 14006 30858
rect 14006 30242 14302 30858
rect 14302 30242 14306 30858
rect 14002 30238 14306 30242
rect 15002 30858 15306 30862
rect 15002 30242 15006 30858
rect 15006 30242 15302 30858
rect 15302 30242 15306 30858
rect 15002 30238 15306 30242
rect 16002 30858 16306 30862
rect 16002 30242 16006 30858
rect 16006 30242 16302 30858
rect 16302 30242 16306 30858
rect 16002 30238 16306 30242
rect 17002 30858 17306 30862
rect 17002 30242 17006 30858
rect 17006 30242 17302 30858
rect 17302 30242 17306 30858
rect 17002 30238 17306 30242
rect 18002 30858 18306 30862
rect 18002 30242 18006 30858
rect 18006 30242 18302 30858
rect 18302 30242 18306 30858
rect 18002 30238 18306 30242
rect 19002 30858 19306 30862
rect 19002 30242 19006 30858
rect 19006 30242 19302 30858
rect 19302 30242 19306 30858
rect 19002 30238 19306 30242
rect 20002 30858 20306 30862
rect 20002 30242 20006 30858
rect 20006 30242 20302 30858
rect 20302 30242 20306 30858
rect 20002 30238 20306 30242
rect 21002 30858 21306 30862
rect 21002 30242 21006 30858
rect 21006 30242 21302 30858
rect 21302 30242 21306 30858
rect 21002 30238 21306 30242
rect 22002 30858 22306 30862
rect 22002 30242 22006 30858
rect 22006 30242 22302 30858
rect 22302 30242 22306 30858
rect 22002 30238 22306 30242
rect 23002 30858 23306 30862
rect 23002 30242 23006 30858
rect 23006 30242 23302 30858
rect 23302 30242 23306 30858
rect 23002 30238 23306 30242
rect 24002 30858 24306 30862
rect 24002 30242 24006 30858
rect 24006 30242 24302 30858
rect 24302 30242 24306 30858
rect 24002 30238 24306 30242
rect 25002 30858 25306 30862
rect 25002 30242 25006 30858
rect 25006 30242 25302 30858
rect 25302 30242 25306 30858
rect 25002 30238 25306 30242
rect 26002 30858 26306 30862
rect 26002 30242 26006 30858
rect 26006 30242 26302 30858
rect 26302 30242 26306 30858
rect 26002 30238 26306 30242
rect 27002 30858 27306 30862
rect 27002 30242 27006 30858
rect 27006 30242 27302 30858
rect 27302 30242 27306 30858
rect 27002 30238 27306 30242
rect 28002 30858 28306 30862
rect 28002 30242 28006 30858
rect 28006 30242 28302 30858
rect 28302 30242 28306 30858
rect 28002 30238 28306 30242
rect 29002 30858 29306 30862
rect 29002 30242 29006 30858
rect 29006 30242 29302 30858
rect 29302 30242 29306 30858
rect 29002 30238 29306 30242
rect 30002 30858 30306 30862
rect 30002 30242 30006 30858
rect 30006 30242 30302 30858
rect 30302 30242 30306 30858
rect 30002 30238 30306 30242
rect 31002 30858 31306 30862
rect 31002 30242 31006 30858
rect 31006 30242 31302 30858
rect 31302 30242 31306 30858
rect 31002 30238 31306 30242
rect 32002 30858 32306 30862
rect 32002 30242 32006 30858
rect 32006 30242 32302 30858
rect 32302 30242 32306 30858
rect 32002 30238 32306 30242
rect 33002 30858 33306 30862
rect 33002 30242 33006 30858
rect 33006 30242 33302 30858
rect 33302 30242 33306 30858
rect 33002 30238 33306 30242
rect 34002 30858 34306 30862
rect 34002 30242 34006 30858
rect 34006 30242 34302 30858
rect 34302 30242 34306 30858
rect 34002 30238 34306 30242
rect -74817 30198 -74513 30202
rect -74817 29902 -74813 30198
rect -74813 29902 -74517 30198
rect -74517 29902 -74513 30198
rect -74817 29898 -74513 29902
rect -74477 30198 -74173 30202
rect -74477 29902 -74473 30198
rect -74473 29902 -74177 30198
rect -74177 29902 -74173 30198
rect -74477 29898 -74173 29902
rect -74137 30198 -73513 30202
rect -74137 29902 -74133 30198
rect -74133 29902 -73517 30198
rect -73517 29902 -73513 30198
rect -74137 29898 -73513 29902
rect -73477 30198 -73173 30202
rect -73477 29902 -73473 30198
rect -73473 29902 -73177 30198
rect -73177 29902 -73173 30198
rect -73477 29898 -73173 29902
rect -73137 30198 -72513 30202
rect -73137 29902 -73133 30198
rect -73133 29902 -72517 30198
rect -72517 29902 -72513 30198
rect -73137 29898 -72513 29902
rect -72477 30198 -72173 30202
rect -72477 29902 -72473 30198
rect -72473 29902 -72177 30198
rect -72177 29902 -72173 30198
rect -72477 29898 -72173 29902
rect -72137 30198 -71513 30202
rect -72137 29902 -72133 30198
rect -72133 29902 -71517 30198
rect -71517 29902 -71513 30198
rect -72137 29898 -71513 29902
rect -71477 30198 -71173 30202
rect -71477 29902 -71473 30198
rect -71473 29902 -71177 30198
rect -71177 29902 -71173 30198
rect -71477 29898 -71173 29902
rect -71137 30198 -70513 30202
rect -71137 29902 -71133 30198
rect -71133 29902 -70517 30198
rect -70517 29902 -70513 30198
rect -71137 29898 -70513 29902
rect -70477 30198 -70173 30202
rect -70477 29902 -70473 30198
rect -70473 29902 -70177 30198
rect -70177 29902 -70173 30198
rect -70477 29898 -70173 29902
rect -70137 30198 -69513 30202
rect -70137 29902 -70133 30198
rect -70133 29902 -69517 30198
rect -69517 29902 -69513 30198
rect -70137 29898 -69513 29902
rect -69477 30198 -69173 30202
rect -69477 29902 -69473 30198
rect -69473 29902 -69177 30198
rect -69177 29902 -69173 30198
rect -69477 29898 -69173 29902
rect -69137 30198 -68513 30202
rect -69137 29902 -69133 30198
rect -69133 29902 -68517 30198
rect -68517 29902 -68513 30198
rect -69137 29898 -68513 29902
rect -68477 30198 -68173 30202
rect -68477 29902 -68473 30198
rect -68473 29902 -68177 30198
rect -68177 29902 -68173 30198
rect -68477 29898 -68173 29902
rect -68137 30198 -67513 30202
rect -68137 29902 -68133 30198
rect -68133 29902 -67517 30198
rect -67517 29902 -67513 30198
rect -68137 29898 -67513 29902
rect -67477 30198 -67173 30202
rect -67477 29902 -67473 30198
rect -67473 29902 -67177 30198
rect -67177 29902 -67173 30198
rect -67477 29898 -67173 29902
rect -67137 30198 -66513 30202
rect -67137 29902 -67133 30198
rect -67133 29902 -66517 30198
rect -66517 29902 -66513 30198
rect -67137 29898 -66513 29902
rect -66477 30198 -66173 30202
rect -66477 29902 -66473 30198
rect -66473 29902 -66177 30198
rect -66177 29902 -66173 30198
rect -66477 29898 -66173 29902
rect -66137 30198 -65513 30202
rect -66137 29902 -66133 30198
rect -66133 29902 -65517 30198
rect -65517 29902 -65513 30198
rect -66137 29898 -65513 29902
rect -65477 30198 -65173 30202
rect -65477 29902 -65473 30198
rect -65473 29902 -65177 30198
rect -65177 29902 -65173 30198
rect -65477 29898 -65173 29902
rect -65137 30198 -64513 30202
rect -65137 29902 -65133 30198
rect -65133 29902 -64517 30198
rect -64517 29902 -64513 30198
rect -65137 29898 -64513 29902
rect -64477 30198 -64173 30202
rect -64477 29902 -64473 30198
rect -64473 29902 -64177 30198
rect -64177 29902 -64173 30198
rect -64477 29898 -64173 29902
rect -64137 30198 -63513 30202
rect -64137 29902 -64133 30198
rect -64133 29902 -63517 30198
rect -63517 29902 -63513 30198
rect -64137 29898 -63513 29902
rect -63477 30198 -63173 30202
rect -63477 29902 -63473 30198
rect -63473 29902 -63177 30198
rect -63177 29902 -63173 30198
rect -63477 29898 -63173 29902
rect -63137 30198 -62513 30202
rect -63137 29902 -63133 30198
rect -63133 29902 -62517 30198
rect -62517 29902 -62513 30198
rect -63137 29898 -62513 29902
rect -62477 30198 -62173 30202
rect -62477 29902 -62473 30198
rect -62473 29902 -62177 30198
rect -62177 29902 -62173 30198
rect -62477 29898 -62173 29902
rect -62137 30198 -61513 30202
rect -62137 29902 -62133 30198
rect -62133 29902 -61517 30198
rect -61517 29902 -61513 30198
rect -62137 29898 -61513 29902
rect -61477 30198 -61173 30202
rect -61477 29902 -61473 30198
rect -61473 29902 -61177 30198
rect -61177 29902 -61173 30198
rect -61477 29898 -61173 29902
rect -61137 30198 -60513 30202
rect -61137 29902 -61133 30198
rect -61133 29902 -60517 30198
rect -60517 29902 -60513 30198
rect -61137 29898 -60513 29902
rect -60477 30198 -60173 30202
rect -60477 29902 -60473 30198
rect -60473 29902 -60177 30198
rect -60177 29902 -60173 30198
rect -60477 29898 -60173 29902
rect -60137 30198 -59513 30202
rect -60137 29902 -60133 30198
rect -60133 29902 -59517 30198
rect -59517 29902 -59513 30198
rect -60137 29898 -59513 29902
rect -59477 30198 -59173 30202
rect -59477 29902 -59473 30198
rect -59473 29902 -59177 30198
rect -59177 29902 -59173 30198
rect -59477 29898 -59173 29902
rect -59137 30198 -58833 30202
rect -59137 29902 -59133 30198
rect -59133 29902 -58837 30198
rect -58837 29902 -58833 30198
rect -59137 29898 -58833 29902
rect 9662 30198 9966 30202
rect 9662 29902 9666 30198
rect 9666 29902 9962 30198
rect 9962 29902 9966 30198
rect 9662 29898 9966 29902
rect 10002 30198 10306 30202
rect 10002 29902 10006 30198
rect 10006 29902 10302 30198
rect 10302 29902 10306 30198
rect 10002 29898 10306 29902
rect 10342 30198 10966 30202
rect 10342 29902 10346 30198
rect 10346 29902 10962 30198
rect 10962 29902 10966 30198
rect 10342 29898 10966 29902
rect 11002 30198 11306 30202
rect 11002 29902 11006 30198
rect 11006 29902 11302 30198
rect 11302 29902 11306 30198
rect 11002 29898 11306 29902
rect 11342 30198 11966 30202
rect 11342 29902 11346 30198
rect 11346 29902 11962 30198
rect 11962 29902 11966 30198
rect 11342 29898 11966 29902
rect 12002 30198 12306 30202
rect 12002 29902 12006 30198
rect 12006 29902 12302 30198
rect 12302 29902 12306 30198
rect 12002 29898 12306 29902
rect 12342 30198 12966 30202
rect 12342 29902 12346 30198
rect 12346 29902 12962 30198
rect 12962 29902 12966 30198
rect 12342 29898 12966 29902
rect 13002 30198 13306 30202
rect 13002 29902 13006 30198
rect 13006 29902 13302 30198
rect 13302 29902 13306 30198
rect 13002 29898 13306 29902
rect 13342 30198 13966 30202
rect 13342 29902 13346 30198
rect 13346 29902 13962 30198
rect 13962 29902 13966 30198
rect 13342 29898 13966 29902
rect 14002 30198 14306 30202
rect 14002 29902 14006 30198
rect 14006 29902 14302 30198
rect 14302 29902 14306 30198
rect 14002 29898 14306 29902
rect 14342 30198 14966 30202
rect 14342 29902 14346 30198
rect 14346 29902 14962 30198
rect 14962 29902 14966 30198
rect 14342 29898 14966 29902
rect 15002 30198 15306 30202
rect 15002 29902 15006 30198
rect 15006 29902 15302 30198
rect 15302 29902 15306 30198
rect 15002 29898 15306 29902
rect 15342 30198 15966 30202
rect 15342 29902 15346 30198
rect 15346 29902 15962 30198
rect 15962 29902 15966 30198
rect 15342 29898 15966 29902
rect 16002 30198 16306 30202
rect 16002 29902 16006 30198
rect 16006 29902 16302 30198
rect 16302 29902 16306 30198
rect 16002 29898 16306 29902
rect 16342 30198 16966 30202
rect 16342 29902 16346 30198
rect 16346 29902 16962 30198
rect 16962 29902 16966 30198
rect 16342 29898 16966 29902
rect 17002 30198 17306 30202
rect 17002 29902 17006 30198
rect 17006 29902 17302 30198
rect 17302 29902 17306 30198
rect 17002 29898 17306 29902
rect 17342 30198 17966 30202
rect 17342 29902 17346 30198
rect 17346 29902 17962 30198
rect 17962 29902 17966 30198
rect 17342 29898 17966 29902
rect 18002 30198 18306 30202
rect 18002 29902 18006 30198
rect 18006 29902 18302 30198
rect 18302 29902 18306 30198
rect 18002 29898 18306 29902
rect 18342 30198 18966 30202
rect 18342 29902 18346 30198
rect 18346 29902 18962 30198
rect 18962 29902 18966 30198
rect 18342 29898 18966 29902
rect 19002 30198 19306 30202
rect 19002 29902 19006 30198
rect 19006 29902 19302 30198
rect 19302 29902 19306 30198
rect 19002 29898 19306 29902
rect 19342 30198 19966 30202
rect 19342 29902 19346 30198
rect 19346 29902 19962 30198
rect 19962 29902 19966 30198
rect 19342 29898 19966 29902
rect 20002 30198 20306 30202
rect 20002 29902 20006 30198
rect 20006 29902 20302 30198
rect 20302 29902 20306 30198
rect 20002 29898 20306 29902
rect 20342 30198 20966 30202
rect 20342 29902 20346 30198
rect 20346 29902 20962 30198
rect 20962 29902 20966 30198
rect 20342 29898 20966 29902
rect 21002 30198 21306 30202
rect 21002 29902 21006 30198
rect 21006 29902 21302 30198
rect 21302 29902 21306 30198
rect 21002 29898 21306 29902
rect 21342 30198 21966 30202
rect 21342 29902 21346 30198
rect 21346 29902 21962 30198
rect 21962 29902 21966 30198
rect 21342 29898 21966 29902
rect 22002 30198 22306 30202
rect 22002 29902 22006 30198
rect 22006 29902 22302 30198
rect 22302 29902 22306 30198
rect 22002 29898 22306 29902
rect 22342 30198 22966 30202
rect 22342 29902 22346 30198
rect 22346 29902 22962 30198
rect 22962 29902 22966 30198
rect 22342 29898 22966 29902
rect 23002 30198 23306 30202
rect 23002 29902 23006 30198
rect 23006 29902 23302 30198
rect 23302 29902 23306 30198
rect 23002 29898 23306 29902
rect 23342 30198 23966 30202
rect 23342 29902 23346 30198
rect 23346 29902 23962 30198
rect 23962 29902 23966 30198
rect 23342 29898 23966 29902
rect 24002 30198 24306 30202
rect 24002 29902 24006 30198
rect 24006 29902 24302 30198
rect 24302 29902 24306 30198
rect 24002 29898 24306 29902
rect 24342 30198 24966 30202
rect 24342 29902 24346 30198
rect 24346 29902 24962 30198
rect 24962 29902 24966 30198
rect 24342 29898 24966 29902
rect 25002 30198 25306 30202
rect 25002 29902 25006 30198
rect 25006 29902 25302 30198
rect 25302 29902 25306 30198
rect 25002 29898 25306 29902
rect 25342 30198 25966 30202
rect 25342 29902 25346 30198
rect 25346 29902 25962 30198
rect 25962 29902 25966 30198
rect 25342 29898 25966 29902
rect 26002 30198 26306 30202
rect 26002 29902 26006 30198
rect 26006 29902 26302 30198
rect 26302 29902 26306 30198
rect 26002 29898 26306 29902
rect 26342 30198 26966 30202
rect 26342 29902 26346 30198
rect 26346 29902 26962 30198
rect 26962 29902 26966 30198
rect 26342 29898 26966 29902
rect 27002 30198 27306 30202
rect 27002 29902 27006 30198
rect 27006 29902 27302 30198
rect 27302 29902 27306 30198
rect 27002 29898 27306 29902
rect 27342 30198 27966 30202
rect 27342 29902 27346 30198
rect 27346 29902 27962 30198
rect 27962 29902 27966 30198
rect 27342 29898 27966 29902
rect 28002 30198 28306 30202
rect 28002 29902 28006 30198
rect 28006 29902 28302 30198
rect 28302 29902 28306 30198
rect 28002 29898 28306 29902
rect 28342 30198 28966 30202
rect 28342 29902 28346 30198
rect 28346 29902 28962 30198
rect 28962 29902 28966 30198
rect 28342 29898 28966 29902
rect 29002 30198 29306 30202
rect 29002 29902 29006 30198
rect 29006 29902 29302 30198
rect 29302 29902 29306 30198
rect 29002 29898 29306 29902
rect 29342 30198 29966 30202
rect 29342 29902 29346 30198
rect 29346 29902 29962 30198
rect 29962 29902 29966 30198
rect 29342 29898 29966 29902
rect 30002 30198 30306 30202
rect 30002 29902 30006 30198
rect 30006 29902 30302 30198
rect 30302 29902 30306 30198
rect 30002 29898 30306 29902
rect 30342 30198 30966 30202
rect 30342 29902 30346 30198
rect 30346 29902 30962 30198
rect 30962 29902 30966 30198
rect 30342 29898 30966 29902
rect 31002 30198 31306 30202
rect 31002 29902 31006 30198
rect 31006 29902 31302 30198
rect 31302 29902 31306 30198
rect 31002 29898 31306 29902
rect 31342 30198 31966 30202
rect 31342 29902 31346 30198
rect 31346 29902 31962 30198
rect 31962 29902 31966 30198
rect 31342 29898 31966 29902
rect 32002 30198 32306 30202
rect 32002 29902 32006 30198
rect 32006 29902 32302 30198
rect 32302 29902 32306 30198
rect 32002 29898 32306 29902
rect 32342 30198 32966 30202
rect 32342 29902 32346 30198
rect 32346 29902 32962 30198
rect 32962 29902 32966 30198
rect 32342 29898 32966 29902
rect 33002 30198 33306 30202
rect 33002 29902 33006 30198
rect 33006 29902 33302 30198
rect 33302 29902 33306 30198
rect 33002 29898 33306 29902
rect 33342 30198 33966 30202
rect 33342 29902 33346 30198
rect 33346 29902 33962 30198
rect 33962 29902 33966 30198
rect 33342 29898 33966 29902
rect 34002 30198 34306 30202
rect 34002 29902 34006 30198
rect 34006 29902 34302 30198
rect 34302 29902 34306 30198
rect 34002 29898 34306 29902
rect 34342 30198 34646 30202
rect 34342 29902 34346 30198
rect 34346 29902 34642 30198
rect 34642 29902 34646 30198
rect 34342 29898 34646 29902
rect -74477 29858 -74173 29862
rect -74477 29242 -74473 29858
rect -74473 29242 -74177 29858
rect -74177 29242 -74173 29858
rect -74477 29238 -74173 29242
rect -73477 29858 -73173 29862
rect -73477 29242 -73473 29858
rect -73473 29242 -73177 29858
rect -73177 29242 -73173 29858
rect -73477 29238 -73173 29242
rect -72477 29858 -72173 29862
rect -72477 29242 -72473 29858
rect -72473 29242 -72177 29858
rect -72177 29242 -72173 29858
rect -72477 29238 -72173 29242
rect -71477 29858 -71173 29862
rect -71477 29242 -71473 29858
rect -71473 29242 -71177 29858
rect -71177 29242 -71173 29858
rect -71477 29238 -71173 29242
rect -70477 29858 -70173 29862
rect -70477 29242 -70473 29858
rect -70473 29242 -70177 29858
rect -70177 29242 -70173 29858
rect -70477 29238 -70173 29242
rect -69477 29858 -69173 29862
rect -69477 29242 -69473 29858
rect -69473 29242 -69177 29858
rect -69177 29242 -69173 29858
rect -69477 29238 -69173 29242
rect -68477 29858 -68173 29862
rect -68477 29242 -68473 29858
rect -68473 29242 -68177 29858
rect -68177 29242 -68173 29858
rect -68477 29238 -68173 29242
rect -67477 29858 -67173 29862
rect -67477 29242 -67473 29858
rect -67473 29242 -67177 29858
rect -67177 29242 -67173 29858
rect -67477 29238 -67173 29242
rect -66477 29858 -66173 29862
rect -66477 29242 -66473 29858
rect -66473 29242 -66177 29858
rect -66177 29242 -66173 29858
rect -66477 29238 -66173 29242
rect -65477 29858 -65173 29862
rect -65477 29242 -65473 29858
rect -65473 29242 -65177 29858
rect -65177 29242 -65173 29858
rect -65477 29238 -65173 29242
rect -64477 29858 -64173 29862
rect -64477 29242 -64473 29858
rect -64473 29242 -64177 29858
rect -64177 29242 -64173 29858
rect -64477 29238 -64173 29242
rect -63477 29858 -63173 29862
rect -63477 29242 -63473 29858
rect -63473 29242 -63177 29858
rect -63177 29242 -63173 29858
rect -63477 29238 -63173 29242
rect -62477 29858 -62173 29862
rect -62477 29242 -62473 29858
rect -62473 29242 -62177 29858
rect -62177 29242 -62173 29858
rect -62477 29238 -62173 29242
rect -61477 29858 -61173 29862
rect -61477 29242 -61473 29858
rect -61473 29242 -61177 29858
rect -61177 29242 -61173 29858
rect -61477 29238 -61173 29242
rect -60477 29858 -60173 29862
rect -60477 29242 -60473 29858
rect -60473 29242 -60177 29858
rect -60177 29242 -60173 29858
rect -60477 29238 -60173 29242
rect -59477 29858 -59173 29862
rect -59477 29242 -59473 29858
rect -59473 29242 -59177 29858
rect -59177 29242 -59173 29858
rect -59477 29238 -59173 29242
rect 10002 29858 10306 29862
rect 10002 29242 10006 29858
rect 10006 29242 10302 29858
rect 10302 29242 10306 29858
rect 10002 29238 10306 29242
rect 11002 29858 11306 29862
rect 11002 29242 11006 29858
rect 11006 29242 11302 29858
rect 11302 29242 11306 29858
rect 11002 29238 11306 29242
rect 12002 29858 12306 29862
rect 12002 29242 12006 29858
rect 12006 29242 12302 29858
rect 12302 29242 12306 29858
rect 12002 29238 12306 29242
rect 13002 29858 13306 29862
rect 13002 29242 13006 29858
rect 13006 29242 13302 29858
rect 13302 29242 13306 29858
rect 13002 29238 13306 29242
rect 14002 29858 14306 29862
rect 14002 29242 14006 29858
rect 14006 29242 14302 29858
rect 14302 29242 14306 29858
rect 14002 29238 14306 29242
rect 15002 29858 15306 29862
rect 15002 29242 15006 29858
rect 15006 29242 15302 29858
rect 15302 29242 15306 29858
rect 15002 29238 15306 29242
rect 16002 29858 16306 29862
rect 16002 29242 16006 29858
rect 16006 29242 16302 29858
rect 16302 29242 16306 29858
rect 16002 29238 16306 29242
rect 17002 29858 17306 29862
rect 17002 29242 17006 29858
rect 17006 29242 17302 29858
rect 17302 29242 17306 29858
rect 17002 29238 17306 29242
rect 18002 29858 18306 29862
rect 18002 29242 18006 29858
rect 18006 29242 18302 29858
rect 18302 29242 18306 29858
rect 18002 29238 18306 29242
rect 19002 29858 19306 29862
rect 19002 29242 19006 29858
rect 19006 29242 19302 29858
rect 19302 29242 19306 29858
rect 19002 29238 19306 29242
rect 20002 29858 20306 29862
rect 20002 29242 20006 29858
rect 20006 29242 20302 29858
rect 20302 29242 20306 29858
rect 20002 29238 20306 29242
rect 21002 29858 21306 29862
rect 21002 29242 21006 29858
rect 21006 29242 21302 29858
rect 21302 29242 21306 29858
rect 21002 29238 21306 29242
rect 22002 29858 22306 29862
rect 22002 29242 22006 29858
rect 22006 29242 22302 29858
rect 22302 29242 22306 29858
rect 22002 29238 22306 29242
rect 23002 29858 23306 29862
rect 23002 29242 23006 29858
rect 23006 29242 23302 29858
rect 23302 29242 23306 29858
rect 23002 29238 23306 29242
rect 24002 29858 24306 29862
rect 24002 29242 24006 29858
rect 24006 29242 24302 29858
rect 24302 29242 24306 29858
rect 24002 29238 24306 29242
rect 25002 29858 25306 29862
rect 25002 29242 25006 29858
rect 25006 29242 25302 29858
rect 25302 29242 25306 29858
rect 25002 29238 25306 29242
rect 26002 29858 26306 29862
rect 26002 29242 26006 29858
rect 26006 29242 26302 29858
rect 26302 29242 26306 29858
rect 26002 29238 26306 29242
rect 27002 29858 27306 29862
rect 27002 29242 27006 29858
rect 27006 29242 27302 29858
rect 27302 29242 27306 29858
rect 27002 29238 27306 29242
rect 28002 29858 28306 29862
rect 28002 29242 28006 29858
rect 28006 29242 28302 29858
rect 28302 29242 28306 29858
rect 28002 29238 28306 29242
rect 29002 29858 29306 29862
rect 29002 29242 29006 29858
rect 29006 29242 29302 29858
rect 29302 29242 29306 29858
rect 29002 29238 29306 29242
rect 30002 29858 30306 29862
rect 30002 29242 30006 29858
rect 30006 29242 30302 29858
rect 30302 29242 30306 29858
rect 30002 29238 30306 29242
rect 31002 29858 31306 29862
rect 31002 29242 31006 29858
rect 31006 29242 31302 29858
rect 31302 29242 31306 29858
rect 31002 29238 31306 29242
rect 32002 29858 32306 29862
rect 32002 29242 32006 29858
rect 32006 29242 32302 29858
rect 32302 29242 32306 29858
rect 32002 29238 32306 29242
rect 33002 29858 33306 29862
rect 33002 29242 33006 29858
rect 33006 29242 33302 29858
rect 33302 29242 33306 29858
rect 33002 29238 33306 29242
rect 34002 29858 34306 29862
rect 34002 29242 34006 29858
rect 34006 29242 34302 29858
rect 34302 29242 34306 29858
rect 34002 29238 34306 29242
rect -74817 29198 -74513 29202
rect -74817 28902 -74813 29198
rect -74813 28902 -74517 29198
rect -74517 28902 -74513 29198
rect -74817 28898 -74513 28902
rect -74477 29198 -74173 29202
rect -74477 28902 -74473 29198
rect -74473 28902 -74177 29198
rect -74177 28902 -74173 29198
rect -74477 28898 -74173 28902
rect -74137 29198 -73513 29202
rect -74137 28902 -74133 29198
rect -74133 28902 -73517 29198
rect -73517 28902 -73513 29198
rect -74137 28898 -73513 28902
rect -73477 29198 -73173 29202
rect -73477 28902 -73473 29198
rect -73473 28902 -73177 29198
rect -73177 28902 -73173 29198
rect -73477 28898 -73173 28902
rect -73137 29198 -72513 29202
rect -73137 28902 -73133 29198
rect -73133 28902 -72517 29198
rect -72517 28902 -72513 29198
rect -73137 28898 -72513 28902
rect -72477 29198 -72173 29202
rect -72477 28902 -72473 29198
rect -72473 28902 -72177 29198
rect -72177 28902 -72173 29198
rect -72477 28898 -72173 28902
rect -72137 29198 -71513 29202
rect -72137 28902 -72133 29198
rect -72133 28902 -71517 29198
rect -71517 28902 -71513 29198
rect -72137 28898 -71513 28902
rect -71477 29198 -71173 29202
rect -71477 28902 -71473 29198
rect -71473 28902 -71177 29198
rect -71177 28902 -71173 29198
rect -71477 28898 -71173 28902
rect -71137 29198 -70513 29202
rect -71137 28902 -71133 29198
rect -71133 28902 -70517 29198
rect -70517 28902 -70513 29198
rect -71137 28898 -70513 28902
rect -70477 29198 -70173 29202
rect -70477 28902 -70473 29198
rect -70473 28902 -70177 29198
rect -70177 28902 -70173 29198
rect -70477 28898 -70173 28902
rect -70137 29198 -69513 29202
rect -70137 28902 -70133 29198
rect -70133 28902 -69517 29198
rect -69517 28902 -69513 29198
rect -70137 28898 -69513 28902
rect -69477 29198 -69173 29202
rect -69477 28902 -69473 29198
rect -69473 28902 -69177 29198
rect -69177 28902 -69173 29198
rect -69477 28898 -69173 28902
rect -69137 29198 -68513 29202
rect -69137 28902 -69133 29198
rect -69133 28902 -68517 29198
rect -68517 28902 -68513 29198
rect -69137 28898 -68513 28902
rect -68477 29198 -68173 29202
rect -68477 28902 -68473 29198
rect -68473 28902 -68177 29198
rect -68177 28902 -68173 29198
rect -68477 28898 -68173 28902
rect -68137 29198 -67513 29202
rect -68137 28902 -68133 29198
rect -68133 28902 -67517 29198
rect -67517 28902 -67513 29198
rect -68137 28898 -67513 28902
rect -67477 29198 -67173 29202
rect -67477 28902 -67473 29198
rect -67473 28902 -67177 29198
rect -67177 28902 -67173 29198
rect -67477 28898 -67173 28902
rect -67137 29198 -66513 29202
rect -67137 28902 -67133 29198
rect -67133 28902 -66517 29198
rect -66517 28902 -66513 29198
rect -67137 28898 -66513 28902
rect -66477 29198 -66173 29202
rect -66477 28902 -66473 29198
rect -66473 28902 -66177 29198
rect -66177 28902 -66173 29198
rect -66477 28898 -66173 28902
rect -66137 29198 -65513 29202
rect -66137 28902 -66133 29198
rect -66133 28902 -65517 29198
rect -65517 28902 -65513 29198
rect -66137 28898 -65513 28902
rect -65477 29198 -65173 29202
rect -65477 28902 -65473 29198
rect -65473 28902 -65177 29198
rect -65177 28902 -65173 29198
rect -65477 28898 -65173 28902
rect -65137 29198 -64513 29202
rect -65137 28902 -65133 29198
rect -65133 28902 -64517 29198
rect -64517 28902 -64513 29198
rect -65137 28898 -64513 28902
rect -64477 29198 -64173 29202
rect -64477 28902 -64473 29198
rect -64473 28902 -64177 29198
rect -64177 28902 -64173 29198
rect -64477 28898 -64173 28902
rect -64137 29198 -63513 29202
rect -64137 28902 -64133 29198
rect -64133 28902 -63517 29198
rect -63517 28902 -63513 29198
rect -64137 28898 -63513 28902
rect -63477 29198 -63173 29202
rect -63477 28902 -63473 29198
rect -63473 28902 -63177 29198
rect -63177 28902 -63173 29198
rect -63477 28898 -63173 28902
rect -63137 29198 -62513 29202
rect -63137 28902 -63133 29198
rect -63133 28902 -62517 29198
rect -62517 28902 -62513 29198
rect -63137 28898 -62513 28902
rect -62477 29198 -62173 29202
rect -62477 28902 -62473 29198
rect -62473 28902 -62177 29198
rect -62177 28902 -62173 29198
rect -62477 28898 -62173 28902
rect -62137 29198 -61513 29202
rect -62137 28902 -62133 29198
rect -62133 28902 -61517 29198
rect -61517 28902 -61513 29198
rect -62137 28898 -61513 28902
rect -61477 29198 -61173 29202
rect -61477 28902 -61473 29198
rect -61473 28902 -61177 29198
rect -61177 28902 -61173 29198
rect -61477 28898 -61173 28902
rect -61137 29198 -60513 29202
rect -61137 28902 -61133 29198
rect -61133 28902 -60517 29198
rect -60517 28902 -60513 29198
rect -61137 28898 -60513 28902
rect -60477 29198 -60173 29202
rect -60477 28902 -60473 29198
rect -60473 28902 -60177 29198
rect -60177 28902 -60173 29198
rect -60477 28898 -60173 28902
rect -60137 29198 -59513 29202
rect -60137 28902 -60133 29198
rect -60133 28902 -59517 29198
rect -59517 28902 -59513 29198
rect -60137 28898 -59513 28902
rect -59477 29198 -59173 29202
rect -59477 28902 -59473 29198
rect -59473 28902 -59177 29198
rect -59177 28902 -59173 29198
rect -59477 28898 -59173 28902
rect -59137 29198 -58833 29202
rect -59137 28902 -59133 29198
rect -59133 28902 -58837 29198
rect -58837 28902 -58833 29198
rect -59137 28898 -58833 28902
rect 9662 29198 9966 29202
rect 9662 28902 9666 29198
rect 9666 28902 9962 29198
rect 9962 28902 9966 29198
rect 9662 28898 9966 28902
rect 10002 29198 10306 29202
rect 10002 28902 10006 29198
rect 10006 28902 10302 29198
rect 10302 28902 10306 29198
rect 10002 28898 10306 28902
rect 10342 29198 10966 29202
rect 10342 28902 10346 29198
rect 10346 28902 10962 29198
rect 10962 28902 10966 29198
rect 10342 28898 10966 28902
rect 11002 29198 11306 29202
rect 11002 28902 11006 29198
rect 11006 28902 11302 29198
rect 11302 28902 11306 29198
rect 11002 28898 11306 28902
rect 11342 29198 11966 29202
rect 11342 28902 11346 29198
rect 11346 28902 11962 29198
rect 11962 28902 11966 29198
rect 11342 28898 11966 28902
rect 12002 29198 12306 29202
rect 12002 28902 12006 29198
rect 12006 28902 12302 29198
rect 12302 28902 12306 29198
rect 12002 28898 12306 28902
rect 12342 29198 12966 29202
rect 12342 28902 12346 29198
rect 12346 28902 12962 29198
rect 12962 28902 12966 29198
rect 12342 28898 12966 28902
rect 13002 29198 13306 29202
rect 13002 28902 13006 29198
rect 13006 28902 13302 29198
rect 13302 28902 13306 29198
rect 13002 28898 13306 28902
rect 13342 29198 13966 29202
rect 13342 28902 13346 29198
rect 13346 28902 13962 29198
rect 13962 28902 13966 29198
rect 13342 28898 13966 28902
rect 14002 29198 14306 29202
rect 14002 28902 14006 29198
rect 14006 28902 14302 29198
rect 14302 28902 14306 29198
rect 14002 28898 14306 28902
rect 14342 29198 14966 29202
rect 14342 28902 14346 29198
rect 14346 28902 14962 29198
rect 14962 28902 14966 29198
rect 14342 28898 14966 28902
rect 15002 29198 15306 29202
rect 15002 28902 15006 29198
rect 15006 28902 15302 29198
rect 15302 28902 15306 29198
rect 15002 28898 15306 28902
rect 15342 29198 15966 29202
rect 15342 28902 15346 29198
rect 15346 28902 15962 29198
rect 15962 28902 15966 29198
rect 15342 28898 15966 28902
rect 16002 29198 16306 29202
rect 16002 28902 16006 29198
rect 16006 28902 16302 29198
rect 16302 28902 16306 29198
rect 16002 28898 16306 28902
rect 16342 29198 16966 29202
rect 16342 28902 16346 29198
rect 16346 28902 16962 29198
rect 16962 28902 16966 29198
rect 16342 28898 16966 28902
rect 17002 29198 17306 29202
rect 17002 28902 17006 29198
rect 17006 28902 17302 29198
rect 17302 28902 17306 29198
rect 17002 28898 17306 28902
rect 17342 29198 17966 29202
rect 17342 28902 17346 29198
rect 17346 28902 17962 29198
rect 17962 28902 17966 29198
rect 17342 28898 17966 28902
rect 18002 29198 18306 29202
rect 18002 28902 18006 29198
rect 18006 28902 18302 29198
rect 18302 28902 18306 29198
rect 18002 28898 18306 28902
rect 18342 29198 18966 29202
rect 18342 28902 18346 29198
rect 18346 28902 18962 29198
rect 18962 28902 18966 29198
rect 18342 28898 18966 28902
rect 19002 29198 19306 29202
rect 19002 28902 19006 29198
rect 19006 28902 19302 29198
rect 19302 28902 19306 29198
rect 19002 28898 19306 28902
rect 19342 29198 19966 29202
rect 19342 28902 19346 29198
rect 19346 28902 19962 29198
rect 19962 28902 19966 29198
rect 19342 28898 19966 28902
rect 20002 29198 20306 29202
rect 20002 28902 20006 29198
rect 20006 28902 20302 29198
rect 20302 28902 20306 29198
rect 20002 28898 20306 28902
rect 20342 29198 20966 29202
rect 20342 28902 20346 29198
rect 20346 28902 20962 29198
rect 20962 28902 20966 29198
rect 20342 28898 20966 28902
rect 21002 29198 21306 29202
rect 21002 28902 21006 29198
rect 21006 28902 21302 29198
rect 21302 28902 21306 29198
rect 21002 28898 21306 28902
rect 21342 29198 21966 29202
rect 21342 28902 21346 29198
rect 21346 28902 21962 29198
rect 21962 28902 21966 29198
rect 21342 28898 21966 28902
rect 22002 29198 22306 29202
rect 22002 28902 22006 29198
rect 22006 28902 22302 29198
rect 22302 28902 22306 29198
rect 22002 28898 22306 28902
rect 22342 29198 22966 29202
rect 22342 28902 22346 29198
rect 22346 28902 22962 29198
rect 22962 28902 22966 29198
rect 22342 28898 22966 28902
rect 23002 29198 23306 29202
rect 23002 28902 23006 29198
rect 23006 28902 23302 29198
rect 23302 28902 23306 29198
rect 23002 28898 23306 28902
rect 23342 29198 23966 29202
rect 23342 28902 23346 29198
rect 23346 28902 23962 29198
rect 23962 28902 23966 29198
rect 23342 28898 23966 28902
rect 24002 29198 24306 29202
rect 24002 28902 24006 29198
rect 24006 28902 24302 29198
rect 24302 28902 24306 29198
rect 24002 28898 24306 28902
rect 24342 29198 24966 29202
rect 24342 28902 24346 29198
rect 24346 28902 24962 29198
rect 24962 28902 24966 29198
rect 24342 28898 24966 28902
rect 25002 29198 25306 29202
rect 25002 28902 25006 29198
rect 25006 28902 25302 29198
rect 25302 28902 25306 29198
rect 25002 28898 25306 28902
rect 25342 29198 25966 29202
rect 25342 28902 25346 29198
rect 25346 28902 25962 29198
rect 25962 28902 25966 29198
rect 25342 28898 25966 28902
rect 26002 29198 26306 29202
rect 26002 28902 26006 29198
rect 26006 28902 26302 29198
rect 26302 28902 26306 29198
rect 26002 28898 26306 28902
rect 26342 29198 26966 29202
rect 26342 28902 26346 29198
rect 26346 28902 26962 29198
rect 26962 28902 26966 29198
rect 26342 28898 26966 28902
rect 27002 29198 27306 29202
rect 27002 28902 27006 29198
rect 27006 28902 27302 29198
rect 27302 28902 27306 29198
rect 27002 28898 27306 28902
rect 27342 29198 27966 29202
rect 27342 28902 27346 29198
rect 27346 28902 27962 29198
rect 27962 28902 27966 29198
rect 27342 28898 27966 28902
rect 28002 29198 28306 29202
rect 28002 28902 28006 29198
rect 28006 28902 28302 29198
rect 28302 28902 28306 29198
rect 28002 28898 28306 28902
rect 28342 29198 28966 29202
rect 28342 28902 28346 29198
rect 28346 28902 28962 29198
rect 28962 28902 28966 29198
rect 28342 28898 28966 28902
rect 29002 29198 29306 29202
rect 29002 28902 29006 29198
rect 29006 28902 29302 29198
rect 29302 28902 29306 29198
rect 29002 28898 29306 28902
rect 29342 29198 29966 29202
rect 29342 28902 29346 29198
rect 29346 28902 29962 29198
rect 29962 28902 29966 29198
rect 29342 28898 29966 28902
rect 30002 29198 30306 29202
rect 30002 28902 30006 29198
rect 30006 28902 30302 29198
rect 30302 28902 30306 29198
rect 30002 28898 30306 28902
rect 30342 29198 30966 29202
rect 30342 28902 30346 29198
rect 30346 28902 30962 29198
rect 30962 28902 30966 29198
rect 30342 28898 30966 28902
rect 31002 29198 31306 29202
rect 31002 28902 31006 29198
rect 31006 28902 31302 29198
rect 31302 28902 31306 29198
rect 31002 28898 31306 28902
rect 31342 29198 31966 29202
rect 31342 28902 31346 29198
rect 31346 28902 31962 29198
rect 31962 28902 31966 29198
rect 31342 28898 31966 28902
rect 32002 29198 32306 29202
rect 32002 28902 32006 29198
rect 32006 28902 32302 29198
rect 32302 28902 32306 29198
rect 32002 28898 32306 28902
rect 32342 29198 32966 29202
rect 32342 28902 32346 29198
rect 32346 28902 32962 29198
rect 32962 28902 32966 29198
rect 32342 28898 32966 28902
rect 33002 29198 33306 29202
rect 33002 28902 33006 29198
rect 33006 28902 33302 29198
rect 33302 28902 33306 29198
rect 33002 28898 33306 28902
rect 33342 29198 33966 29202
rect 33342 28902 33346 29198
rect 33346 28902 33962 29198
rect 33962 28902 33966 29198
rect 33342 28898 33966 28902
rect 34002 29198 34306 29202
rect 34002 28902 34006 29198
rect 34006 28902 34302 29198
rect 34302 28902 34306 29198
rect 34002 28898 34306 28902
rect 34342 29198 34646 29202
rect 34342 28902 34346 29198
rect 34346 28902 34642 29198
rect 34642 28902 34646 29198
rect 34342 28898 34646 28902
rect -74477 28858 -74173 28862
rect -74477 28562 -74473 28858
rect -74473 28562 -74177 28858
rect -74177 28562 -74173 28858
rect -74477 28558 -74173 28562
rect -73477 28858 -73173 28862
rect -73477 28562 -73473 28858
rect -73473 28562 -73177 28858
rect -73177 28562 -73173 28858
rect -73477 28558 -73173 28562
rect -72477 28858 -72173 28862
rect -72477 28562 -72473 28858
rect -72473 28562 -72177 28858
rect -72177 28562 -72173 28858
rect -72477 28558 -72173 28562
rect -71477 28858 -71173 28862
rect -71477 28562 -71473 28858
rect -71473 28562 -71177 28858
rect -71177 28562 -71173 28858
rect -71477 28558 -71173 28562
rect -70477 28858 -70173 28862
rect -70477 28562 -70473 28858
rect -70473 28562 -70177 28858
rect -70177 28562 -70173 28858
rect -70477 28558 -70173 28562
rect -69477 28858 -69173 28862
rect -69477 28562 -69473 28858
rect -69473 28562 -69177 28858
rect -69177 28562 -69173 28858
rect -69477 28558 -69173 28562
rect -68477 28858 -68173 28862
rect -68477 28562 -68473 28858
rect -68473 28562 -68177 28858
rect -68177 28562 -68173 28858
rect -68477 28558 -68173 28562
rect -67477 28858 -67173 28862
rect -67477 28562 -67473 28858
rect -67473 28562 -67177 28858
rect -67177 28562 -67173 28858
rect -67477 28558 -67173 28562
rect -66477 28858 -66173 28862
rect -66477 28562 -66473 28858
rect -66473 28562 -66177 28858
rect -66177 28562 -66173 28858
rect -66477 28558 -66173 28562
rect -65477 28858 -65173 28862
rect -65477 28562 -65473 28858
rect -65473 28562 -65177 28858
rect -65177 28562 -65173 28858
rect -65477 28558 -65173 28562
rect -64477 28858 -64173 28862
rect -64477 28562 -64473 28858
rect -64473 28562 -64177 28858
rect -64177 28562 -64173 28858
rect -64477 28558 -64173 28562
rect -63477 28858 -63173 28862
rect -63477 28562 -63473 28858
rect -63473 28562 -63177 28858
rect -63177 28562 -63173 28858
rect -63477 28558 -63173 28562
rect -62477 28858 -62173 28862
rect -62477 28562 -62473 28858
rect -62473 28562 -62177 28858
rect -62177 28562 -62173 28858
rect -62477 28558 -62173 28562
rect -61477 28858 -61173 28862
rect -61477 28562 -61473 28858
rect -61473 28562 -61177 28858
rect -61177 28562 -61173 28858
rect -61477 28558 -61173 28562
rect -60477 28858 -60173 28862
rect -60477 28562 -60473 28858
rect -60473 28562 -60177 28858
rect -60177 28562 -60173 28858
rect -60477 28558 -60173 28562
rect -59477 28858 -59173 28862
rect -59477 28562 -59473 28858
rect -59473 28562 -59177 28858
rect -59177 28562 -59173 28858
rect -59477 28558 -59173 28562
rect 10002 28858 10306 28862
rect 10002 28562 10006 28858
rect 10006 28562 10302 28858
rect 10302 28562 10306 28858
rect 10002 28558 10306 28562
rect 11002 28858 11306 28862
rect 11002 28562 11006 28858
rect 11006 28562 11302 28858
rect 11302 28562 11306 28858
rect 11002 28558 11306 28562
rect 12002 28858 12306 28862
rect 12002 28562 12006 28858
rect 12006 28562 12302 28858
rect 12302 28562 12306 28858
rect 12002 28558 12306 28562
rect 13002 28858 13306 28862
rect 13002 28562 13006 28858
rect 13006 28562 13302 28858
rect 13302 28562 13306 28858
rect 13002 28558 13306 28562
rect 14002 28858 14306 28862
rect 14002 28562 14006 28858
rect 14006 28562 14302 28858
rect 14302 28562 14306 28858
rect 14002 28558 14306 28562
rect 15002 28858 15306 28862
rect 15002 28562 15006 28858
rect 15006 28562 15302 28858
rect 15302 28562 15306 28858
rect 15002 28558 15306 28562
rect 16002 28858 16306 28862
rect 16002 28562 16006 28858
rect 16006 28562 16302 28858
rect 16302 28562 16306 28858
rect 16002 28558 16306 28562
rect 17002 28858 17306 28862
rect 17002 28562 17006 28858
rect 17006 28562 17302 28858
rect 17302 28562 17306 28858
rect 17002 28558 17306 28562
rect 18002 28858 18306 28862
rect 18002 28562 18006 28858
rect 18006 28562 18302 28858
rect 18302 28562 18306 28858
rect 18002 28558 18306 28562
rect 19002 28858 19306 28862
rect 19002 28562 19006 28858
rect 19006 28562 19302 28858
rect 19302 28562 19306 28858
rect 19002 28558 19306 28562
rect 20002 28858 20306 28862
rect 20002 28562 20006 28858
rect 20006 28562 20302 28858
rect 20302 28562 20306 28858
rect 20002 28558 20306 28562
rect 21002 28858 21306 28862
rect 21002 28562 21006 28858
rect 21006 28562 21302 28858
rect 21302 28562 21306 28858
rect 21002 28558 21306 28562
rect 22002 28858 22306 28862
rect 22002 28562 22006 28858
rect 22006 28562 22302 28858
rect 22302 28562 22306 28858
rect 22002 28558 22306 28562
rect 23002 28858 23306 28862
rect 23002 28562 23006 28858
rect 23006 28562 23302 28858
rect 23302 28562 23306 28858
rect 23002 28558 23306 28562
rect 24002 28858 24306 28862
rect 24002 28562 24006 28858
rect 24006 28562 24302 28858
rect 24302 28562 24306 28858
rect 24002 28558 24306 28562
rect 25002 28858 25306 28862
rect 25002 28562 25006 28858
rect 25006 28562 25302 28858
rect 25302 28562 25306 28858
rect 25002 28558 25306 28562
rect 26002 28858 26306 28862
rect 26002 28562 26006 28858
rect 26006 28562 26302 28858
rect 26302 28562 26306 28858
rect 26002 28558 26306 28562
rect 27002 28858 27306 28862
rect 27002 28562 27006 28858
rect 27006 28562 27302 28858
rect 27302 28562 27306 28858
rect 27002 28558 27306 28562
rect 28002 28858 28306 28862
rect 28002 28562 28006 28858
rect 28006 28562 28302 28858
rect 28302 28562 28306 28858
rect 28002 28558 28306 28562
rect 29002 28858 29306 28862
rect 29002 28562 29006 28858
rect 29006 28562 29302 28858
rect 29302 28562 29306 28858
rect 29002 28558 29306 28562
rect 30002 28858 30306 28862
rect 30002 28562 30006 28858
rect 30006 28562 30302 28858
rect 30302 28562 30306 28858
rect 30002 28558 30306 28562
rect 31002 28858 31306 28862
rect 31002 28562 31006 28858
rect 31006 28562 31302 28858
rect 31302 28562 31306 28858
rect 31002 28558 31306 28562
rect 32002 28858 32306 28862
rect 32002 28562 32006 28858
rect 32006 28562 32302 28858
rect 32302 28562 32306 28858
rect 32002 28558 32306 28562
rect 33002 28858 33306 28862
rect 33002 28562 33006 28858
rect 33006 28562 33302 28858
rect 33302 28562 33306 28858
rect 33002 28558 33306 28562
rect 34002 28858 34306 28862
rect 34002 28562 34006 28858
rect 34006 28562 34302 28858
rect 34302 28562 34306 28858
rect 34002 28558 34306 28562
rect -72782 25943 -60878 25947
rect -72782 16047 -72778 25943
rect -72778 16047 -60882 25943
rect -60882 16047 -60878 25943
rect -72782 16043 -60878 16047
rect 20318 25948 32222 25952
rect 20318 16052 20322 25948
rect 20322 16052 32218 25948
rect 32218 16052 32222 25948
rect 20318 16048 32222 16052
rect -21210 15118 -19306 15122
rect -21210 13862 -21206 15118
rect -21206 13862 -19310 15118
rect -19310 13862 -19306 15118
rect -21210 13858 -19306 13862
rect -42382 13798 -40718 13802
rect -42382 7902 -42378 13798
rect -42378 7902 -40722 13798
rect -40722 7902 -40718 13798
rect -42382 7898 -40718 7902
rect 168 13798 1832 13802
rect 168 7902 172 13798
rect 172 7902 1828 13798
rect 1828 7902 1832 13798
rect 168 7898 1832 7902
rect -42382 2308 -40718 2312
rect -42382 -2308 -42378 2308
rect -42378 -2308 -40722 2308
rect -40722 -2308 -40718 2308
rect -42382 -2312 -40718 -2308
rect 168 2308 1832 2312
rect 168 -2308 172 2308
rect 172 -2308 1828 2308
rect 1828 -2308 1832 2308
rect 168 -2312 1832 -2308
rect -42382 -7902 -40718 -7898
rect -42382 -13798 -42378 -7902
rect -42378 -13798 -40722 -7902
rect -40722 -13798 -40718 -7902
rect -42382 -13802 -40718 -13798
rect 168 -7902 1832 -7898
rect 168 -13798 172 -7902
rect 172 -13798 1828 -7902
rect 1828 -13798 1832 -7902
rect 168 -13802 1832 -13798
rect -72782 -16052 -60878 -16048
rect -72782 -25948 -72778 -16052
rect -72778 -25948 -60882 -16052
rect -60882 -25948 -60878 -16052
rect -72782 -25952 -60878 -25948
rect 20318 -16052 32222 -16048
rect 20318 -25948 20322 -16052
rect 20322 -25948 32218 -16052
rect 32218 -25948 32222 -16052
rect 20318 -25952 32222 -25948
rect -74477 -28562 -74173 -28558
rect -74477 -28858 -74473 -28562
rect -74473 -28858 -74177 -28562
rect -74177 -28858 -74173 -28562
rect -74477 -28862 -74173 -28858
rect -73477 -28562 -73173 -28558
rect -73477 -28858 -73473 -28562
rect -73473 -28858 -73177 -28562
rect -73177 -28858 -73173 -28562
rect -73477 -28862 -73173 -28858
rect -72477 -28562 -72173 -28558
rect -72477 -28858 -72473 -28562
rect -72473 -28858 -72177 -28562
rect -72177 -28858 -72173 -28562
rect -72477 -28862 -72173 -28858
rect -71477 -28562 -71173 -28558
rect -71477 -28858 -71473 -28562
rect -71473 -28858 -71177 -28562
rect -71177 -28858 -71173 -28562
rect -71477 -28862 -71173 -28858
rect -70477 -28562 -70173 -28558
rect -70477 -28858 -70473 -28562
rect -70473 -28858 -70177 -28562
rect -70177 -28858 -70173 -28562
rect -70477 -28862 -70173 -28858
rect -69477 -28562 -69173 -28558
rect -69477 -28858 -69473 -28562
rect -69473 -28858 -69177 -28562
rect -69177 -28858 -69173 -28562
rect -69477 -28862 -69173 -28858
rect -68477 -28562 -68173 -28558
rect -68477 -28858 -68473 -28562
rect -68473 -28858 -68177 -28562
rect -68177 -28858 -68173 -28562
rect -68477 -28862 -68173 -28858
rect -67477 -28562 -67173 -28558
rect -67477 -28858 -67473 -28562
rect -67473 -28858 -67177 -28562
rect -67177 -28858 -67173 -28562
rect -67477 -28862 -67173 -28858
rect -66477 -28562 -66173 -28558
rect -66477 -28858 -66473 -28562
rect -66473 -28858 -66177 -28562
rect -66177 -28858 -66173 -28562
rect -66477 -28862 -66173 -28858
rect -65477 -28562 -65173 -28558
rect -65477 -28858 -65473 -28562
rect -65473 -28858 -65177 -28562
rect -65177 -28858 -65173 -28562
rect -65477 -28862 -65173 -28858
rect -64477 -28562 -64173 -28558
rect -64477 -28858 -64473 -28562
rect -64473 -28858 -64177 -28562
rect -64177 -28858 -64173 -28562
rect -64477 -28862 -64173 -28858
rect -63477 -28562 -63173 -28558
rect -63477 -28858 -63473 -28562
rect -63473 -28858 -63177 -28562
rect -63177 -28858 -63173 -28562
rect -63477 -28862 -63173 -28858
rect -62477 -28562 -62173 -28558
rect -62477 -28858 -62473 -28562
rect -62473 -28858 -62177 -28562
rect -62177 -28858 -62173 -28562
rect -62477 -28862 -62173 -28858
rect -61477 -28562 -61173 -28558
rect -61477 -28858 -61473 -28562
rect -61473 -28858 -61177 -28562
rect -61177 -28858 -61173 -28562
rect -61477 -28862 -61173 -28858
rect -60477 -28562 -60173 -28558
rect -60477 -28858 -60473 -28562
rect -60473 -28858 -60177 -28562
rect -60177 -28858 -60173 -28562
rect -60477 -28862 -60173 -28858
rect -59477 -28562 -59173 -28558
rect -59477 -28858 -59473 -28562
rect -59473 -28858 -59177 -28562
rect -59177 -28858 -59173 -28562
rect -59477 -28862 -59173 -28858
rect -58477 -28562 -58173 -28558
rect -58477 -28858 -58473 -28562
rect -58473 -28858 -58177 -28562
rect -58177 -28858 -58173 -28562
rect -58477 -28862 -58173 -28858
rect -57477 -28562 -57173 -28558
rect -57477 -28858 -57473 -28562
rect -57473 -28858 -57177 -28562
rect -57177 -28858 -57173 -28562
rect -57477 -28862 -57173 -28858
rect -56477 -28562 -56173 -28558
rect -56477 -28858 -56473 -28562
rect -56473 -28858 -56177 -28562
rect -56177 -28858 -56173 -28562
rect -56477 -28862 -56173 -28858
rect -55477 -28562 -55173 -28558
rect -55477 -28858 -55473 -28562
rect -55473 -28858 -55177 -28562
rect -55177 -28858 -55173 -28562
rect -55477 -28862 -55173 -28858
rect -54477 -28562 -54173 -28558
rect -54477 -28858 -54473 -28562
rect -54473 -28858 -54177 -28562
rect -54177 -28858 -54173 -28562
rect -54477 -28862 -54173 -28858
rect -53477 -28562 -53173 -28558
rect -53477 -28858 -53473 -28562
rect -53473 -28858 -53177 -28562
rect -53177 -28858 -53173 -28562
rect -53477 -28862 -53173 -28858
rect -52477 -28562 -52173 -28558
rect -52477 -28858 -52473 -28562
rect -52473 -28858 -52177 -28562
rect -52177 -28858 -52173 -28562
rect -52477 -28862 -52173 -28858
rect -51477 -28562 -51173 -28558
rect -51477 -28858 -51473 -28562
rect -51473 -28858 -51177 -28562
rect -51177 -28858 -51173 -28562
rect -51477 -28862 -51173 -28858
rect -50477 -28562 -50173 -28558
rect -50477 -28858 -50473 -28562
rect -50473 -28858 -50177 -28562
rect -50177 -28858 -50173 -28562
rect -50477 -28862 -50173 -28858
rect -49477 -28562 -49173 -28558
rect -49477 -28858 -49473 -28562
rect -49473 -28858 -49177 -28562
rect -49177 -28858 -49173 -28562
rect -49477 -28862 -49173 -28858
rect 8623 -28562 8927 -28558
rect 8623 -28858 8627 -28562
rect 8627 -28858 8923 -28562
rect 8923 -28858 8927 -28562
rect 8623 -28862 8927 -28858
rect 9623 -28562 9927 -28558
rect 9623 -28858 9627 -28562
rect 9627 -28858 9923 -28562
rect 9923 -28858 9927 -28562
rect 9623 -28862 9927 -28858
rect 10623 -28562 10927 -28558
rect 10623 -28858 10627 -28562
rect 10627 -28858 10923 -28562
rect 10923 -28858 10927 -28562
rect 10623 -28862 10927 -28858
rect 11623 -28562 11927 -28558
rect 11623 -28858 11627 -28562
rect 11627 -28858 11923 -28562
rect 11923 -28858 11927 -28562
rect 11623 -28862 11927 -28858
rect 12623 -28562 12927 -28558
rect 12623 -28858 12627 -28562
rect 12627 -28858 12923 -28562
rect 12923 -28858 12927 -28562
rect 12623 -28862 12927 -28858
rect 13623 -28562 13927 -28558
rect 13623 -28858 13627 -28562
rect 13627 -28858 13923 -28562
rect 13923 -28858 13927 -28562
rect 13623 -28862 13927 -28858
rect 14623 -28562 14927 -28558
rect 14623 -28858 14627 -28562
rect 14627 -28858 14923 -28562
rect 14923 -28858 14927 -28562
rect 14623 -28862 14927 -28858
rect 15623 -28562 15927 -28558
rect 15623 -28858 15627 -28562
rect 15627 -28858 15923 -28562
rect 15923 -28858 15927 -28562
rect 15623 -28862 15927 -28858
rect 16623 -28562 16927 -28558
rect 16623 -28858 16627 -28562
rect 16627 -28858 16923 -28562
rect 16923 -28858 16927 -28562
rect 16623 -28862 16927 -28858
rect 17623 -28562 17927 -28558
rect 17623 -28858 17627 -28562
rect 17627 -28858 17923 -28562
rect 17923 -28858 17927 -28562
rect 17623 -28862 17927 -28858
rect 18623 -28562 18927 -28558
rect 18623 -28858 18627 -28562
rect 18627 -28858 18923 -28562
rect 18923 -28858 18927 -28562
rect 18623 -28862 18927 -28858
rect 19623 -28562 19927 -28558
rect 19623 -28858 19627 -28562
rect 19627 -28858 19923 -28562
rect 19923 -28858 19927 -28562
rect 19623 -28862 19927 -28858
rect 20623 -28562 20927 -28558
rect 20623 -28858 20627 -28562
rect 20627 -28858 20923 -28562
rect 20923 -28858 20927 -28562
rect 20623 -28862 20927 -28858
rect 21623 -28562 21927 -28558
rect 21623 -28858 21627 -28562
rect 21627 -28858 21923 -28562
rect 21923 -28858 21927 -28562
rect 21623 -28862 21927 -28858
rect 22623 -28562 22927 -28558
rect 22623 -28858 22627 -28562
rect 22627 -28858 22923 -28562
rect 22923 -28858 22927 -28562
rect 22623 -28862 22927 -28858
rect 23623 -28562 23927 -28558
rect 23623 -28858 23627 -28562
rect 23627 -28858 23923 -28562
rect 23923 -28858 23927 -28562
rect 23623 -28862 23927 -28858
rect 24623 -28562 24927 -28558
rect 24623 -28858 24627 -28562
rect 24627 -28858 24923 -28562
rect 24923 -28858 24927 -28562
rect 24623 -28862 24927 -28858
rect 25623 -28562 25927 -28558
rect 25623 -28858 25627 -28562
rect 25627 -28858 25923 -28562
rect 25923 -28858 25927 -28562
rect 25623 -28862 25927 -28858
rect 26623 -28562 26927 -28558
rect 26623 -28858 26627 -28562
rect 26627 -28858 26923 -28562
rect 26923 -28858 26927 -28562
rect 26623 -28862 26927 -28858
rect 27623 -28562 27927 -28558
rect 27623 -28858 27627 -28562
rect 27627 -28858 27923 -28562
rect 27923 -28858 27927 -28562
rect 27623 -28862 27927 -28858
rect 28623 -28562 28927 -28558
rect 28623 -28858 28627 -28562
rect 28627 -28858 28923 -28562
rect 28923 -28858 28927 -28562
rect 28623 -28862 28927 -28858
rect 29623 -28562 29927 -28558
rect 29623 -28858 29627 -28562
rect 29627 -28858 29923 -28562
rect 29923 -28858 29927 -28562
rect 29623 -28862 29927 -28858
rect 30623 -28562 30927 -28558
rect 30623 -28858 30627 -28562
rect 30627 -28858 30923 -28562
rect 30923 -28858 30927 -28562
rect 30623 -28862 30927 -28858
rect 31623 -28562 31927 -28558
rect 31623 -28858 31627 -28562
rect 31627 -28858 31923 -28562
rect 31923 -28858 31927 -28562
rect 31623 -28862 31927 -28858
rect 32623 -28562 32927 -28558
rect 32623 -28858 32627 -28562
rect 32627 -28858 32923 -28562
rect 32923 -28858 32927 -28562
rect 32623 -28862 32927 -28858
rect 33623 -28562 33927 -28558
rect 33623 -28858 33627 -28562
rect 33627 -28858 33923 -28562
rect 33923 -28858 33927 -28562
rect 33623 -28862 33927 -28858
rect -74817 -28902 -74513 -28898
rect -74817 -29198 -74813 -28902
rect -74813 -29198 -74517 -28902
rect -74517 -29198 -74513 -28902
rect -74817 -29202 -74513 -29198
rect -74477 -28902 -74173 -28898
rect -74477 -29198 -74473 -28902
rect -74473 -29198 -74177 -28902
rect -74177 -29198 -74173 -28902
rect -74477 -29202 -74173 -29198
rect -74137 -28902 -73513 -28898
rect -74137 -29198 -74133 -28902
rect -74133 -29198 -73517 -28902
rect -73517 -29198 -73513 -28902
rect -74137 -29202 -73513 -29198
rect -73477 -28902 -73173 -28898
rect -73477 -29198 -73473 -28902
rect -73473 -29198 -73177 -28902
rect -73177 -29198 -73173 -28902
rect -73477 -29202 -73173 -29198
rect -73137 -28902 -72513 -28898
rect -73137 -29198 -73133 -28902
rect -73133 -29198 -72517 -28902
rect -72517 -29198 -72513 -28902
rect -73137 -29202 -72513 -29198
rect -72477 -28902 -72173 -28898
rect -72477 -29198 -72473 -28902
rect -72473 -29198 -72177 -28902
rect -72177 -29198 -72173 -28902
rect -72477 -29202 -72173 -29198
rect -72137 -28902 -71513 -28898
rect -72137 -29198 -72133 -28902
rect -72133 -29198 -71517 -28902
rect -71517 -29198 -71513 -28902
rect -72137 -29202 -71513 -29198
rect -71477 -28902 -71173 -28898
rect -71477 -29198 -71473 -28902
rect -71473 -29198 -71177 -28902
rect -71177 -29198 -71173 -28902
rect -71477 -29202 -71173 -29198
rect -71137 -28902 -70513 -28898
rect -71137 -29198 -71133 -28902
rect -71133 -29198 -70517 -28902
rect -70517 -29198 -70513 -28902
rect -71137 -29202 -70513 -29198
rect -70477 -28902 -70173 -28898
rect -70477 -29198 -70473 -28902
rect -70473 -29198 -70177 -28902
rect -70177 -29198 -70173 -28902
rect -70477 -29202 -70173 -29198
rect -70137 -28902 -69513 -28898
rect -70137 -29198 -70133 -28902
rect -70133 -29198 -69517 -28902
rect -69517 -29198 -69513 -28902
rect -70137 -29202 -69513 -29198
rect -69477 -28902 -69173 -28898
rect -69477 -29198 -69473 -28902
rect -69473 -29198 -69177 -28902
rect -69177 -29198 -69173 -28902
rect -69477 -29202 -69173 -29198
rect -69137 -28902 -68513 -28898
rect -69137 -29198 -69133 -28902
rect -69133 -29198 -68517 -28902
rect -68517 -29198 -68513 -28902
rect -69137 -29202 -68513 -29198
rect -68477 -28902 -68173 -28898
rect -68477 -29198 -68473 -28902
rect -68473 -29198 -68177 -28902
rect -68177 -29198 -68173 -28902
rect -68477 -29202 -68173 -29198
rect -68137 -28902 -67513 -28898
rect -68137 -29198 -68133 -28902
rect -68133 -29198 -67517 -28902
rect -67517 -29198 -67513 -28902
rect -68137 -29202 -67513 -29198
rect -67477 -28902 -67173 -28898
rect -67477 -29198 -67473 -28902
rect -67473 -29198 -67177 -28902
rect -67177 -29198 -67173 -28902
rect -67477 -29202 -67173 -29198
rect -67137 -28902 -66513 -28898
rect -67137 -29198 -67133 -28902
rect -67133 -29198 -66517 -28902
rect -66517 -29198 -66513 -28902
rect -67137 -29202 -66513 -29198
rect -66477 -28902 -66173 -28898
rect -66477 -29198 -66473 -28902
rect -66473 -29198 -66177 -28902
rect -66177 -29198 -66173 -28902
rect -66477 -29202 -66173 -29198
rect -66137 -28902 -65513 -28898
rect -66137 -29198 -66133 -28902
rect -66133 -29198 -65517 -28902
rect -65517 -29198 -65513 -28902
rect -66137 -29202 -65513 -29198
rect -65477 -28902 -65173 -28898
rect -65477 -29198 -65473 -28902
rect -65473 -29198 -65177 -28902
rect -65177 -29198 -65173 -28902
rect -65477 -29202 -65173 -29198
rect -65137 -28902 -64513 -28898
rect -65137 -29198 -65133 -28902
rect -65133 -29198 -64517 -28902
rect -64517 -29198 -64513 -28902
rect -65137 -29202 -64513 -29198
rect -64477 -28902 -64173 -28898
rect -64477 -29198 -64473 -28902
rect -64473 -29198 -64177 -28902
rect -64177 -29198 -64173 -28902
rect -64477 -29202 -64173 -29198
rect -64137 -28902 -63513 -28898
rect -64137 -29198 -64133 -28902
rect -64133 -29198 -63517 -28902
rect -63517 -29198 -63513 -28902
rect -64137 -29202 -63513 -29198
rect -63477 -28902 -63173 -28898
rect -63477 -29198 -63473 -28902
rect -63473 -29198 -63177 -28902
rect -63177 -29198 -63173 -28902
rect -63477 -29202 -63173 -29198
rect -63137 -28902 -62513 -28898
rect -63137 -29198 -63133 -28902
rect -63133 -29198 -62517 -28902
rect -62517 -29198 -62513 -28902
rect -63137 -29202 -62513 -29198
rect -62477 -28902 -62173 -28898
rect -62477 -29198 -62473 -28902
rect -62473 -29198 -62177 -28902
rect -62177 -29198 -62173 -28902
rect -62477 -29202 -62173 -29198
rect -62137 -28902 -61513 -28898
rect -62137 -29198 -62133 -28902
rect -62133 -29198 -61517 -28902
rect -61517 -29198 -61513 -28902
rect -62137 -29202 -61513 -29198
rect -61477 -28902 -61173 -28898
rect -61477 -29198 -61473 -28902
rect -61473 -29198 -61177 -28902
rect -61177 -29198 -61173 -28902
rect -61477 -29202 -61173 -29198
rect -61137 -28902 -60513 -28898
rect -61137 -29198 -61133 -28902
rect -61133 -29198 -60517 -28902
rect -60517 -29198 -60513 -28902
rect -61137 -29202 -60513 -29198
rect -60477 -28902 -60173 -28898
rect -60477 -29198 -60473 -28902
rect -60473 -29198 -60177 -28902
rect -60177 -29198 -60173 -28902
rect -60477 -29202 -60173 -29198
rect -60137 -28902 -59513 -28898
rect -60137 -29198 -60133 -28902
rect -60133 -29198 -59517 -28902
rect -59517 -29198 -59513 -28902
rect -60137 -29202 -59513 -29198
rect -59477 -28902 -59173 -28898
rect -59477 -29198 -59473 -28902
rect -59473 -29198 -59177 -28902
rect -59177 -29198 -59173 -28902
rect -59477 -29202 -59173 -29198
rect -59137 -28902 -58513 -28898
rect -59137 -29198 -59133 -28902
rect -59133 -29198 -58517 -28902
rect -58517 -29198 -58513 -28902
rect -59137 -29202 -58513 -29198
rect -58477 -28902 -58173 -28898
rect -58477 -29198 -58473 -28902
rect -58473 -29198 -58177 -28902
rect -58177 -29198 -58173 -28902
rect -58477 -29202 -58173 -29198
rect -58137 -28902 -57513 -28898
rect -58137 -29198 -58133 -28902
rect -58133 -29198 -57517 -28902
rect -57517 -29198 -57513 -28902
rect -58137 -29202 -57513 -29198
rect -57477 -28902 -57173 -28898
rect -57477 -29198 -57473 -28902
rect -57473 -29198 -57177 -28902
rect -57177 -29198 -57173 -28902
rect -57477 -29202 -57173 -29198
rect -57137 -28902 -56513 -28898
rect -57137 -29198 -57133 -28902
rect -57133 -29198 -56517 -28902
rect -56517 -29198 -56513 -28902
rect -57137 -29202 -56513 -29198
rect -56477 -28902 -56173 -28898
rect -56477 -29198 -56473 -28902
rect -56473 -29198 -56177 -28902
rect -56177 -29198 -56173 -28902
rect -56477 -29202 -56173 -29198
rect -56137 -28902 -55513 -28898
rect -56137 -29198 -56133 -28902
rect -56133 -29198 -55517 -28902
rect -55517 -29198 -55513 -28902
rect -56137 -29202 -55513 -29198
rect -55477 -28902 -55173 -28898
rect -55477 -29198 -55473 -28902
rect -55473 -29198 -55177 -28902
rect -55177 -29198 -55173 -28902
rect -55477 -29202 -55173 -29198
rect -55137 -28902 -54513 -28898
rect -55137 -29198 -55133 -28902
rect -55133 -29198 -54517 -28902
rect -54517 -29198 -54513 -28902
rect -55137 -29202 -54513 -29198
rect -54477 -28902 -54173 -28898
rect -54477 -29198 -54473 -28902
rect -54473 -29198 -54177 -28902
rect -54177 -29198 -54173 -28902
rect -54477 -29202 -54173 -29198
rect -54137 -28902 -53513 -28898
rect -54137 -29198 -54133 -28902
rect -54133 -29198 -53517 -28902
rect -53517 -29198 -53513 -28902
rect -54137 -29202 -53513 -29198
rect -53477 -28902 -53173 -28898
rect -53477 -29198 -53473 -28902
rect -53473 -29198 -53177 -28902
rect -53177 -29198 -53173 -28902
rect -53477 -29202 -53173 -29198
rect -53137 -28902 -52513 -28898
rect -53137 -29198 -53133 -28902
rect -53133 -29198 -52517 -28902
rect -52517 -29198 -52513 -28902
rect -53137 -29202 -52513 -29198
rect -52477 -28902 -52173 -28898
rect -52477 -29198 -52473 -28902
rect -52473 -29198 -52177 -28902
rect -52177 -29198 -52173 -28902
rect -52477 -29202 -52173 -29198
rect -52137 -28902 -51513 -28898
rect -52137 -29198 -52133 -28902
rect -52133 -29198 -51517 -28902
rect -51517 -29198 -51513 -28902
rect -52137 -29202 -51513 -29198
rect -51477 -28902 -51173 -28898
rect -51477 -29198 -51473 -28902
rect -51473 -29198 -51177 -28902
rect -51177 -29198 -51173 -28902
rect -51477 -29202 -51173 -29198
rect -51137 -28902 -50513 -28898
rect -51137 -29198 -51133 -28902
rect -51133 -29198 -50517 -28902
rect -50517 -29198 -50513 -28902
rect -51137 -29202 -50513 -29198
rect -50477 -28902 -50173 -28898
rect -50477 -29198 -50473 -28902
rect -50473 -29198 -50177 -28902
rect -50177 -29198 -50173 -28902
rect -50477 -29202 -50173 -29198
rect -50137 -28902 -49513 -28898
rect -50137 -29198 -50133 -28902
rect -50133 -29198 -49517 -28902
rect -49517 -29198 -49513 -28902
rect -50137 -29202 -49513 -29198
rect -49477 -28902 -49173 -28898
rect -49477 -29198 -49473 -28902
rect -49473 -29198 -49177 -28902
rect -49177 -29198 -49173 -28902
rect -49477 -29202 -49173 -29198
rect -49137 -28902 -48833 -28898
rect -49137 -29198 -49133 -28902
rect -49133 -29198 -48837 -28902
rect -48837 -29198 -48833 -28902
rect -49137 -29202 -48833 -29198
rect 8283 -28902 8587 -28898
rect 8283 -29198 8287 -28902
rect 8287 -29198 8583 -28902
rect 8583 -29198 8587 -28902
rect 8283 -29202 8587 -29198
rect 8623 -28902 8927 -28898
rect 8623 -29198 8627 -28902
rect 8627 -29198 8923 -28902
rect 8923 -29198 8927 -28902
rect 8623 -29202 8927 -29198
rect 8963 -28902 9587 -28898
rect 8963 -29198 8967 -28902
rect 8967 -29198 9583 -28902
rect 9583 -29198 9587 -28902
rect 8963 -29202 9587 -29198
rect 9623 -28902 9927 -28898
rect 9623 -29198 9627 -28902
rect 9627 -29198 9923 -28902
rect 9923 -29198 9927 -28902
rect 9623 -29202 9927 -29198
rect 9963 -28902 10587 -28898
rect 9963 -29198 9967 -28902
rect 9967 -29198 10583 -28902
rect 10583 -29198 10587 -28902
rect 9963 -29202 10587 -29198
rect 10623 -28902 10927 -28898
rect 10623 -29198 10627 -28902
rect 10627 -29198 10923 -28902
rect 10923 -29198 10927 -28902
rect 10623 -29202 10927 -29198
rect 10963 -28902 11587 -28898
rect 10963 -29198 10967 -28902
rect 10967 -29198 11583 -28902
rect 11583 -29198 11587 -28902
rect 10963 -29202 11587 -29198
rect 11623 -28902 11927 -28898
rect 11623 -29198 11627 -28902
rect 11627 -29198 11923 -28902
rect 11923 -29198 11927 -28902
rect 11623 -29202 11927 -29198
rect 11963 -28902 12587 -28898
rect 11963 -29198 11967 -28902
rect 11967 -29198 12583 -28902
rect 12583 -29198 12587 -28902
rect 11963 -29202 12587 -29198
rect 12623 -28902 12927 -28898
rect 12623 -29198 12627 -28902
rect 12627 -29198 12923 -28902
rect 12923 -29198 12927 -28902
rect 12623 -29202 12927 -29198
rect 12963 -28902 13587 -28898
rect 12963 -29198 12967 -28902
rect 12967 -29198 13583 -28902
rect 13583 -29198 13587 -28902
rect 12963 -29202 13587 -29198
rect 13623 -28902 13927 -28898
rect 13623 -29198 13627 -28902
rect 13627 -29198 13923 -28902
rect 13923 -29198 13927 -28902
rect 13623 -29202 13927 -29198
rect 13963 -28902 14587 -28898
rect 13963 -29198 13967 -28902
rect 13967 -29198 14583 -28902
rect 14583 -29198 14587 -28902
rect 13963 -29202 14587 -29198
rect 14623 -28902 14927 -28898
rect 14623 -29198 14627 -28902
rect 14627 -29198 14923 -28902
rect 14923 -29198 14927 -28902
rect 14623 -29202 14927 -29198
rect 14963 -28902 15587 -28898
rect 14963 -29198 14967 -28902
rect 14967 -29198 15583 -28902
rect 15583 -29198 15587 -28902
rect 14963 -29202 15587 -29198
rect 15623 -28902 15927 -28898
rect 15623 -29198 15627 -28902
rect 15627 -29198 15923 -28902
rect 15923 -29198 15927 -28902
rect 15623 -29202 15927 -29198
rect 15963 -28902 16587 -28898
rect 15963 -29198 15967 -28902
rect 15967 -29198 16583 -28902
rect 16583 -29198 16587 -28902
rect 15963 -29202 16587 -29198
rect 16623 -28902 16927 -28898
rect 16623 -29198 16627 -28902
rect 16627 -29198 16923 -28902
rect 16923 -29198 16927 -28902
rect 16623 -29202 16927 -29198
rect 16963 -28902 17587 -28898
rect 16963 -29198 16967 -28902
rect 16967 -29198 17583 -28902
rect 17583 -29198 17587 -28902
rect 16963 -29202 17587 -29198
rect 17623 -28902 17927 -28898
rect 17623 -29198 17627 -28902
rect 17627 -29198 17923 -28902
rect 17923 -29198 17927 -28902
rect 17623 -29202 17927 -29198
rect 17963 -28902 18587 -28898
rect 17963 -29198 17967 -28902
rect 17967 -29198 18583 -28902
rect 18583 -29198 18587 -28902
rect 17963 -29202 18587 -29198
rect 18623 -28902 18927 -28898
rect 18623 -29198 18627 -28902
rect 18627 -29198 18923 -28902
rect 18923 -29198 18927 -28902
rect 18623 -29202 18927 -29198
rect 18963 -28902 19587 -28898
rect 18963 -29198 18967 -28902
rect 18967 -29198 19583 -28902
rect 19583 -29198 19587 -28902
rect 18963 -29202 19587 -29198
rect 19623 -28902 19927 -28898
rect 19623 -29198 19627 -28902
rect 19627 -29198 19923 -28902
rect 19923 -29198 19927 -28902
rect 19623 -29202 19927 -29198
rect 19963 -28902 20587 -28898
rect 19963 -29198 19967 -28902
rect 19967 -29198 20583 -28902
rect 20583 -29198 20587 -28902
rect 19963 -29202 20587 -29198
rect 20623 -28902 20927 -28898
rect 20623 -29198 20627 -28902
rect 20627 -29198 20923 -28902
rect 20923 -29198 20927 -28902
rect 20623 -29202 20927 -29198
rect 20963 -28902 21587 -28898
rect 20963 -29198 20967 -28902
rect 20967 -29198 21583 -28902
rect 21583 -29198 21587 -28902
rect 20963 -29202 21587 -29198
rect 21623 -28902 21927 -28898
rect 21623 -29198 21627 -28902
rect 21627 -29198 21923 -28902
rect 21923 -29198 21927 -28902
rect 21623 -29202 21927 -29198
rect 21963 -28902 22587 -28898
rect 21963 -29198 21967 -28902
rect 21967 -29198 22583 -28902
rect 22583 -29198 22587 -28902
rect 21963 -29202 22587 -29198
rect 22623 -28902 22927 -28898
rect 22623 -29198 22627 -28902
rect 22627 -29198 22923 -28902
rect 22923 -29198 22927 -28902
rect 22623 -29202 22927 -29198
rect 22963 -28902 23587 -28898
rect 22963 -29198 22967 -28902
rect 22967 -29198 23583 -28902
rect 23583 -29198 23587 -28902
rect 22963 -29202 23587 -29198
rect 23623 -28902 23927 -28898
rect 23623 -29198 23627 -28902
rect 23627 -29198 23923 -28902
rect 23923 -29198 23927 -28902
rect 23623 -29202 23927 -29198
rect 23963 -28902 24587 -28898
rect 23963 -29198 23967 -28902
rect 23967 -29198 24583 -28902
rect 24583 -29198 24587 -28902
rect 23963 -29202 24587 -29198
rect 24623 -28902 24927 -28898
rect 24623 -29198 24627 -28902
rect 24627 -29198 24923 -28902
rect 24923 -29198 24927 -28902
rect 24623 -29202 24927 -29198
rect 24963 -28902 25587 -28898
rect 24963 -29198 24967 -28902
rect 24967 -29198 25583 -28902
rect 25583 -29198 25587 -28902
rect 24963 -29202 25587 -29198
rect 25623 -28902 25927 -28898
rect 25623 -29198 25627 -28902
rect 25627 -29198 25923 -28902
rect 25923 -29198 25927 -28902
rect 25623 -29202 25927 -29198
rect 25963 -28902 26587 -28898
rect 25963 -29198 25967 -28902
rect 25967 -29198 26583 -28902
rect 26583 -29198 26587 -28902
rect 25963 -29202 26587 -29198
rect 26623 -28902 26927 -28898
rect 26623 -29198 26627 -28902
rect 26627 -29198 26923 -28902
rect 26923 -29198 26927 -28902
rect 26623 -29202 26927 -29198
rect 26963 -28902 27587 -28898
rect 26963 -29198 26967 -28902
rect 26967 -29198 27583 -28902
rect 27583 -29198 27587 -28902
rect 26963 -29202 27587 -29198
rect 27623 -28902 27927 -28898
rect 27623 -29198 27627 -28902
rect 27627 -29198 27923 -28902
rect 27923 -29198 27927 -28902
rect 27623 -29202 27927 -29198
rect 27963 -28902 28587 -28898
rect 27963 -29198 27967 -28902
rect 27967 -29198 28583 -28902
rect 28583 -29198 28587 -28902
rect 27963 -29202 28587 -29198
rect 28623 -28902 28927 -28898
rect 28623 -29198 28627 -28902
rect 28627 -29198 28923 -28902
rect 28923 -29198 28927 -28902
rect 28623 -29202 28927 -29198
rect 28963 -28902 29587 -28898
rect 28963 -29198 28967 -28902
rect 28967 -29198 29583 -28902
rect 29583 -29198 29587 -28902
rect 28963 -29202 29587 -29198
rect 29623 -28902 29927 -28898
rect 29623 -29198 29627 -28902
rect 29627 -29198 29923 -28902
rect 29923 -29198 29927 -28902
rect 29623 -29202 29927 -29198
rect 29963 -28902 30587 -28898
rect 29963 -29198 29967 -28902
rect 29967 -29198 30583 -28902
rect 30583 -29198 30587 -28902
rect 29963 -29202 30587 -29198
rect 30623 -28902 30927 -28898
rect 30623 -29198 30627 -28902
rect 30627 -29198 30923 -28902
rect 30923 -29198 30927 -28902
rect 30623 -29202 30927 -29198
rect 30963 -28902 31587 -28898
rect 30963 -29198 30967 -28902
rect 30967 -29198 31583 -28902
rect 31583 -29198 31587 -28902
rect 30963 -29202 31587 -29198
rect 31623 -28902 31927 -28898
rect 31623 -29198 31627 -28902
rect 31627 -29198 31923 -28902
rect 31923 -29198 31927 -28902
rect 31623 -29202 31927 -29198
rect 31963 -28902 32587 -28898
rect 31963 -29198 31967 -28902
rect 31967 -29198 32583 -28902
rect 32583 -29198 32587 -28902
rect 31963 -29202 32587 -29198
rect 32623 -28902 32927 -28898
rect 32623 -29198 32627 -28902
rect 32627 -29198 32923 -28902
rect 32923 -29198 32927 -28902
rect 32623 -29202 32927 -29198
rect 32963 -28902 33587 -28898
rect 32963 -29198 32967 -28902
rect 32967 -29198 33583 -28902
rect 33583 -29198 33587 -28902
rect 32963 -29202 33587 -29198
rect 33623 -28902 33927 -28898
rect 33623 -29198 33627 -28902
rect 33627 -29198 33923 -28902
rect 33923 -29198 33927 -28902
rect 33623 -29202 33927 -29198
rect 33963 -28902 34267 -28898
rect 33963 -29198 33967 -28902
rect 33967 -29198 34263 -28902
rect 34263 -29198 34267 -28902
rect 33963 -29202 34267 -29198
rect -74477 -29242 -74173 -29238
rect -74477 -29858 -74473 -29242
rect -74473 -29858 -74177 -29242
rect -74177 -29858 -74173 -29242
rect -74477 -29862 -74173 -29858
rect -73477 -29242 -73173 -29238
rect -73477 -29858 -73473 -29242
rect -73473 -29858 -73177 -29242
rect -73177 -29858 -73173 -29242
rect -73477 -29862 -73173 -29858
rect -72477 -29242 -72173 -29238
rect -72477 -29858 -72473 -29242
rect -72473 -29858 -72177 -29242
rect -72177 -29858 -72173 -29242
rect -72477 -29862 -72173 -29858
rect -71477 -29242 -71173 -29238
rect -71477 -29858 -71473 -29242
rect -71473 -29858 -71177 -29242
rect -71177 -29858 -71173 -29242
rect -71477 -29862 -71173 -29858
rect -70477 -29242 -70173 -29238
rect -70477 -29858 -70473 -29242
rect -70473 -29858 -70177 -29242
rect -70177 -29858 -70173 -29242
rect -70477 -29862 -70173 -29858
rect -69477 -29242 -69173 -29238
rect -69477 -29858 -69473 -29242
rect -69473 -29858 -69177 -29242
rect -69177 -29858 -69173 -29242
rect -69477 -29862 -69173 -29858
rect -68477 -29242 -68173 -29238
rect -68477 -29858 -68473 -29242
rect -68473 -29858 -68177 -29242
rect -68177 -29858 -68173 -29242
rect -68477 -29862 -68173 -29858
rect -67477 -29242 -67173 -29238
rect -67477 -29858 -67473 -29242
rect -67473 -29858 -67177 -29242
rect -67177 -29858 -67173 -29242
rect -67477 -29862 -67173 -29858
rect -66477 -29242 -66173 -29238
rect -66477 -29858 -66473 -29242
rect -66473 -29858 -66177 -29242
rect -66177 -29858 -66173 -29242
rect -66477 -29862 -66173 -29858
rect -65477 -29242 -65173 -29238
rect -65477 -29858 -65473 -29242
rect -65473 -29858 -65177 -29242
rect -65177 -29858 -65173 -29242
rect -65477 -29862 -65173 -29858
rect -64477 -29242 -64173 -29238
rect -64477 -29858 -64473 -29242
rect -64473 -29858 -64177 -29242
rect -64177 -29858 -64173 -29242
rect -64477 -29862 -64173 -29858
rect -63477 -29242 -63173 -29238
rect -63477 -29858 -63473 -29242
rect -63473 -29858 -63177 -29242
rect -63177 -29858 -63173 -29242
rect -63477 -29862 -63173 -29858
rect -62477 -29242 -62173 -29238
rect -62477 -29858 -62473 -29242
rect -62473 -29858 -62177 -29242
rect -62177 -29858 -62173 -29242
rect -62477 -29862 -62173 -29858
rect -61477 -29242 -61173 -29238
rect -61477 -29858 -61473 -29242
rect -61473 -29858 -61177 -29242
rect -61177 -29858 -61173 -29242
rect -61477 -29862 -61173 -29858
rect -60477 -29242 -60173 -29238
rect -60477 -29858 -60473 -29242
rect -60473 -29858 -60177 -29242
rect -60177 -29858 -60173 -29242
rect -60477 -29862 -60173 -29858
rect -59477 -29242 -59173 -29238
rect -59477 -29858 -59473 -29242
rect -59473 -29858 -59177 -29242
rect -59177 -29858 -59173 -29242
rect -59477 -29862 -59173 -29858
rect -58477 -29242 -58173 -29238
rect -58477 -29858 -58473 -29242
rect -58473 -29858 -58177 -29242
rect -58177 -29858 -58173 -29242
rect -58477 -29862 -58173 -29858
rect -57477 -29242 -57173 -29238
rect -57477 -29858 -57473 -29242
rect -57473 -29858 -57177 -29242
rect -57177 -29858 -57173 -29242
rect -57477 -29862 -57173 -29858
rect -56477 -29242 -56173 -29238
rect -56477 -29858 -56473 -29242
rect -56473 -29858 -56177 -29242
rect -56177 -29858 -56173 -29242
rect -56477 -29862 -56173 -29858
rect -55477 -29242 -55173 -29238
rect -55477 -29858 -55473 -29242
rect -55473 -29858 -55177 -29242
rect -55177 -29858 -55173 -29242
rect -55477 -29862 -55173 -29858
rect -54477 -29242 -54173 -29238
rect -54477 -29858 -54473 -29242
rect -54473 -29858 -54177 -29242
rect -54177 -29858 -54173 -29242
rect -54477 -29862 -54173 -29858
rect -53477 -29242 -53173 -29238
rect -53477 -29858 -53473 -29242
rect -53473 -29858 -53177 -29242
rect -53177 -29858 -53173 -29242
rect -53477 -29862 -53173 -29858
rect -52477 -29242 -52173 -29238
rect -52477 -29858 -52473 -29242
rect -52473 -29858 -52177 -29242
rect -52177 -29858 -52173 -29242
rect -52477 -29862 -52173 -29858
rect -51477 -29242 -51173 -29238
rect -51477 -29858 -51473 -29242
rect -51473 -29858 -51177 -29242
rect -51177 -29858 -51173 -29242
rect -51477 -29862 -51173 -29858
rect -50477 -29242 -50173 -29238
rect -50477 -29858 -50473 -29242
rect -50473 -29858 -50177 -29242
rect -50177 -29858 -50173 -29242
rect -50477 -29862 -50173 -29858
rect -49477 -29242 -49173 -29238
rect -49477 -29858 -49473 -29242
rect -49473 -29858 -49177 -29242
rect -49177 -29858 -49173 -29242
rect -49477 -29862 -49173 -29858
rect 8623 -29242 8927 -29238
rect 8623 -29858 8627 -29242
rect 8627 -29858 8923 -29242
rect 8923 -29858 8927 -29242
rect 8623 -29862 8927 -29858
rect 9623 -29242 9927 -29238
rect 9623 -29858 9627 -29242
rect 9627 -29858 9923 -29242
rect 9923 -29858 9927 -29242
rect 9623 -29862 9927 -29858
rect 10623 -29242 10927 -29238
rect 10623 -29858 10627 -29242
rect 10627 -29858 10923 -29242
rect 10923 -29858 10927 -29242
rect 10623 -29862 10927 -29858
rect 11623 -29242 11927 -29238
rect 11623 -29858 11627 -29242
rect 11627 -29858 11923 -29242
rect 11923 -29858 11927 -29242
rect 11623 -29862 11927 -29858
rect 12623 -29242 12927 -29238
rect 12623 -29858 12627 -29242
rect 12627 -29858 12923 -29242
rect 12923 -29858 12927 -29242
rect 12623 -29862 12927 -29858
rect 13623 -29242 13927 -29238
rect 13623 -29858 13627 -29242
rect 13627 -29858 13923 -29242
rect 13923 -29858 13927 -29242
rect 13623 -29862 13927 -29858
rect 14623 -29242 14927 -29238
rect 14623 -29858 14627 -29242
rect 14627 -29858 14923 -29242
rect 14923 -29858 14927 -29242
rect 14623 -29862 14927 -29858
rect 15623 -29242 15927 -29238
rect 15623 -29858 15627 -29242
rect 15627 -29858 15923 -29242
rect 15923 -29858 15927 -29242
rect 15623 -29862 15927 -29858
rect 16623 -29242 16927 -29238
rect 16623 -29858 16627 -29242
rect 16627 -29858 16923 -29242
rect 16923 -29858 16927 -29242
rect 16623 -29862 16927 -29858
rect 17623 -29242 17927 -29238
rect 17623 -29858 17627 -29242
rect 17627 -29858 17923 -29242
rect 17923 -29858 17927 -29242
rect 17623 -29862 17927 -29858
rect 18623 -29242 18927 -29238
rect 18623 -29858 18627 -29242
rect 18627 -29858 18923 -29242
rect 18923 -29858 18927 -29242
rect 18623 -29862 18927 -29858
rect 19623 -29242 19927 -29238
rect 19623 -29858 19627 -29242
rect 19627 -29858 19923 -29242
rect 19923 -29858 19927 -29242
rect 19623 -29862 19927 -29858
rect 20623 -29242 20927 -29238
rect 20623 -29858 20627 -29242
rect 20627 -29858 20923 -29242
rect 20923 -29858 20927 -29242
rect 20623 -29862 20927 -29858
rect 21623 -29242 21927 -29238
rect 21623 -29858 21627 -29242
rect 21627 -29858 21923 -29242
rect 21923 -29858 21927 -29242
rect 21623 -29862 21927 -29858
rect 22623 -29242 22927 -29238
rect 22623 -29858 22627 -29242
rect 22627 -29858 22923 -29242
rect 22923 -29858 22927 -29242
rect 22623 -29862 22927 -29858
rect 23623 -29242 23927 -29238
rect 23623 -29858 23627 -29242
rect 23627 -29858 23923 -29242
rect 23923 -29858 23927 -29242
rect 23623 -29862 23927 -29858
rect 24623 -29242 24927 -29238
rect 24623 -29858 24627 -29242
rect 24627 -29858 24923 -29242
rect 24923 -29858 24927 -29242
rect 24623 -29862 24927 -29858
rect 25623 -29242 25927 -29238
rect 25623 -29858 25627 -29242
rect 25627 -29858 25923 -29242
rect 25923 -29858 25927 -29242
rect 25623 -29862 25927 -29858
rect 26623 -29242 26927 -29238
rect 26623 -29858 26627 -29242
rect 26627 -29858 26923 -29242
rect 26923 -29858 26927 -29242
rect 26623 -29862 26927 -29858
rect 27623 -29242 27927 -29238
rect 27623 -29858 27627 -29242
rect 27627 -29858 27923 -29242
rect 27923 -29858 27927 -29242
rect 27623 -29862 27927 -29858
rect 28623 -29242 28927 -29238
rect 28623 -29858 28627 -29242
rect 28627 -29858 28923 -29242
rect 28923 -29858 28927 -29242
rect 28623 -29862 28927 -29858
rect 29623 -29242 29927 -29238
rect 29623 -29858 29627 -29242
rect 29627 -29858 29923 -29242
rect 29923 -29858 29927 -29242
rect 29623 -29862 29927 -29858
rect 30623 -29242 30927 -29238
rect 30623 -29858 30627 -29242
rect 30627 -29858 30923 -29242
rect 30923 -29858 30927 -29242
rect 30623 -29862 30927 -29858
rect 31623 -29242 31927 -29238
rect 31623 -29858 31627 -29242
rect 31627 -29858 31923 -29242
rect 31923 -29858 31927 -29242
rect 31623 -29862 31927 -29858
rect 32623 -29242 32927 -29238
rect 32623 -29858 32627 -29242
rect 32627 -29858 32923 -29242
rect 32923 -29858 32927 -29242
rect 32623 -29862 32927 -29858
rect 33623 -29242 33927 -29238
rect 33623 -29858 33627 -29242
rect 33627 -29858 33923 -29242
rect 33923 -29858 33927 -29242
rect 33623 -29862 33927 -29858
rect -74817 -29902 -74513 -29898
rect -74817 -30198 -74813 -29902
rect -74813 -30198 -74517 -29902
rect -74517 -30198 -74513 -29902
rect -74817 -30202 -74513 -30198
rect -74477 -29902 -74173 -29898
rect -74477 -30198 -74473 -29902
rect -74473 -30198 -74177 -29902
rect -74177 -30198 -74173 -29902
rect -74477 -30202 -74173 -30198
rect -74137 -29902 -73513 -29898
rect -74137 -30198 -74133 -29902
rect -74133 -30198 -73517 -29902
rect -73517 -30198 -73513 -29902
rect -74137 -30202 -73513 -30198
rect -73477 -29902 -73173 -29898
rect -73477 -30198 -73473 -29902
rect -73473 -30198 -73177 -29902
rect -73177 -30198 -73173 -29902
rect -73477 -30202 -73173 -30198
rect -73137 -29902 -72513 -29898
rect -73137 -30198 -73133 -29902
rect -73133 -30198 -72517 -29902
rect -72517 -30198 -72513 -29902
rect -73137 -30202 -72513 -30198
rect -72477 -29902 -72173 -29898
rect -72477 -30198 -72473 -29902
rect -72473 -30198 -72177 -29902
rect -72177 -30198 -72173 -29902
rect -72477 -30202 -72173 -30198
rect -72137 -29902 -71513 -29898
rect -72137 -30198 -72133 -29902
rect -72133 -30198 -71517 -29902
rect -71517 -30198 -71513 -29902
rect -72137 -30202 -71513 -30198
rect -71477 -29902 -71173 -29898
rect -71477 -30198 -71473 -29902
rect -71473 -30198 -71177 -29902
rect -71177 -30198 -71173 -29902
rect -71477 -30202 -71173 -30198
rect -71137 -29902 -70513 -29898
rect -71137 -30198 -71133 -29902
rect -71133 -30198 -70517 -29902
rect -70517 -30198 -70513 -29902
rect -71137 -30202 -70513 -30198
rect -70477 -29902 -70173 -29898
rect -70477 -30198 -70473 -29902
rect -70473 -30198 -70177 -29902
rect -70177 -30198 -70173 -29902
rect -70477 -30202 -70173 -30198
rect -70137 -29902 -69513 -29898
rect -70137 -30198 -70133 -29902
rect -70133 -30198 -69517 -29902
rect -69517 -30198 -69513 -29902
rect -70137 -30202 -69513 -30198
rect -69477 -29902 -69173 -29898
rect -69477 -30198 -69473 -29902
rect -69473 -30198 -69177 -29902
rect -69177 -30198 -69173 -29902
rect -69477 -30202 -69173 -30198
rect -69137 -29902 -68513 -29898
rect -69137 -30198 -69133 -29902
rect -69133 -30198 -68517 -29902
rect -68517 -30198 -68513 -29902
rect -69137 -30202 -68513 -30198
rect -68477 -29902 -68173 -29898
rect -68477 -30198 -68473 -29902
rect -68473 -30198 -68177 -29902
rect -68177 -30198 -68173 -29902
rect -68477 -30202 -68173 -30198
rect -68137 -29902 -67513 -29898
rect -68137 -30198 -68133 -29902
rect -68133 -30198 -67517 -29902
rect -67517 -30198 -67513 -29902
rect -68137 -30202 -67513 -30198
rect -67477 -29902 -67173 -29898
rect -67477 -30198 -67473 -29902
rect -67473 -30198 -67177 -29902
rect -67177 -30198 -67173 -29902
rect -67477 -30202 -67173 -30198
rect -67137 -29902 -66513 -29898
rect -67137 -30198 -67133 -29902
rect -67133 -30198 -66517 -29902
rect -66517 -30198 -66513 -29902
rect -67137 -30202 -66513 -30198
rect -66477 -29902 -66173 -29898
rect -66477 -30198 -66473 -29902
rect -66473 -30198 -66177 -29902
rect -66177 -30198 -66173 -29902
rect -66477 -30202 -66173 -30198
rect -66137 -29902 -65513 -29898
rect -66137 -30198 -66133 -29902
rect -66133 -30198 -65517 -29902
rect -65517 -30198 -65513 -29902
rect -66137 -30202 -65513 -30198
rect -65477 -29902 -65173 -29898
rect -65477 -30198 -65473 -29902
rect -65473 -30198 -65177 -29902
rect -65177 -30198 -65173 -29902
rect -65477 -30202 -65173 -30198
rect -65137 -29902 -64513 -29898
rect -65137 -30198 -65133 -29902
rect -65133 -30198 -64517 -29902
rect -64517 -30198 -64513 -29902
rect -65137 -30202 -64513 -30198
rect -64477 -29902 -64173 -29898
rect -64477 -30198 -64473 -29902
rect -64473 -30198 -64177 -29902
rect -64177 -30198 -64173 -29902
rect -64477 -30202 -64173 -30198
rect -64137 -29902 -63513 -29898
rect -64137 -30198 -64133 -29902
rect -64133 -30198 -63517 -29902
rect -63517 -30198 -63513 -29902
rect -64137 -30202 -63513 -30198
rect -63477 -29902 -63173 -29898
rect -63477 -30198 -63473 -29902
rect -63473 -30198 -63177 -29902
rect -63177 -30198 -63173 -29902
rect -63477 -30202 -63173 -30198
rect -63137 -29902 -62513 -29898
rect -63137 -30198 -63133 -29902
rect -63133 -30198 -62517 -29902
rect -62517 -30198 -62513 -29902
rect -63137 -30202 -62513 -30198
rect -62477 -29902 -62173 -29898
rect -62477 -30198 -62473 -29902
rect -62473 -30198 -62177 -29902
rect -62177 -30198 -62173 -29902
rect -62477 -30202 -62173 -30198
rect -62137 -29902 -61513 -29898
rect -62137 -30198 -62133 -29902
rect -62133 -30198 -61517 -29902
rect -61517 -30198 -61513 -29902
rect -62137 -30202 -61513 -30198
rect -61477 -29902 -61173 -29898
rect -61477 -30198 -61473 -29902
rect -61473 -30198 -61177 -29902
rect -61177 -30198 -61173 -29902
rect -61477 -30202 -61173 -30198
rect -61137 -29902 -60513 -29898
rect -61137 -30198 -61133 -29902
rect -61133 -30198 -60517 -29902
rect -60517 -30198 -60513 -29902
rect -61137 -30202 -60513 -30198
rect -60477 -29902 -60173 -29898
rect -60477 -30198 -60473 -29902
rect -60473 -30198 -60177 -29902
rect -60177 -30198 -60173 -29902
rect -60477 -30202 -60173 -30198
rect -60137 -29902 -59513 -29898
rect -60137 -30198 -60133 -29902
rect -60133 -30198 -59517 -29902
rect -59517 -30198 -59513 -29902
rect -60137 -30202 -59513 -30198
rect -59477 -29902 -59173 -29898
rect -59477 -30198 -59473 -29902
rect -59473 -30198 -59177 -29902
rect -59177 -30198 -59173 -29902
rect -59477 -30202 -59173 -30198
rect -59137 -29902 -58513 -29898
rect -59137 -30198 -59133 -29902
rect -59133 -30198 -58517 -29902
rect -58517 -30198 -58513 -29902
rect -59137 -30202 -58513 -30198
rect -58477 -29902 -58173 -29898
rect -58477 -30198 -58473 -29902
rect -58473 -30198 -58177 -29902
rect -58177 -30198 -58173 -29902
rect -58477 -30202 -58173 -30198
rect -58137 -29902 -57513 -29898
rect -58137 -30198 -58133 -29902
rect -58133 -30198 -57517 -29902
rect -57517 -30198 -57513 -29902
rect -58137 -30202 -57513 -30198
rect -57477 -29902 -57173 -29898
rect -57477 -30198 -57473 -29902
rect -57473 -30198 -57177 -29902
rect -57177 -30198 -57173 -29902
rect -57477 -30202 -57173 -30198
rect -57137 -29902 -56513 -29898
rect -57137 -30198 -57133 -29902
rect -57133 -30198 -56517 -29902
rect -56517 -30198 -56513 -29902
rect -57137 -30202 -56513 -30198
rect -56477 -29902 -56173 -29898
rect -56477 -30198 -56473 -29902
rect -56473 -30198 -56177 -29902
rect -56177 -30198 -56173 -29902
rect -56477 -30202 -56173 -30198
rect -56137 -29902 -55513 -29898
rect -56137 -30198 -56133 -29902
rect -56133 -30198 -55517 -29902
rect -55517 -30198 -55513 -29902
rect -56137 -30202 -55513 -30198
rect -55477 -29902 -55173 -29898
rect -55477 -30198 -55473 -29902
rect -55473 -30198 -55177 -29902
rect -55177 -30198 -55173 -29902
rect -55477 -30202 -55173 -30198
rect -55137 -29902 -54513 -29898
rect -55137 -30198 -55133 -29902
rect -55133 -30198 -54517 -29902
rect -54517 -30198 -54513 -29902
rect -55137 -30202 -54513 -30198
rect -54477 -29902 -54173 -29898
rect -54477 -30198 -54473 -29902
rect -54473 -30198 -54177 -29902
rect -54177 -30198 -54173 -29902
rect -54477 -30202 -54173 -30198
rect -54137 -29902 -53513 -29898
rect -54137 -30198 -54133 -29902
rect -54133 -30198 -53517 -29902
rect -53517 -30198 -53513 -29902
rect -54137 -30202 -53513 -30198
rect -53477 -29902 -53173 -29898
rect -53477 -30198 -53473 -29902
rect -53473 -30198 -53177 -29902
rect -53177 -30198 -53173 -29902
rect -53477 -30202 -53173 -30198
rect -53137 -29902 -52513 -29898
rect -53137 -30198 -53133 -29902
rect -53133 -30198 -52517 -29902
rect -52517 -30198 -52513 -29902
rect -53137 -30202 -52513 -30198
rect -52477 -29902 -52173 -29898
rect -52477 -30198 -52473 -29902
rect -52473 -30198 -52177 -29902
rect -52177 -30198 -52173 -29902
rect -52477 -30202 -52173 -30198
rect -52137 -29902 -51513 -29898
rect -52137 -30198 -52133 -29902
rect -52133 -30198 -51517 -29902
rect -51517 -30198 -51513 -29902
rect -52137 -30202 -51513 -30198
rect -51477 -29902 -51173 -29898
rect -51477 -30198 -51473 -29902
rect -51473 -30198 -51177 -29902
rect -51177 -30198 -51173 -29902
rect -51477 -30202 -51173 -30198
rect -51137 -29902 -50513 -29898
rect -51137 -30198 -51133 -29902
rect -51133 -30198 -50517 -29902
rect -50517 -30198 -50513 -29902
rect -51137 -30202 -50513 -30198
rect -50477 -29902 -50173 -29898
rect -50477 -30198 -50473 -29902
rect -50473 -30198 -50177 -29902
rect -50177 -30198 -50173 -29902
rect -50477 -30202 -50173 -30198
rect -50137 -29902 -49513 -29898
rect -50137 -30198 -50133 -29902
rect -50133 -30198 -49517 -29902
rect -49517 -30198 -49513 -29902
rect -50137 -30202 -49513 -30198
rect -49477 -29902 -49173 -29898
rect -49477 -30198 -49473 -29902
rect -49473 -30198 -49177 -29902
rect -49177 -30198 -49173 -29902
rect -49477 -30202 -49173 -30198
rect -49137 -29902 -48833 -29898
rect -49137 -30198 -49133 -29902
rect -49133 -30198 -48837 -29902
rect -48837 -30198 -48833 -29902
rect -49137 -30202 -48833 -30198
rect 8283 -29902 8587 -29898
rect 8283 -30198 8287 -29902
rect 8287 -30198 8583 -29902
rect 8583 -30198 8587 -29902
rect 8283 -30202 8587 -30198
rect 8623 -29902 8927 -29898
rect 8623 -30198 8627 -29902
rect 8627 -30198 8923 -29902
rect 8923 -30198 8927 -29902
rect 8623 -30202 8927 -30198
rect 8963 -29902 9587 -29898
rect 8963 -30198 8967 -29902
rect 8967 -30198 9583 -29902
rect 9583 -30198 9587 -29902
rect 8963 -30202 9587 -30198
rect 9623 -29902 9927 -29898
rect 9623 -30198 9627 -29902
rect 9627 -30198 9923 -29902
rect 9923 -30198 9927 -29902
rect 9623 -30202 9927 -30198
rect 9963 -29902 10587 -29898
rect 9963 -30198 9967 -29902
rect 9967 -30198 10583 -29902
rect 10583 -30198 10587 -29902
rect 9963 -30202 10587 -30198
rect 10623 -29902 10927 -29898
rect 10623 -30198 10627 -29902
rect 10627 -30198 10923 -29902
rect 10923 -30198 10927 -29902
rect 10623 -30202 10927 -30198
rect 10963 -29902 11587 -29898
rect 10963 -30198 10967 -29902
rect 10967 -30198 11583 -29902
rect 11583 -30198 11587 -29902
rect 10963 -30202 11587 -30198
rect 11623 -29902 11927 -29898
rect 11623 -30198 11627 -29902
rect 11627 -30198 11923 -29902
rect 11923 -30198 11927 -29902
rect 11623 -30202 11927 -30198
rect 11963 -29902 12587 -29898
rect 11963 -30198 11967 -29902
rect 11967 -30198 12583 -29902
rect 12583 -30198 12587 -29902
rect 11963 -30202 12587 -30198
rect 12623 -29902 12927 -29898
rect 12623 -30198 12627 -29902
rect 12627 -30198 12923 -29902
rect 12923 -30198 12927 -29902
rect 12623 -30202 12927 -30198
rect 12963 -29902 13587 -29898
rect 12963 -30198 12967 -29902
rect 12967 -30198 13583 -29902
rect 13583 -30198 13587 -29902
rect 12963 -30202 13587 -30198
rect 13623 -29902 13927 -29898
rect 13623 -30198 13627 -29902
rect 13627 -30198 13923 -29902
rect 13923 -30198 13927 -29902
rect 13623 -30202 13927 -30198
rect 13963 -29902 14587 -29898
rect 13963 -30198 13967 -29902
rect 13967 -30198 14583 -29902
rect 14583 -30198 14587 -29902
rect 13963 -30202 14587 -30198
rect 14623 -29902 14927 -29898
rect 14623 -30198 14627 -29902
rect 14627 -30198 14923 -29902
rect 14923 -30198 14927 -29902
rect 14623 -30202 14927 -30198
rect 14963 -29902 15587 -29898
rect 14963 -30198 14967 -29902
rect 14967 -30198 15583 -29902
rect 15583 -30198 15587 -29902
rect 14963 -30202 15587 -30198
rect 15623 -29902 15927 -29898
rect 15623 -30198 15627 -29902
rect 15627 -30198 15923 -29902
rect 15923 -30198 15927 -29902
rect 15623 -30202 15927 -30198
rect 15963 -29902 16587 -29898
rect 15963 -30198 15967 -29902
rect 15967 -30198 16583 -29902
rect 16583 -30198 16587 -29902
rect 15963 -30202 16587 -30198
rect 16623 -29902 16927 -29898
rect 16623 -30198 16627 -29902
rect 16627 -30198 16923 -29902
rect 16923 -30198 16927 -29902
rect 16623 -30202 16927 -30198
rect 16963 -29902 17587 -29898
rect 16963 -30198 16967 -29902
rect 16967 -30198 17583 -29902
rect 17583 -30198 17587 -29902
rect 16963 -30202 17587 -30198
rect 17623 -29902 17927 -29898
rect 17623 -30198 17627 -29902
rect 17627 -30198 17923 -29902
rect 17923 -30198 17927 -29902
rect 17623 -30202 17927 -30198
rect 17963 -29902 18587 -29898
rect 17963 -30198 17967 -29902
rect 17967 -30198 18583 -29902
rect 18583 -30198 18587 -29902
rect 17963 -30202 18587 -30198
rect 18623 -29902 18927 -29898
rect 18623 -30198 18627 -29902
rect 18627 -30198 18923 -29902
rect 18923 -30198 18927 -29902
rect 18623 -30202 18927 -30198
rect 18963 -29902 19587 -29898
rect 18963 -30198 18967 -29902
rect 18967 -30198 19583 -29902
rect 19583 -30198 19587 -29902
rect 18963 -30202 19587 -30198
rect 19623 -29902 19927 -29898
rect 19623 -30198 19627 -29902
rect 19627 -30198 19923 -29902
rect 19923 -30198 19927 -29902
rect 19623 -30202 19927 -30198
rect 19963 -29902 20587 -29898
rect 19963 -30198 19967 -29902
rect 19967 -30198 20583 -29902
rect 20583 -30198 20587 -29902
rect 19963 -30202 20587 -30198
rect 20623 -29902 20927 -29898
rect 20623 -30198 20627 -29902
rect 20627 -30198 20923 -29902
rect 20923 -30198 20927 -29902
rect 20623 -30202 20927 -30198
rect 20963 -29902 21587 -29898
rect 20963 -30198 20967 -29902
rect 20967 -30198 21583 -29902
rect 21583 -30198 21587 -29902
rect 20963 -30202 21587 -30198
rect 21623 -29902 21927 -29898
rect 21623 -30198 21627 -29902
rect 21627 -30198 21923 -29902
rect 21923 -30198 21927 -29902
rect 21623 -30202 21927 -30198
rect 21963 -29902 22587 -29898
rect 21963 -30198 21967 -29902
rect 21967 -30198 22583 -29902
rect 22583 -30198 22587 -29902
rect 21963 -30202 22587 -30198
rect 22623 -29902 22927 -29898
rect 22623 -30198 22627 -29902
rect 22627 -30198 22923 -29902
rect 22923 -30198 22927 -29902
rect 22623 -30202 22927 -30198
rect 22963 -29902 23587 -29898
rect 22963 -30198 22967 -29902
rect 22967 -30198 23583 -29902
rect 23583 -30198 23587 -29902
rect 22963 -30202 23587 -30198
rect 23623 -29902 23927 -29898
rect 23623 -30198 23627 -29902
rect 23627 -30198 23923 -29902
rect 23923 -30198 23927 -29902
rect 23623 -30202 23927 -30198
rect 23963 -29902 24587 -29898
rect 23963 -30198 23967 -29902
rect 23967 -30198 24583 -29902
rect 24583 -30198 24587 -29902
rect 23963 -30202 24587 -30198
rect 24623 -29902 24927 -29898
rect 24623 -30198 24627 -29902
rect 24627 -30198 24923 -29902
rect 24923 -30198 24927 -29902
rect 24623 -30202 24927 -30198
rect 24963 -29902 25587 -29898
rect 24963 -30198 24967 -29902
rect 24967 -30198 25583 -29902
rect 25583 -30198 25587 -29902
rect 24963 -30202 25587 -30198
rect 25623 -29902 25927 -29898
rect 25623 -30198 25627 -29902
rect 25627 -30198 25923 -29902
rect 25923 -30198 25927 -29902
rect 25623 -30202 25927 -30198
rect 25963 -29902 26587 -29898
rect 25963 -30198 25967 -29902
rect 25967 -30198 26583 -29902
rect 26583 -30198 26587 -29902
rect 25963 -30202 26587 -30198
rect 26623 -29902 26927 -29898
rect 26623 -30198 26627 -29902
rect 26627 -30198 26923 -29902
rect 26923 -30198 26927 -29902
rect 26623 -30202 26927 -30198
rect 26963 -29902 27587 -29898
rect 26963 -30198 26967 -29902
rect 26967 -30198 27583 -29902
rect 27583 -30198 27587 -29902
rect 26963 -30202 27587 -30198
rect 27623 -29902 27927 -29898
rect 27623 -30198 27627 -29902
rect 27627 -30198 27923 -29902
rect 27923 -30198 27927 -29902
rect 27623 -30202 27927 -30198
rect 27963 -29902 28587 -29898
rect 27963 -30198 27967 -29902
rect 27967 -30198 28583 -29902
rect 28583 -30198 28587 -29902
rect 27963 -30202 28587 -30198
rect 28623 -29902 28927 -29898
rect 28623 -30198 28627 -29902
rect 28627 -30198 28923 -29902
rect 28923 -30198 28927 -29902
rect 28623 -30202 28927 -30198
rect 28963 -29902 29587 -29898
rect 28963 -30198 28967 -29902
rect 28967 -30198 29583 -29902
rect 29583 -30198 29587 -29902
rect 28963 -30202 29587 -30198
rect 29623 -29902 29927 -29898
rect 29623 -30198 29627 -29902
rect 29627 -30198 29923 -29902
rect 29923 -30198 29927 -29902
rect 29623 -30202 29927 -30198
rect 29963 -29902 30587 -29898
rect 29963 -30198 29967 -29902
rect 29967 -30198 30583 -29902
rect 30583 -30198 30587 -29902
rect 29963 -30202 30587 -30198
rect 30623 -29902 30927 -29898
rect 30623 -30198 30627 -29902
rect 30627 -30198 30923 -29902
rect 30923 -30198 30927 -29902
rect 30623 -30202 30927 -30198
rect 30963 -29902 31587 -29898
rect 30963 -30198 30967 -29902
rect 30967 -30198 31583 -29902
rect 31583 -30198 31587 -29902
rect 30963 -30202 31587 -30198
rect 31623 -29902 31927 -29898
rect 31623 -30198 31627 -29902
rect 31627 -30198 31923 -29902
rect 31923 -30198 31927 -29902
rect 31623 -30202 31927 -30198
rect 31963 -29902 32587 -29898
rect 31963 -30198 31967 -29902
rect 31967 -30198 32583 -29902
rect 32583 -30198 32587 -29902
rect 31963 -30202 32587 -30198
rect 32623 -29902 32927 -29898
rect 32623 -30198 32627 -29902
rect 32627 -30198 32923 -29902
rect 32923 -30198 32927 -29902
rect 32623 -30202 32927 -30198
rect 32963 -29902 33587 -29898
rect 32963 -30198 32967 -29902
rect 32967 -30198 33583 -29902
rect 33583 -30198 33587 -29902
rect 32963 -30202 33587 -30198
rect 33623 -29902 33927 -29898
rect 33623 -30198 33627 -29902
rect 33627 -30198 33923 -29902
rect 33923 -30198 33927 -29902
rect 33623 -30202 33927 -30198
rect 33963 -29902 34267 -29898
rect 33963 -30198 33967 -29902
rect 33967 -30198 34263 -29902
rect 34263 -30198 34267 -29902
rect 33963 -30202 34267 -30198
rect -74477 -30242 -74173 -30238
rect -74477 -30858 -74473 -30242
rect -74473 -30858 -74177 -30242
rect -74177 -30858 -74173 -30242
rect -74477 -30862 -74173 -30858
rect -73477 -30242 -73173 -30238
rect -73477 -30858 -73473 -30242
rect -73473 -30858 -73177 -30242
rect -73177 -30858 -73173 -30242
rect -73477 -30862 -73173 -30858
rect -72477 -30242 -72173 -30238
rect -72477 -30858 -72473 -30242
rect -72473 -30858 -72177 -30242
rect -72177 -30858 -72173 -30242
rect -72477 -30862 -72173 -30858
rect -71477 -30242 -71173 -30238
rect -71477 -30858 -71473 -30242
rect -71473 -30858 -71177 -30242
rect -71177 -30858 -71173 -30242
rect -71477 -30862 -71173 -30858
rect -70477 -30242 -70173 -30238
rect -70477 -30858 -70473 -30242
rect -70473 -30858 -70177 -30242
rect -70177 -30858 -70173 -30242
rect -70477 -30862 -70173 -30858
rect -69477 -30242 -69173 -30238
rect -69477 -30858 -69473 -30242
rect -69473 -30858 -69177 -30242
rect -69177 -30858 -69173 -30242
rect -69477 -30862 -69173 -30858
rect -68477 -30242 -68173 -30238
rect -68477 -30858 -68473 -30242
rect -68473 -30858 -68177 -30242
rect -68177 -30858 -68173 -30242
rect -68477 -30862 -68173 -30858
rect -67477 -30242 -67173 -30238
rect -67477 -30858 -67473 -30242
rect -67473 -30858 -67177 -30242
rect -67177 -30858 -67173 -30242
rect -67477 -30862 -67173 -30858
rect -66477 -30242 -66173 -30238
rect -66477 -30858 -66473 -30242
rect -66473 -30858 -66177 -30242
rect -66177 -30858 -66173 -30242
rect -66477 -30862 -66173 -30858
rect -65477 -30242 -65173 -30238
rect -65477 -30858 -65473 -30242
rect -65473 -30858 -65177 -30242
rect -65177 -30858 -65173 -30242
rect -65477 -30862 -65173 -30858
rect -64477 -30242 -64173 -30238
rect -64477 -30858 -64473 -30242
rect -64473 -30858 -64177 -30242
rect -64177 -30858 -64173 -30242
rect -64477 -30862 -64173 -30858
rect -63477 -30242 -63173 -30238
rect -63477 -30858 -63473 -30242
rect -63473 -30858 -63177 -30242
rect -63177 -30858 -63173 -30242
rect -63477 -30862 -63173 -30858
rect -62477 -30242 -62173 -30238
rect -62477 -30858 -62473 -30242
rect -62473 -30858 -62177 -30242
rect -62177 -30858 -62173 -30242
rect -62477 -30862 -62173 -30858
rect -61477 -30242 -61173 -30238
rect -61477 -30858 -61473 -30242
rect -61473 -30858 -61177 -30242
rect -61177 -30858 -61173 -30242
rect -61477 -30862 -61173 -30858
rect -60477 -30242 -60173 -30238
rect -60477 -30858 -60473 -30242
rect -60473 -30858 -60177 -30242
rect -60177 -30858 -60173 -30242
rect -60477 -30862 -60173 -30858
rect -59477 -30242 -59173 -30238
rect -59477 -30858 -59473 -30242
rect -59473 -30858 -59177 -30242
rect -59177 -30858 -59173 -30242
rect -59477 -30862 -59173 -30858
rect -58477 -30242 -58173 -30238
rect -58477 -30858 -58473 -30242
rect -58473 -30858 -58177 -30242
rect -58177 -30858 -58173 -30242
rect -58477 -30862 -58173 -30858
rect -57477 -30242 -57173 -30238
rect -57477 -30858 -57473 -30242
rect -57473 -30858 -57177 -30242
rect -57177 -30858 -57173 -30242
rect -57477 -30862 -57173 -30858
rect -56477 -30242 -56173 -30238
rect -56477 -30858 -56473 -30242
rect -56473 -30858 -56177 -30242
rect -56177 -30858 -56173 -30242
rect -56477 -30862 -56173 -30858
rect -55477 -30242 -55173 -30238
rect -55477 -30858 -55473 -30242
rect -55473 -30858 -55177 -30242
rect -55177 -30858 -55173 -30242
rect -55477 -30862 -55173 -30858
rect -54477 -30242 -54173 -30238
rect -54477 -30858 -54473 -30242
rect -54473 -30858 -54177 -30242
rect -54177 -30858 -54173 -30242
rect -54477 -30862 -54173 -30858
rect -53477 -30242 -53173 -30238
rect -53477 -30858 -53473 -30242
rect -53473 -30858 -53177 -30242
rect -53177 -30858 -53173 -30242
rect -53477 -30862 -53173 -30858
rect -52477 -30242 -52173 -30238
rect -52477 -30858 -52473 -30242
rect -52473 -30858 -52177 -30242
rect -52177 -30858 -52173 -30242
rect -52477 -30862 -52173 -30858
rect -51477 -30242 -51173 -30238
rect -51477 -30858 -51473 -30242
rect -51473 -30858 -51177 -30242
rect -51177 -30858 -51173 -30242
rect -51477 -30862 -51173 -30858
rect -50477 -30242 -50173 -30238
rect -50477 -30858 -50473 -30242
rect -50473 -30858 -50177 -30242
rect -50177 -30858 -50173 -30242
rect -50477 -30862 -50173 -30858
rect -49477 -30242 -49173 -30238
rect -49477 -30858 -49473 -30242
rect -49473 -30858 -49177 -30242
rect -49177 -30858 -49173 -30242
rect -49477 -30862 -49173 -30858
rect 8623 -30242 8927 -30238
rect 8623 -30858 8627 -30242
rect 8627 -30858 8923 -30242
rect 8923 -30858 8927 -30242
rect 8623 -30862 8927 -30858
rect 9623 -30242 9927 -30238
rect 9623 -30858 9627 -30242
rect 9627 -30858 9923 -30242
rect 9923 -30858 9927 -30242
rect 9623 -30862 9927 -30858
rect 10623 -30242 10927 -30238
rect 10623 -30858 10627 -30242
rect 10627 -30858 10923 -30242
rect 10923 -30858 10927 -30242
rect 10623 -30862 10927 -30858
rect 11623 -30242 11927 -30238
rect 11623 -30858 11627 -30242
rect 11627 -30858 11923 -30242
rect 11923 -30858 11927 -30242
rect 11623 -30862 11927 -30858
rect 12623 -30242 12927 -30238
rect 12623 -30858 12627 -30242
rect 12627 -30858 12923 -30242
rect 12923 -30858 12927 -30242
rect 12623 -30862 12927 -30858
rect 13623 -30242 13927 -30238
rect 13623 -30858 13627 -30242
rect 13627 -30858 13923 -30242
rect 13923 -30858 13927 -30242
rect 13623 -30862 13927 -30858
rect 14623 -30242 14927 -30238
rect 14623 -30858 14627 -30242
rect 14627 -30858 14923 -30242
rect 14923 -30858 14927 -30242
rect 14623 -30862 14927 -30858
rect 15623 -30242 15927 -30238
rect 15623 -30858 15627 -30242
rect 15627 -30858 15923 -30242
rect 15923 -30858 15927 -30242
rect 15623 -30862 15927 -30858
rect 16623 -30242 16927 -30238
rect 16623 -30858 16627 -30242
rect 16627 -30858 16923 -30242
rect 16923 -30858 16927 -30242
rect 16623 -30862 16927 -30858
rect 17623 -30242 17927 -30238
rect 17623 -30858 17627 -30242
rect 17627 -30858 17923 -30242
rect 17923 -30858 17927 -30242
rect 17623 -30862 17927 -30858
rect 18623 -30242 18927 -30238
rect 18623 -30858 18627 -30242
rect 18627 -30858 18923 -30242
rect 18923 -30858 18927 -30242
rect 18623 -30862 18927 -30858
rect 19623 -30242 19927 -30238
rect 19623 -30858 19627 -30242
rect 19627 -30858 19923 -30242
rect 19923 -30858 19927 -30242
rect 19623 -30862 19927 -30858
rect 20623 -30242 20927 -30238
rect 20623 -30858 20627 -30242
rect 20627 -30858 20923 -30242
rect 20923 -30858 20927 -30242
rect 20623 -30862 20927 -30858
rect 21623 -30242 21927 -30238
rect 21623 -30858 21627 -30242
rect 21627 -30858 21923 -30242
rect 21923 -30858 21927 -30242
rect 21623 -30862 21927 -30858
rect 22623 -30242 22927 -30238
rect 22623 -30858 22627 -30242
rect 22627 -30858 22923 -30242
rect 22923 -30858 22927 -30242
rect 22623 -30862 22927 -30858
rect 23623 -30242 23927 -30238
rect 23623 -30858 23627 -30242
rect 23627 -30858 23923 -30242
rect 23923 -30858 23927 -30242
rect 23623 -30862 23927 -30858
rect 24623 -30242 24927 -30238
rect 24623 -30858 24627 -30242
rect 24627 -30858 24923 -30242
rect 24923 -30858 24927 -30242
rect 24623 -30862 24927 -30858
rect 25623 -30242 25927 -30238
rect 25623 -30858 25627 -30242
rect 25627 -30858 25923 -30242
rect 25923 -30858 25927 -30242
rect 25623 -30862 25927 -30858
rect 26623 -30242 26927 -30238
rect 26623 -30858 26627 -30242
rect 26627 -30858 26923 -30242
rect 26923 -30858 26927 -30242
rect 26623 -30862 26927 -30858
rect 27623 -30242 27927 -30238
rect 27623 -30858 27627 -30242
rect 27627 -30858 27923 -30242
rect 27923 -30858 27927 -30242
rect 27623 -30862 27927 -30858
rect 28623 -30242 28927 -30238
rect 28623 -30858 28627 -30242
rect 28627 -30858 28923 -30242
rect 28923 -30858 28927 -30242
rect 28623 -30862 28927 -30858
rect 29623 -30242 29927 -30238
rect 29623 -30858 29627 -30242
rect 29627 -30858 29923 -30242
rect 29923 -30858 29927 -30242
rect 29623 -30862 29927 -30858
rect 30623 -30242 30927 -30238
rect 30623 -30858 30627 -30242
rect 30627 -30858 30923 -30242
rect 30923 -30858 30927 -30242
rect 30623 -30862 30927 -30858
rect 31623 -30242 31927 -30238
rect 31623 -30858 31627 -30242
rect 31627 -30858 31923 -30242
rect 31923 -30858 31927 -30242
rect 31623 -30862 31927 -30858
rect 32623 -30242 32927 -30238
rect 32623 -30858 32627 -30242
rect 32627 -30858 32923 -30242
rect 32923 -30858 32927 -30242
rect 32623 -30862 32927 -30858
rect 33623 -30242 33927 -30238
rect 33623 -30858 33627 -30242
rect 33627 -30858 33923 -30242
rect 33923 -30858 33927 -30242
rect 33623 -30862 33927 -30858
rect -74817 -30902 -74513 -30898
rect -74817 -31198 -74813 -30902
rect -74813 -31198 -74517 -30902
rect -74517 -31198 -74513 -30902
rect -74817 -31202 -74513 -31198
rect -74477 -30902 -74173 -30898
rect -74477 -31198 -74473 -30902
rect -74473 -31198 -74177 -30902
rect -74177 -31198 -74173 -30902
rect -74477 -31202 -74173 -31198
rect -74137 -30902 -73513 -30898
rect -74137 -31198 -74133 -30902
rect -74133 -31198 -73517 -30902
rect -73517 -31198 -73513 -30902
rect -74137 -31202 -73513 -31198
rect -73477 -30902 -73173 -30898
rect -73477 -31198 -73473 -30902
rect -73473 -31198 -73177 -30902
rect -73177 -31198 -73173 -30902
rect -73477 -31202 -73173 -31198
rect -73137 -30902 -72513 -30898
rect -73137 -31198 -73133 -30902
rect -73133 -31198 -72517 -30902
rect -72517 -31198 -72513 -30902
rect -73137 -31202 -72513 -31198
rect -72477 -30902 -72173 -30898
rect -72477 -31198 -72473 -30902
rect -72473 -31198 -72177 -30902
rect -72177 -31198 -72173 -30902
rect -72477 -31202 -72173 -31198
rect -72137 -30902 -71513 -30898
rect -72137 -31198 -72133 -30902
rect -72133 -31198 -71517 -30902
rect -71517 -31198 -71513 -30902
rect -72137 -31202 -71513 -31198
rect -71477 -30902 -71173 -30898
rect -71477 -31198 -71473 -30902
rect -71473 -31198 -71177 -30902
rect -71177 -31198 -71173 -30902
rect -71477 -31202 -71173 -31198
rect -71137 -30902 -70513 -30898
rect -71137 -31198 -71133 -30902
rect -71133 -31198 -70517 -30902
rect -70517 -31198 -70513 -30902
rect -71137 -31202 -70513 -31198
rect -70477 -30902 -70173 -30898
rect -70477 -31198 -70473 -30902
rect -70473 -31198 -70177 -30902
rect -70177 -31198 -70173 -30902
rect -70477 -31202 -70173 -31198
rect -70137 -30902 -69513 -30898
rect -70137 -31198 -70133 -30902
rect -70133 -31198 -69517 -30902
rect -69517 -31198 -69513 -30902
rect -70137 -31202 -69513 -31198
rect -69477 -30902 -69173 -30898
rect -69477 -31198 -69473 -30902
rect -69473 -31198 -69177 -30902
rect -69177 -31198 -69173 -30902
rect -69477 -31202 -69173 -31198
rect -69137 -30902 -68513 -30898
rect -69137 -31198 -69133 -30902
rect -69133 -31198 -68517 -30902
rect -68517 -31198 -68513 -30902
rect -69137 -31202 -68513 -31198
rect -68477 -30902 -68173 -30898
rect -68477 -31198 -68473 -30902
rect -68473 -31198 -68177 -30902
rect -68177 -31198 -68173 -30902
rect -68477 -31202 -68173 -31198
rect -68137 -30902 -67513 -30898
rect -68137 -31198 -68133 -30902
rect -68133 -31198 -67517 -30902
rect -67517 -31198 -67513 -30902
rect -68137 -31202 -67513 -31198
rect -67477 -30902 -67173 -30898
rect -67477 -31198 -67473 -30902
rect -67473 -31198 -67177 -30902
rect -67177 -31198 -67173 -30902
rect -67477 -31202 -67173 -31198
rect -67137 -30902 -66513 -30898
rect -67137 -31198 -67133 -30902
rect -67133 -31198 -66517 -30902
rect -66517 -31198 -66513 -30902
rect -67137 -31202 -66513 -31198
rect -66477 -30902 -66173 -30898
rect -66477 -31198 -66473 -30902
rect -66473 -31198 -66177 -30902
rect -66177 -31198 -66173 -30902
rect -66477 -31202 -66173 -31198
rect -66137 -30902 -65513 -30898
rect -66137 -31198 -66133 -30902
rect -66133 -31198 -65517 -30902
rect -65517 -31198 -65513 -30902
rect -66137 -31202 -65513 -31198
rect -65477 -30902 -65173 -30898
rect -65477 -31198 -65473 -30902
rect -65473 -31198 -65177 -30902
rect -65177 -31198 -65173 -30902
rect -65477 -31202 -65173 -31198
rect -65137 -30902 -64513 -30898
rect -65137 -31198 -65133 -30902
rect -65133 -31198 -64517 -30902
rect -64517 -31198 -64513 -30902
rect -65137 -31202 -64513 -31198
rect -64477 -30902 -64173 -30898
rect -64477 -31198 -64473 -30902
rect -64473 -31198 -64177 -30902
rect -64177 -31198 -64173 -30902
rect -64477 -31202 -64173 -31198
rect -64137 -30902 -63513 -30898
rect -64137 -31198 -64133 -30902
rect -64133 -31198 -63517 -30902
rect -63517 -31198 -63513 -30902
rect -64137 -31202 -63513 -31198
rect -63477 -30902 -63173 -30898
rect -63477 -31198 -63473 -30902
rect -63473 -31198 -63177 -30902
rect -63177 -31198 -63173 -30902
rect -63477 -31202 -63173 -31198
rect -63137 -30902 -62513 -30898
rect -63137 -31198 -63133 -30902
rect -63133 -31198 -62517 -30902
rect -62517 -31198 -62513 -30902
rect -63137 -31202 -62513 -31198
rect -62477 -30902 -62173 -30898
rect -62477 -31198 -62473 -30902
rect -62473 -31198 -62177 -30902
rect -62177 -31198 -62173 -30902
rect -62477 -31202 -62173 -31198
rect -62137 -30902 -61513 -30898
rect -62137 -31198 -62133 -30902
rect -62133 -31198 -61517 -30902
rect -61517 -31198 -61513 -30902
rect -62137 -31202 -61513 -31198
rect -61477 -30902 -61173 -30898
rect -61477 -31198 -61473 -30902
rect -61473 -31198 -61177 -30902
rect -61177 -31198 -61173 -30902
rect -61477 -31202 -61173 -31198
rect -61137 -30902 -60513 -30898
rect -61137 -31198 -61133 -30902
rect -61133 -31198 -60517 -30902
rect -60517 -31198 -60513 -30902
rect -61137 -31202 -60513 -31198
rect -60477 -30902 -60173 -30898
rect -60477 -31198 -60473 -30902
rect -60473 -31198 -60177 -30902
rect -60177 -31198 -60173 -30902
rect -60477 -31202 -60173 -31198
rect -60137 -30902 -59513 -30898
rect -60137 -31198 -60133 -30902
rect -60133 -31198 -59517 -30902
rect -59517 -31198 -59513 -30902
rect -60137 -31202 -59513 -31198
rect -59477 -30902 -59173 -30898
rect -59477 -31198 -59473 -30902
rect -59473 -31198 -59177 -30902
rect -59177 -31198 -59173 -30902
rect -59477 -31202 -59173 -31198
rect -59137 -30902 -58513 -30898
rect -59137 -31198 -59133 -30902
rect -59133 -31198 -58517 -30902
rect -58517 -31198 -58513 -30902
rect -59137 -31202 -58513 -31198
rect -58477 -30902 -58173 -30898
rect -58477 -31198 -58473 -30902
rect -58473 -31198 -58177 -30902
rect -58177 -31198 -58173 -30902
rect -58477 -31202 -58173 -31198
rect -58137 -30902 -57513 -30898
rect -58137 -31198 -58133 -30902
rect -58133 -31198 -57517 -30902
rect -57517 -31198 -57513 -30902
rect -58137 -31202 -57513 -31198
rect -57477 -30902 -57173 -30898
rect -57477 -31198 -57473 -30902
rect -57473 -31198 -57177 -30902
rect -57177 -31198 -57173 -30902
rect -57477 -31202 -57173 -31198
rect -57137 -30902 -56513 -30898
rect -57137 -31198 -57133 -30902
rect -57133 -31198 -56517 -30902
rect -56517 -31198 -56513 -30902
rect -57137 -31202 -56513 -31198
rect -56477 -30902 -56173 -30898
rect -56477 -31198 -56473 -30902
rect -56473 -31198 -56177 -30902
rect -56177 -31198 -56173 -30902
rect -56477 -31202 -56173 -31198
rect -56137 -30902 -55513 -30898
rect -56137 -31198 -56133 -30902
rect -56133 -31198 -55517 -30902
rect -55517 -31198 -55513 -30902
rect -56137 -31202 -55513 -31198
rect -55477 -30902 -55173 -30898
rect -55477 -31198 -55473 -30902
rect -55473 -31198 -55177 -30902
rect -55177 -31198 -55173 -30902
rect -55477 -31202 -55173 -31198
rect -55137 -30902 -54513 -30898
rect -55137 -31198 -55133 -30902
rect -55133 -31198 -54517 -30902
rect -54517 -31198 -54513 -30902
rect -55137 -31202 -54513 -31198
rect -54477 -30902 -54173 -30898
rect -54477 -31198 -54473 -30902
rect -54473 -31198 -54177 -30902
rect -54177 -31198 -54173 -30902
rect -54477 -31202 -54173 -31198
rect -54137 -30902 -53513 -30898
rect -54137 -31198 -54133 -30902
rect -54133 -31198 -53517 -30902
rect -53517 -31198 -53513 -30902
rect -54137 -31202 -53513 -31198
rect -53477 -30902 -53173 -30898
rect -53477 -31198 -53473 -30902
rect -53473 -31198 -53177 -30902
rect -53177 -31198 -53173 -30902
rect -53477 -31202 -53173 -31198
rect -53137 -30902 -52513 -30898
rect -53137 -31198 -53133 -30902
rect -53133 -31198 -52517 -30902
rect -52517 -31198 -52513 -30902
rect -53137 -31202 -52513 -31198
rect -52477 -30902 -52173 -30898
rect -52477 -31198 -52473 -30902
rect -52473 -31198 -52177 -30902
rect -52177 -31198 -52173 -30902
rect -52477 -31202 -52173 -31198
rect -52137 -30902 -51513 -30898
rect -52137 -31198 -52133 -30902
rect -52133 -31198 -51517 -30902
rect -51517 -31198 -51513 -30902
rect -52137 -31202 -51513 -31198
rect -51477 -30902 -51173 -30898
rect -51477 -31198 -51473 -30902
rect -51473 -31198 -51177 -30902
rect -51177 -31198 -51173 -30902
rect -51477 -31202 -51173 -31198
rect -51137 -30902 -50513 -30898
rect -51137 -31198 -51133 -30902
rect -51133 -31198 -50517 -30902
rect -50517 -31198 -50513 -30902
rect -51137 -31202 -50513 -31198
rect -50477 -30902 -50173 -30898
rect -50477 -31198 -50473 -30902
rect -50473 -31198 -50177 -30902
rect -50177 -31198 -50173 -30902
rect -50477 -31202 -50173 -31198
rect -50137 -30902 -49513 -30898
rect -50137 -31198 -50133 -30902
rect -50133 -31198 -49517 -30902
rect -49517 -31198 -49513 -30902
rect -50137 -31202 -49513 -31198
rect -49477 -30902 -49173 -30898
rect -49477 -31198 -49473 -30902
rect -49473 -31198 -49177 -30902
rect -49177 -31198 -49173 -30902
rect -49477 -31202 -49173 -31198
rect -49137 -30902 -48833 -30898
rect -49137 -31198 -49133 -30902
rect -49133 -31198 -48837 -30902
rect -48837 -31198 -48833 -30902
rect -49137 -31202 -48833 -31198
rect 8283 -30902 8587 -30898
rect 8283 -31198 8287 -30902
rect 8287 -31198 8583 -30902
rect 8583 -31198 8587 -30902
rect 8283 -31202 8587 -31198
rect 8623 -30902 8927 -30898
rect 8623 -31198 8627 -30902
rect 8627 -31198 8923 -30902
rect 8923 -31198 8927 -30902
rect 8623 -31202 8927 -31198
rect 8963 -30902 9587 -30898
rect 8963 -31198 8967 -30902
rect 8967 -31198 9583 -30902
rect 9583 -31198 9587 -30902
rect 8963 -31202 9587 -31198
rect 9623 -30902 9927 -30898
rect 9623 -31198 9627 -30902
rect 9627 -31198 9923 -30902
rect 9923 -31198 9927 -30902
rect 9623 -31202 9927 -31198
rect 9963 -30902 10587 -30898
rect 9963 -31198 9967 -30902
rect 9967 -31198 10583 -30902
rect 10583 -31198 10587 -30902
rect 9963 -31202 10587 -31198
rect 10623 -30902 10927 -30898
rect 10623 -31198 10627 -30902
rect 10627 -31198 10923 -30902
rect 10923 -31198 10927 -30902
rect 10623 -31202 10927 -31198
rect 10963 -30902 11587 -30898
rect 10963 -31198 10967 -30902
rect 10967 -31198 11583 -30902
rect 11583 -31198 11587 -30902
rect 10963 -31202 11587 -31198
rect 11623 -30902 11927 -30898
rect 11623 -31198 11627 -30902
rect 11627 -31198 11923 -30902
rect 11923 -31198 11927 -30902
rect 11623 -31202 11927 -31198
rect 11963 -30902 12587 -30898
rect 11963 -31198 11967 -30902
rect 11967 -31198 12583 -30902
rect 12583 -31198 12587 -30902
rect 11963 -31202 12587 -31198
rect 12623 -30902 12927 -30898
rect 12623 -31198 12627 -30902
rect 12627 -31198 12923 -30902
rect 12923 -31198 12927 -30902
rect 12623 -31202 12927 -31198
rect 12963 -30902 13587 -30898
rect 12963 -31198 12967 -30902
rect 12967 -31198 13583 -30902
rect 13583 -31198 13587 -30902
rect 12963 -31202 13587 -31198
rect 13623 -30902 13927 -30898
rect 13623 -31198 13627 -30902
rect 13627 -31198 13923 -30902
rect 13923 -31198 13927 -30902
rect 13623 -31202 13927 -31198
rect 13963 -30902 14587 -30898
rect 13963 -31198 13967 -30902
rect 13967 -31198 14583 -30902
rect 14583 -31198 14587 -30902
rect 13963 -31202 14587 -31198
rect 14623 -30902 14927 -30898
rect 14623 -31198 14627 -30902
rect 14627 -31198 14923 -30902
rect 14923 -31198 14927 -30902
rect 14623 -31202 14927 -31198
rect 14963 -30902 15587 -30898
rect 14963 -31198 14967 -30902
rect 14967 -31198 15583 -30902
rect 15583 -31198 15587 -30902
rect 14963 -31202 15587 -31198
rect 15623 -30902 15927 -30898
rect 15623 -31198 15627 -30902
rect 15627 -31198 15923 -30902
rect 15923 -31198 15927 -30902
rect 15623 -31202 15927 -31198
rect 15963 -30902 16587 -30898
rect 15963 -31198 15967 -30902
rect 15967 -31198 16583 -30902
rect 16583 -31198 16587 -30902
rect 15963 -31202 16587 -31198
rect 16623 -30902 16927 -30898
rect 16623 -31198 16627 -30902
rect 16627 -31198 16923 -30902
rect 16923 -31198 16927 -30902
rect 16623 -31202 16927 -31198
rect 16963 -30902 17587 -30898
rect 16963 -31198 16967 -30902
rect 16967 -31198 17583 -30902
rect 17583 -31198 17587 -30902
rect 16963 -31202 17587 -31198
rect 17623 -30902 17927 -30898
rect 17623 -31198 17627 -30902
rect 17627 -31198 17923 -30902
rect 17923 -31198 17927 -30902
rect 17623 -31202 17927 -31198
rect 17963 -30902 18587 -30898
rect 17963 -31198 17967 -30902
rect 17967 -31198 18583 -30902
rect 18583 -31198 18587 -30902
rect 17963 -31202 18587 -31198
rect 18623 -30902 18927 -30898
rect 18623 -31198 18627 -30902
rect 18627 -31198 18923 -30902
rect 18923 -31198 18927 -30902
rect 18623 -31202 18927 -31198
rect 18963 -30902 19587 -30898
rect 18963 -31198 18967 -30902
rect 18967 -31198 19583 -30902
rect 19583 -31198 19587 -30902
rect 18963 -31202 19587 -31198
rect 19623 -30902 19927 -30898
rect 19623 -31198 19627 -30902
rect 19627 -31198 19923 -30902
rect 19923 -31198 19927 -30902
rect 19623 -31202 19927 -31198
rect 19963 -30902 20587 -30898
rect 19963 -31198 19967 -30902
rect 19967 -31198 20583 -30902
rect 20583 -31198 20587 -30902
rect 19963 -31202 20587 -31198
rect 20623 -30902 20927 -30898
rect 20623 -31198 20627 -30902
rect 20627 -31198 20923 -30902
rect 20923 -31198 20927 -30902
rect 20623 -31202 20927 -31198
rect 20963 -30902 21587 -30898
rect 20963 -31198 20967 -30902
rect 20967 -31198 21583 -30902
rect 21583 -31198 21587 -30902
rect 20963 -31202 21587 -31198
rect 21623 -30902 21927 -30898
rect 21623 -31198 21627 -30902
rect 21627 -31198 21923 -30902
rect 21923 -31198 21927 -30902
rect 21623 -31202 21927 -31198
rect 21963 -30902 22587 -30898
rect 21963 -31198 21967 -30902
rect 21967 -31198 22583 -30902
rect 22583 -31198 22587 -30902
rect 21963 -31202 22587 -31198
rect 22623 -30902 22927 -30898
rect 22623 -31198 22627 -30902
rect 22627 -31198 22923 -30902
rect 22923 -31198 22927 -30902
rect 22623 -31202 22927 -31198
rect 22963 -30902 23587 -30898
rect 22963 -31198 22967 -30902
rect 22967 -31198 23583 -30902
rect 23583 -31198 23587 -30902
rect 22963 -31202 23587 -31198
rect 23623 -30902 23927 -30898
rect 23623 -31198 23627 -30902
rect 23627 -31198 23923 -30902
rect 23923 -31198 23927 -30902
rect 23623 -31202 23927 -31198
rect 23963 -30902 24587 -30898
rect 23963 -31198 23967 -30902
rect 23967 -31198 24583 -30902
rect 24583 -31198 24587 -30902
rect 23963 -31202 24587 -31198
rect 24623 -30902 24927 -30898
rect 24623 -31198 24627 -30902
rect 24627 -31198 24923 -30902
rect 24923 -31198 24927 -30902
rect 24623 -31202 24927 -31198
rect 24963 -30902 25587 -30898
rect 24963 -31198 24967 -30902
rect 24967 -31198 25583 -30902
rect 25583 -31198 25587 -30902
rect 24963 -31202 25587 -31198
rect 25623 -30902 25927 -30898
rect 25623 -31198 25627 -30902
rect 25627 -31198 25923 -30902
rect 25923 -31198 25927 -30902
rect 25623 -31202 25927 -31198
rect 25963 -30902 26587 -30898
rect 25963 -31198 25967 -30902
rect 25967 -31198 26583 -30902
rect 26583 -31198 26587 -30902
rect 25963 -31202 26587 -31198
rect 26623 -30902 26927 -30898
rect 26623 -31198 26627 -30902
rect 26627 -31198 26923 -30902
rect 26923 -31198 26927 -30902
rect 26623 -31202 26927 -31198
rect 26963 -30902 27587 -30898
rect 26963 -31198 26967 -30902
rect 26967 -31198 27583 -30902
rect 27583 -31198 27587 -30902
rect 26963 -31202 27587 -31198
rect 27623 -30902 27927 -30898
rect 27623 -31198 27627 -30902
rect 27627 -31198 27923 -30902
rect 27923 -31198 27927 -30902
rect 27623 -31202 27927 -31198
rect 27963 -30902 28587 -30898
rect 27963 -31198 27967 -30902
rect 27967 -31198 28583 -30902
rect 28583 -31198 28587 -30902
rect 27963 -31202 28587 -31198
rect 28623 -30902 28927 -30898
rect 28623 -31198 28627 -30902
rect 28627 -31198 28923 -30902
rect 28923 -31198 28927 -30902
rect 28623 -31202 28927 -31198
rect 28963 -30902 29587 -30898
rect 28963 -31198 28967 -30902
rect 28967 -31198 29583 -30902
rect 29583 -31198 29587 -30902
rect 28963 -31202 29587 -31198
rect 29623 -30902 29927 -30898
rect 29623 -31198 29627 -30902
rect 29627 -31198 29923 -30902
rect 29923 -31198 29927 -30902
rect 29623 -31202 29927 -31198
rect 29963 -30902 30587 -30898
rect 29963 -31198 29967 -30902
rect 29967 -31198 30583 -30902
rect 30583 -31198 30587 -30902
rect 29963 -31202 30587 -31198
rect 30623 -30902 30927 -30898
rect 30623 -31198 30627 -30902
rect 30627 -31198 30923 -30902
rect 30923 -31198 30927 -30902
rect 30623 -31202 30927 -31198
rect 30963 -30902 31587 -30898
rect 30963 -31198 30967 -30902
rect 30967 -31198 31583 -30902
rect 31583 -31198 31587 -30902
rect 30963 -31202 31587 -31198
rect 31623 -30902 31927 -30898
rect 31623 -31198 31627 -30902
rect 31627 -31198 31923 -30902
rect 31923 -31198 31927 -30902
rect 31623 -31202 31927 -31198
rect 31963 -30902 32587 -30898
rect 31963 -31198 31967 -30902
rect 31967 -31198 32583 -30902
rect 32583 -31198 32587 -30902
rect 31963 -31202 32587 -31198
rect 32623 -30902 32927 -30898
rect 32623 -31198 32627 -30902
rect 32627 -31198 32923 -30902
rect 32923 -31198 32927 -30902
rect 32623 -31202 32927 -31198
rect 32963 -30902 33587 -30898
rect 32963 -31198 32967 -30902
rect 32967 -31198 33583 -30902
rect 33583 -31198 33587 -30902
rect 32963 -31202 33587 -31198
rect 33623 -30902 33927 -30898
rect 33623 -31198 33627 -30902
rect 33627 -31198 33923 -30902
rect 33923 -31198 33927 -30902
rect 33623 -31202 33927 -31198
rect 33963 -30902 34267 -30898
rect 33963 -31198 33967 -30902
rect 33967 -31198 34263 -30902
rect 34263 -31198 34267 -30902
rect 33963 -31202 34267 -31198
rect -74477 -31242 -74173 -31238
rect -74477 -31858 -74473 -31242
rect -74473 -31858 -74177 -31242
rect -74177 -31858 -74173 -31242
rect -74477 -31862 -74173 -31858
rect -73477 -31242 -73173 -31238
rect -73477 -31858 -73473 -31242
rect -73473 -31858 -73177 -31242
rect -73177 -31858 -73173 -31242
rect -73477 -31862 -73173 -31858
rect -72477 -31242 -72173 -31238
rect -72477 -31858 -72473 -31242
rect -72473 -31858 -72177 -31242
rect -72177 -31858 -72173 -31242
rect -72477 -31862 -72173 -31858
rect -71477 -31242 -71173 -31238
rect -71477 -31858 -71473 -31242
rect -71473 -31858 -71177 -31242
rect -71177 -31858 -71173 -31242
rect -71477 -31862 -71173 -31858
rect -70477 -31242 -70173 -31238
rect -70477 -31858 -70473 -31242
rect -70473 -31858 -70177 -31242
rect -70177 -31858 -70173 -31242
rect -70477 -31862 -70173 -31858
rect -69477 -31242 -69173 -31238
rect -69477 -31858 -69473 -31242
rect -69473 -31858 -69177 -31242
rect -69177 -31858 -69173 -31242
rect -69477 -31862 -69173 -31858
rect -68477 -31242 -68173 -31238
rect -68477 -31858 -68473 -31242
rect -68473 -31858 -68177 -31242
rect -68177 -31858 -68173 -31242
rect -68477 -31862 -68173 -31858
rect -67477 -31242 -67173 -31238
rect -67477 -31858 -67473 -31242
rect -67473 -31858 -67177 -31242
rect -67177 -31858 -67173 -31242
rect -67477 -31862 -67173 -31858
rect -66477 -31242 -66173 -31238
rect -66477 -31858 -66473 -31242
rect -66473 -31858 -66177 -31242
rect -66177 -31858 -66173 -31242
rect -66477 -31862 -66173 -31858
rect -65477 -31242 -65173 -31238
rect -65477 -31858 -65473 -31242
rect -65473 -31858 -65177 -31242
rect -65177 -31858 -65173 -31242
rect -65477 -31862 -65173 -31858
rect -64477 -31242 -64173 -31238
rect -64477 -31858 -64473 -31242
rect -64473 -31858 -64177 -31242
rect -64177 -31858 -64173 -31242
rect -64477 -31862 -64173 -31858
rect -63477 -31242 -63173 -31238
rect -63477 -31858 -63473 -31242
rect -63473 -31858 -63177 -31242
rect -63177 -31858 -63173 -31242
rect -63477 -31862 -63173 -31858
rect -62477 -31242 -62173 -31238
rect -62477 -31858 -62473 -31242
rect -62473 -31858 -62177 -31242
rect -62177 -31858 -62173 -31242
rect -62477 -31862 -62173 -31858
rect -61477 -31242 -61173 -31238
rect -61477 -31858 -61473 -31242
rect -61473 -31858 -61177 -31242
rect -61177 -31858 -61173 -31242
rect -61477 -31862 -61173 -31858
rect -60477 -31242 -60173 -31238
rect -60477 -31858 -60473 -31242
rect -60473 -31858 -60177 -31242
rect -60177 -31858 -60173 -31242
rect -60477 -31862 -60173 -31858
rect -59477 -31242 -59173 -31238
rect -59477 -31858 -59473 -31242
rect -59473 -31858 -59177 -31242
rect -59177 -31858 -59173 -31242
rect -59477 -31862 -59173 -31858
rect -58477 -31242 -58173 -31238
rect -58477 -31858 -58473 -31242
rect -58473 -31858 -58177 -31242
rect -58177 -31858 -58173 -31242
rect -58477 -31862 -58173 -31858
rect -57477 -31242 -57173 -31238
rect -57477 -31858 -57473 -31242
rect -57473 -31858 -57177 -31242
rect -57177 -31858 -57173 -31242
rect -57477 -31862 -57173 -31858
rect -56477 -31242 -56173 -31238
rect -56477 -31858 -56473 -31242
rect -56473 -31858 -56177 -31242
rect -56177 -31858 -56173 -31242
rect -56477 -31862 -56173 -31858
rect -55477 -31242 -55173 -31238
rect -55477 -31858 -55473 -31242
rect -55473 -31858 -55177 -31242
rect -55177 -31858 -55173 -31242
rect -55477 -31862 -55173 -31858
rect -54477 -31242 -54173 -31238
rect -54477 -31858 -54473 -31242
rect -54473 -31858 -54177 -31242
rect -54177 -31858 -54173 -31242
rect -54477 -31862 -54173 -31858
rect -53477 -31242 -53173 -31238
rect -53477 -31858 -53473 -31242
rect -53473 -31858 -53177 -31242
rect -53177 -31858 -53173 -31242
rect -53477 -31862 -53173 -31858
rect -52477 -31242 -52173 -31238
rect -52477 -31858 -52473 -31242
rect -52473 -31858 -52177 -31242
rect -52177 -31858 -52173 -31242
rect -52477 -31862 -52173 -31858
rect -51477 -31242 -51173 -31238
rect -51477 -31858 -51473 -31242
rect -51473 -31858 -51177 -31242
rect -51177 -31858 -51173 -31242
rect -51477 -31862 -51173 -31858
rect -50477 -31242 -50173 -31238
rect -50477 -31858 -50473 -31242
rect -50473 -31858 -50177 -31242
rect -50177 -31858 -50173 -31242
rect -50477 -31862 -50173 -31858
rect -49477 -31242 -49173 -31238
rect -49477 -31858 -49473 -31242
rect -49473 -31858 -49177 -31242
rect -49177 -31858 -49173 -31242
rect -49477 -31862 -49173 -31858
rect 8623 -31242 8927 -31238
rect 8623 -31858 8627 -31242
rect 8627 -31858 8923 -31242
rect 8923 -31858 8927 -31242
rect 8623 -31862 8927 -31858
rect 9623 -31242 9927 -31238
rect 9623 -31858 9627 -31242
rect 9627 -31858 9923 -31242
rect 9923 -31858 9927 -31242
rect 9623 -31862 9927 -31858
rect 10623 -31242 10927 -31238
rect 10623 -31858 10627 -31242
rect 10627 -31858 10923 -31242
rect 10923 -31858 10927 -31242
rect 10623 -31862 10927 -31858
rect 11623 -31242 11927 -31238
rect 11623 -31858 11627 -31242
rect 11627 -31858 11923 -31242
rect 11923 -31858 11927 -31242
rect 11623 -31862 11927 -31858
rect 12623 -31242 12927 -31238
rect 12623 -31858 12627 -31242
rect 12627 -31858 12923 -31242
rect 12923 -31858 12927 -31242
rect 12623 -31862 12927 -31858
rect 13623 -31242 13927 -31238
rect 13623 -31858 13627 -31242
rect 13627 -31858 13923 -31242
rect 13923 -31858 13927 -31242
rect 13623 -31862 13927 -31858
rect 14623 -31242 14927 -31238
rect 14623 -31858 14627 -31242
rect 14627 -31858 14923 -31242
rect 14923 -31858 14927 -31242
rect 14623 -31862 14927 -31858
rect 15623 -31242 15927 -31238
rect 15623 -31858 15627 -31242
rect 15627 -31858 15923 -31242
rect 15923 -31858 15927 -31242
rect 15623 -31862 15927 -31858
rect 16623 -31242 16927 -31238
rect 16623 -31858 16627 -31242
rect 16627 -31858 16923 -31242
rect 16923 -31858 16927 -31242
rect 16623 -31862 16927 -31858
rect 17623 -31242 17927 -31238
rect 17623 -31858 17627 -31242
rect 17627 -31858 17923 -31242
rect 17923 -31858 17927 -31242
rect 17623 -31862 17927 -31858
rect 18623 -31242 18927 -31238
rect 18623 -31858 18627 -31242
rect 18627 -31858 18923 -31242
rect 18923 -31858 18927 -31242
rect 18623 -31862 18927 -31858
rect 19623 -31242 19927 -31238
rect 19623 -31858 19627 -31242
rect 19627 -31858 19923 -31242
rect 19923 -31858 19927 -31242
rect 19623 -31862 19927 -31858
rect 20623 -31242 20927 -31238
rect 20623 -31858 20627 -31242
rect 20627 -31858 20923 -31242
rect 20923 -31858 20927 -31242
rect 20623 -31862 20927 -31858
rect 21623 -31242 21927 -31238
rect 21623 -31858 21627 -31242
rect 21627 -31858 21923 -31242
rect 21923 -31858 21927 -31242
rect 21623 -31862 21927 -31858
rect 22623 -31242 22927 -31238
rect 22623 -31858 22627 -31242
rect 22627 -31858 22923 -31242
rect 22923 -31858 22927 -31242
rect 22623 -31862 22927 -31858
rect 23623 -31242 23927 -31238
rect 23623 -31858 23627 -31242
rect 23627 -31858 23923 -31242
rect 23923 -31858 23927 -31242
rect 23623 -31862 23927 -31858
rect 24623 -31242 24927 -31238
rect 24623 -31858 24627 -31242
rect 24627 -31858 24923 -31242
rect 24923 -31858 24927 -31242
rect 24623 -31862 24927 -31858
rect 25623 -31242 25927 -31238
rect 25623 -31858 25627 -31242
rect 25627 -31858 25923 -31242
rect 25923 -31858 25927 -31242
rect 25623 -31862 25927 -31858
rect 26623 -31242 26927 -31238
rect 26623 -31858 26627 -31242
rect 26627 -31858 26923 -31242
rect 26923 -31858 26927 -31242
rect 26623 -31862 26927 -31858
rect 27623 -31242 27927 -31238
rect 27623 -31858 27627 -31242
rect 27627 -31858 27923 -31242
rect 27923 -31858 27927 -31242
rect 27623 -31862 27927 -31858
rect 28623 -31242 28927 -31238
rect 28623 -31858 28627 -31242
rect 28627 -31858 28923 -31242
rect 28923 -31858 28927 -31242
rect 28623 -31862 28927 -31858
rect 29623 -31242 29927 -31238
rect 29623 -31858 29627 -31242
rect 29627 -31858 29923 -31242
rect 29923 -31858 29927 -31242
rect 29623 -31862 29927 -31858
rect 30623 -31242 30927 -31238
rect 30623 -31858 30627 -31242
rect 30627 -31858 30923 -31242
rect 30923 -31858 30927 -31242
rect 30623 -31862 30927 -31858
rect 31623 -31242 31927 -31238
rect 31623 -31858 31627 -31242
rect 31627 -31858 31923 -31242
rect 31923 -31858 31927 -31242
rect 31623 -31862 31927 -31858
rect 32623 -31242 32927 -31238
rect 32623 -31858 32627 -31242
rect 32627 -31858 32923 -31242
rect 32923 -31858 32927 -31242
rect 32623 -31862 32927 -31858
rect 33623 -31242 33927 -31238
rect 33623 -31858 33627 -31242
rect 33627 -31858 33923 -31242
rect 33923 -31858 33927 -31242
rect 33623 -31862 33927 -31858
rect -74817 -31902 -74513 -31898
rect -74817 -32198 -74813 -31902
rect -74813 -32198 -74517 -31902
rect -74517 -32198 -74513 -31902
rect -74817 -32202 -74513 -32198
rect -74477 -31902 -74173 -31898
rect -74477 -32198 -74473 -31902
rect -74473 -32198 -74177 -31902
rect -74177 -32198 -74173 -31902
rect -74477 -32202 -74173 -32198
rect -74137 -31902 -73513 -31898
rect -74137 -32198 -74133 -31902
rect -74133 -32198 -73517 -31902
rect -73517 -32198 -73513 -31902
rect -74137 -32202 -73513 -32198
rect -73477 -31902 -73173 -31898
rect -73477 -32198 -73473 -31902
rect -73473 -32198 -73177 -31902
rect -73177 -32198 -73173 -31902
rect -73477 -32202 -73173 -32198
rect -73137 -31902 -72513 -31898
rect -73137 -32198 -73133 -31902
rect -73133 -32198 -72517 -31902
rect -72517 -32198 -72513 -31902
rect -73137 -32202 -72513 -32198
rect -72477 -31902 -72173 -31898
rect -72477 -32198 -72473 -31902
rect -72473 -32198 -72177 -31902
rect -72177 -32198 -72173 -31902
rect -72477 -32202 -72173 -32198
rect -72137 -31902 -71513 -31898
rect -72137 -32198 -72133 -31902
rect -72133 -32198 -71517 -31902
rect -71517 -32198 -71513 -31902
rect -72137 -32202 -71513 -32198
rect -71477 -31902 -71173 -31898
rect -71477 -32198 -71473 -31902
rect -71473 -32198 -71177 -31902
rect -71177 -32198 -71173 -31902
rect -71477 -32202 -71173 -32198
rect -71137 -31902 -70513 -31898
rect -71137 -32198 -71133 -31902
rect -71133 -32198 -70517 -31902
rect -70517 -32198 -70513 -31902
rect -71137 -32202 -70513 -32198
rect -70477 -31902 -70173 -31898
rect -70477 -32198 -70473 -31902
rect -70473 -32198 -70177 -31902
rect -70177 -32198 -70173 -31902
rect -70477 -32202 -70173 -32198
rect -70137 -31902 -69513 -31898
rect -70137 -32198 -70133 -31902
rect -70133 -32198 -69517 -31902
rect -69517 -32198 -69513 -31902
rect -70137 -32202 -69513 -32198
rect -69477 -31902 -69173 -31898
rect -69477 -32198 -69473 -31902
rect -69473 -32198 -69177 -31902
rect -69177 -32198 -69173 -31902
rect -69477 -32202 -69173 -32198
rect -69137 -31902 -68513 -31898
rect -69137 -32198 -69133 -31902
rect -69133 -32198 -68517 -31902
rect -68517 -32198 -68513 -31902
rect -69137 -32202 -68513 -32198
rect -68477 -31902 -68173 -31898
rect -68477 -32198 -68473 -31902
rect -68473 -32198 -68177 -31902
rect -68177 -32198 -68173 -31902
rect -68477 -32202 -68173 -32198
rect -68137 -31902 -67513 -31898
rect -68137 -32198 -68133 -31902
rect -68133 -32198 -67517 -31902
rect -67517 -32198 -67513 -31902
rect -68137 -32202 -67513 -32198
rect -67477 -31902 -67173 -31898
rect -67477 -32198 -67473 -31902
rect -67473 -32198 -67177 -31902
rect -67177 -32198 -67173 -31902
rect -67477 -32202 -67173 -32198
rect -67137 -31902 -66513 -31898
rect -67137 -32198 -67133 -31902
rect -67133 -32198 -66517 -31902
rect -66517 -32198 -66513 -31902
rect -67137 -32202 -66513 -32198
rect -66477 -31902 -66173 -31898
rect -66477 -32198 -66473 -31902
rect -66473 -32198 -66177 -31902
rect -66177 -32198 -66173 -31902
rect -66477 -32202 -66173 -32198
rect -66137 -31902 -65513 -31898
rect -66137 -32198 -66133 -31902
rect -66133 -32198 -65517 -31902
rect -65517 -32198 -65513 -31902
rect -66137 -32202 -65513 -32198
rect -65477 -31902 -65173 -31898
rect -65477 -32198 -65473 -31902
rect -65473 -32198 -65177 -31902
rect -65177 -32198 -65173 -31902
rect -65477 -32202 -65173 -32198
rect -65137 -31902 -64513 -31898
rect -65137 -32198 -65133 -31902
rect -65133 -32198 -64517 -31902
rect -64517 -32198 -64513 -31902
rect -65137 -32202 -64513 -32198
rect -64477 -31902 -64173 -31898
rect -64477 -32198 -64473 -31902
rect -64473 -32198 -64177 -31902
rect -64177 -32198 -64173 -31902
rect -64477 -32202 -64173 -32198
rect -64137 -31902 -63513 -31898
rect -64137 -32198 -64133 -31902
rect -64133 -32198 -63517 -31902
rect -63517 -32198 -63513 -31902
rect -64137 -32202 -63513 -32198
rect -63477 -31902 -63173 -31898
rect -63477 -32198 -63473 -31902
rect -63473 -32198 -63177 -31902
rect -63177 -32198 -63173 -31902
rect -63477 -32202 -63173 -32198
rect -63137 -31902 -62513 -31898
rect -63137 -32198 -63133 -31902
rect -63133 -32198 -62517 -31902
rect -62517 -32198 -62513 -31902
rect -63137 -32202 -62513 -32198
rect -62477 -31902 -62173 -31898
rect -62477 -32198 -62473 -31902
rect -62473 -32198 -62177 -31902
rect -62177 -32198 -62173 -31902
rect -62477 -32202 -62173 -32198
rect -62137 -31902 -61513 -31898
rect -62137 -32198 -62133 -31902
rect -62133 -32198 -61517 -31902
rect -61517 -32198 -61513 -31902
rect -62137 -32202 -61513 -32198
rect -61477 -31902 -61173 -31898
rect -61477 -32198 -61473 -31902
rect -61473 -32198 -61177 -31902
rect -61177 -32198 -61173 -31902
rect -61477 -32202 -61173 -32198
rect -61137 -31902 -60513 -31898
rect -61137 -32198 -61133 -31902
rect -61133 -32198 -60517 -31902
rect -60517 -32198 -60513 -31902
rect -61137 -32202 -60513 -32198
rect -60477 -31902 -60173 -31898
rect -60477 -32198 -60473 -31902
rect -60473 -32198 -60177 -31902
rect -60177 -32198 -60173 -31902
rect -60477 -32202 -60173 -32198
rect -60137 -31902 -59513 -31898
rect -60137 -32198 -60133 -31902
rect -60133 -32198 -59517 -31902
rect -59517 -32198 -59513 -31902
rect -60137 -32202 -59513 -32198
rect -59477 -31902 -59173 -31898
rect -59477 -32198 -59473 -31902
rect -59473 -32198 -59177 -31902
rect -59177 -32198 -59173 -31902
rect -59477 -32202 -59173 -32198
rect -59137 -31902 -58513 -31898
rect -59137 -32198 -59133 -31902
rect -59133 -32198 -58517 -31902
rect -58517 -32198 -58513 -31902
rect -59137 -32202 -58513 -32198
rect -58477 -31902 -58173 -31898
rect -58477 -32198 -58473 -31902
rect -58473 -32198 -58177 -31902
rect -58177 -32198 -58173 -31902
rect -58477 -32202 -58173 -32198
rect -58137 -31902 -57513 -31898
rect -58137 -32198 -58133 -31902
rect -58133 -32198 -57517 -31902
rect -57517 -32198 -57513 -31902
rect -58137 -32202 -57513 -32198
rect -57477 -31902 -57173 -31898
rect -57477 -32198 -57473 -31902
rect -57473 -32198 -57177 -31902
rect -57177 -32198 -57173 -31902
rect -57477 -32202 -57173 -32198
rect -57137 -31902 -56513 -31898
rect -57137 -32198 -57133 -31902
rect -57133 -32198 -56517 -31902
rect -56517 -32198 -56513 -31902
rect -57137 -32202 -56513 -32198
rect -56477 -31902 -56173 -31898
rect -56477 -32198 -56473 -31902
rect -56473 -32198 -56177 -31902
rect -56177 -32198 -56173 -31902
rect -56477 -32202 -56173 -32198
rect -56137 -31902 -55513 -31898
rect -56137 -32198 -56133 -31902
rect -56133 -32198 -55517 -31902
rect -55517 -32198 -55513 -31902
rect -56137 -32202 -55513 -32198
rect -55477 -31902 -55173 -31898
rect -55477 -32198 -55473 -31902
rect -55473 -32198 -55177 -31902
rect -55177 -32198 -55173 -31902
rect -55477 -32202 -55173 -32198
rect -55137 -31902 -54513 -31898
rect -55137 -32198 -55133 -31902
rect -55133 -32198 -54517 -31902
rect -54517 -32198 -54513 -31902
rect -55137 -32202 -54513 -32198
rect -54477 -31902 -54173 -31898
rect -54477 -32198 -54473 -31902
rect -54473 -32198 -54177 -31902
rect -54177 -32198 -54173 -31902
rect -54477 -32202 -54173 -32198
rect -54137 -31902 -53513 -31898
rect -54137 -32198 -54133 -31902
rect -54133 -32198 -53517 -31902
rect -53517 -32198 -53513 -31902
rect -54137 -32202 -53513 -32198
rect -53477 -31902 -53173 -31898
rect -53477 -32198 -53473 -31902
rect -53473 -32198 -53177 -31902
rect -53177 -32198 -53173 -31902
rect -53477 -32202 -53173 -32198
rect -53137 -31902 -52513 -31898
rect -53137 -32198 -53133 -31902
rect -53133 -32198 -52517 -31902
rect -52517 -32198 -52513 -31902
rect -53137 -32202 -52513 -32198
rect -52477 -31902 -52173 -31898
rect -52477 -32198 -52473 -31902
rect -52473 -32198 -52177 -31902
rect -52177 -32198 -52173 -31902
rect -52477 -32202 -52173 -32198
rect -52137 -31902 -51513 -31898
rect -52137 -32198 -52133 -31902
rect -52133 -32198 -51517 -31902
rect -51517 -32198 -51513 -31902
rect -52137 -32202 -51513 -32198
rect -51477 -31902 -51173 -31898
rect -51477 -32198 -51473 -31902
rect -51473 -32198 -51177 -31902
rect -51177 -32198 -51173 -31902
rect -51477 -32202 -51173 -32198
rect -51137 -31902 -50513 -31898
rect -51137 -32198 -51133 -31902
rect -51133 -32198 -50517 -31902
rect -50517 -32198 -50513 -31902
rect -51137 -32202 -50513 -32198
rect -50477 -31902 -50173 -31898
rect -50477 -32198 -50473 -31902
rect -50473 -32198 -50177 -31902
rect -50177 -32198 -50173 -31902
rect -50477 -32202 -50173 -32198
rect -50137 -31902 -49513 -31898
rect -50137 -32198 -50133 -31902
rect -50133 -32198 -49517 -31902
rect -49517 -32198 -49513 -31902
rect -50137 -32202 -49513 -32198
rect -49477 -31902 -49173 -31898
rect -49477 -32198 -49473 -31902
rect -49473 -32198 -49177 -31902
rect -49177 -32198 -49173 -31902
rect -49477 -32202 -49173 -32198
rect -49137 -31902 -48833 -31898
rect -49137 -32198 -49133 -31902
rect -49133 -32198 -48837 -31902
rect -48837 -32198 -48833 -31902
rect -49137 -32202 -48833 -32198
rect 8283 -31902 8587 -31898
rect 8283 -32198 8287 -31902
rect 8287 -32198 8583 -31902
rect 8583 -32198 8587 -31902
rect 8283 -32202 8587 -32198
rect 8623 -31902 8927 -31898
rect 8623 -32198 8627 -31902
rect 8627 -32198 8923 -31902
rect 8923 -32198 8927 -31902
rect 8623 -32202 8927 -32198
rect 8963 -31902 9587 -31898
rect 8963 -32198 8967 -31902
rect 8967 -32198 9583 -31902
rect 9583 -32198 9587 -31902
rect 8963 -32202 9587 -32198
rect 9623 -31902 9927 -31898
rect 9623 -32198 9627 -31902
rect 9627 -32198 9923 -31902
rect 9923 -32198 9927 -31902
rect 9623 -32202 9927 -32198
rect 9963 -31902 10587 -31898
rect 9963 -32198 9967 -31902
rect 9967 -32198 10583 -31902
rect 10583 -32198 10587 -31902
rect 9963 -32202 10587 -32198
rect 10623 -31902 10927 -31898
rect 10623 -32198 10627 -31902
rect 10627 -32198 10923 -31902
rect 10923 -32198 10927 -31902
rect 10623 -32202 10927 -32198
rect 10963 -31902 11587 -31898
rect 10963 -32198 10967 -31902
rect 10967 -32198 11583 -31902
rect 11583 -32198 11587 -31902
rect 10963 -32202 11587 -32198
rect 11623 -31902 11927 -31898
rect 11623 -32198 11627 -31902
rect 11627 -32198 11923 -31902
rect 11923 -32198 11927 -31902
rect 11623 -32202 11927 -32198
rect 11963 -31902 12587 -31898
rect 11963 -32198 11967 -31902
rect 11967 -32198 12583 -31902
rect 12583 -32198 12587 -31902
rect 11963 -32202 12587 -32198
rect 12623 -31902 12927 -31898
rect 12623 -32198 12627 -31902
rect 12627 -32198 12923 -31902
rect 12923 -32198 12927 -31902
rect 12623 -32202 12927 -32198
rect 12963 -31902 13587 -31898
rect 12963 -32198 12967 -31902
rect 12967 -32198 13583 -31902
rect 13583 -32198 13587 -31902
rect 12963 -32202 13587 -32198
rect 13623 -31902 13927 -31898
rect 13623 -32198 13627 -31902
rect 13627 -32198 13923 -31902
rect 13923 -32198 13927 -31902
rect 13623 -32202 13927 -32198
rect 13963 -31902 14587 -31898
rect 13963 -32198 13967 -31902
rect 13967 -32198 14583 -31902
rect 14583 -32198 14587 -31902
rect 13963 -32202 14587 -32198
rect 14623 -31902 14927 -31898
rect 14623 -32198 14627 -31902
rect 14627 -32198 14923 -31902
rect 14923 -32198 14927 -31902
rect 14623 -32202 14927 -32198
rect 14963 -31902 15587 -31898
rect 14963 -32198 14967 -31902
rect 14967 -32198 15583 -31902
rect 15583 -32198 15587 -31902
rect 14963 -32202 15587 -32198
rect 15623 -31902 15927 -31898
rect 15623 -32198 15627 -31902
rect 15627 -32198 15923 -31902
rect 15923 -32198 15927 -31902
rect 15623 -32202 15927 -32198
rect 15963 -31902 16587 -31898
rect 15963 -32198 15967 -31902
rect 15967 -32198 16583 -31902
rect 16583 -32198 16587 -31902
rect 15963 -32202 16587 -32198
rect 16623 -31902 16927 -31898
rect 16623 -32198 16627 -31902
rect 16627 -32198 16923 -31902
rect 16923 -32198 16927 -31902
rect 16623 -32202 16927 -32198
rect 16963 -31902 17587 -31898
rect 16963 -32198 16967 -31902
rect 16967 -32198 17583 -31902
rect 17583 -32198 17587 -31902
rect 16963 -32202 17587 -32198
rect 17623 -31902 17927 -31898
rect 17623 -32198 17627 -31902
rect 17627 -32198 17923 -31902
rect 17923 -32198 17927 -31902
rect 17623 -32202 17927 -32198
rect 17963 -31902 18587 -31898
rect 17963 -32198 17967 -31902
rect 17967 -32198 18583 -31902
rect 18583 -32198 18587 -31902
rect 17963 -32202 18587 -32198
rect 18623 -31902 18927 -31898
rect 18623 -32198 18627 -31902
rect 18627 -32198 18923 -31902
rect 18923 -32198 18927 -31902
rect 18623 -32202 18927 -32198
rect 18963 -31902 19587 -31898
rect 18963 -32198 18967 -31902
rect 18967 -32198 19583 -31902
rect 19583 -32198 19587 -31902
rect 18963 -32202 19587 -32198
rect 19623 -31902 19927 -31898
rect 19623 -32198 19627 -31902
rect 19627 -32198 19923 -31902
rect 19923 -32198 19927 -31902
rect 19623 -32202 19927 -32198
rect 19963 -31902 20587 -31898
rect 19963 -32198 19967 -31902
rect 19967 -32198 20583 -31902
rect 20583 -32198 20587 -31902
rect 19963 -32202 20587 -32198
rect 20623 -31902 20927 -31898
rect 20623 -32198 20627 -31902
rect 20627 -32198 20923 -31902
rect 20923 -32198 20927 -31902
rect 20623 -32202 20927 -32198
rect 20963 -31902 21587 -31898
rect 20963 -32198 20967 -31902
rect 20967 -32198 21583 -31902
rect 21583 -32198 21587 -31902
rect 20963 -32202 21587 -32198
rect 21623 -31902 21927 -31898
rect 21623 -32198 21627 -31902
rect 21627 -32198 21923 -31902
rect 21923 -32198 21927 -31902
rect 21623 -32202 21927 -32198
rect 21963 -31902 22587 -31898
rect 21963 -32198 21967 -31902
rect 21967 -32198 22583 -31902
rect 22583 -32198 22587 -31902
rect 21963 -32202 22587 -32198
rect 22623 -31902 22927 -31898
rect 22623 -32198 22627 -31902
rect 22627 -32198 22923 -31902
rect 22923 -32198 22927 -31902
rect 22623 -32202 22927 -32198
rect 22963 -31902 23587 -31898
rect 22963 -32198 22967 -31902
rect 22967 -32198 23583 -31902
rect 23583 -32198 23587 -31902
rect 22963 -32202 23587 -32198
rect 23623 -31902 23927 -31898
rect 23623 -32198 23627 -31902
rect 23627 -32198 23923 -31902
rect 23923 -32198 23927 -31902
rect 23623 -32202 23927 -32198
rect 23963 -31902 24587 -31898
rect 23963 -32198 23967 -31902
rect 23967 -32198 24583 -31902
rect 24583 -32198 24587 -31902
rect 23963 -32202 24587 -32198
rect 24623 -31902 24927 -31898
rect 24623 -32198 24627 -31902
rect 24627 -32198 24923 -31902
rect 24923 -32198 24927 -31902
rect 24623 -32202 24927 -32198
rect 24963 -31902 25587 -31898
rect 24963 -32198 24967 -31902
rect 24967 -32198 25583 -31902
rect 25583 -32198 25587 -31902
rect 24963 -32202 25587 -32198
rect 25623 -31902 25927 -31898
rect 25623 -32198 25627 -31902
rect 25627 -32198 25923 -31902
rect 25923 -32198 25927 -31902
rect 25623 -32202 25927 -32198
rect 25963 -31902 26587 -31898
rect 25963 -32198 25967 -31902
rect 25967 -32198 26583 -31902
rect 26583 -32198 26587 -31902
rect 25963 -32202 26587 -32198
rect 26623 -31902 26927 -31898
rect 26623 -32198 26627 -31902
rect 26627 -32198 26923 -31902
rect 26923 -32198 26927 -31902
rect 26623 -32202 26927 -32198
rect 26963 -31902 27587 -31898
rect 26963 -32198 26967 -31902
rect 26967 -32198 27583 -31902
rect 27583 -32198 27587 -31902
rect 26963 -32202 27587 -32198
rect 27623 -31902 27927 -31898
rect 27623 -32198 27627 -31902
rect 27627 -32198 27923 -31902
rect 27923 -32198 27927 -31902
rect 27623 -32202 27927 -32198
rect 27963 -31902 28587 -31898
rect 27963 -32198 27967 -31902
rect 27967 -32198 28583 -31902
rect 28583 -32198 28587 -31902
rect 27963 -32202 28587 -32198
rect 28623 -31902 28927 -31898
rect 28623 -32198 28627 -31902
rect 28627 -32198 28923 -31902
rect 28923 -32198 28927 -31902
rect 28623 -32202 28927 -32198
rect 28963 -31902 29587 -31898
rect 28963 -32198 28967 -31902
rect 28967 -32198 29583 -31902
rect 29583 -32198 29587 -31902
rect 28963 -32202 29587 -32198
rect 29623 -31902 29927 -31898
rect 29623 -32198 29627 -31902
rect 29627 -32198 29923 -31902
rect 29923 -32198 29927 -31902
rect 29623 -32202 29927 -32198
rect 29963 -31902 30587 -31898
rect 29963 -32198 29967 -31902
rect 29967 -32198 30583 -31902
rect 30583 -32198 30587 -31902
rect 29963 -32202 30587 -32198
rect 30623 -31902 30927 -31898
rect 30623 -32198 30627 -31902
rect 30627 -32198 30923 -31902
rect 30923 -32198 30927 -31902
rect 30623 -32202 30927 -32198
rect 30963 -31902 31587 -31898
rect 30963 -32198 30967 -31902
rect 30967 -32198 31583 -31902
rect 31583 -32198 31587 -31902
rect 30963 -32202 31587 -32198
rect 31623 -31902 31927 -31898
rect 31623 -32198 31627 -31902
rect 31627 -32198 31923 -31902
rect 31923 -32198 31927 -31902
rect 31623 -32202 31927 -32198
rect 31963 -31902 32587 -31898
rect 31963 -32198 31967 -31902
rect 31967 -32198 32583 -31902
rect 32583 -32198 32587 -31902
rect 31963 -32202 32587 -32198
rect 32623 -31902 32927 -31898
rect 32623 -32198 32627 -31902
rect 32627 -32198 32923 -31902
rect 32923 -32198 32927 -31902
rect 32623 -32202 32927 -32198
rect 32963 -31902 33587 -31898
rect 32963 -32198 32967 -31902
rect 32967 -32198 33583 -31902
rect 33583 -32198 33587 -31902
rect 32963 -32202 33587 -32198
rect 33623 -31902 33927 -31898
rect 33623 -32198 33627 -31902
rect 33627 -32198 33923 -31902
rect 33923 -32198 33927 -31902
rect 33623 -32202 33927 -32198
rect 33963 -31902 34267 -31898
rect 33963 -32198 33967 -31902
rect 33967 -32198 34263 -31902
rect 34263 -32198 34267 -31902
rect 33963 -32202 34267 -32198
rect -74477 -32242 -74173 -32238
rect -74477 -32858 -74473 -32242
rect -74473 -32858 -74177 -32242
rect -74177 -32858 -74173 -32242
rect -74477 -32862 -74173 -32858
rect -73477 -32242 -73173 -32238
rect -73477 -32858 -73473 -32242
rect -73473 -32858 -73177 -32242
rect -73177 -32858 -73173 -32242
rect -73477 -32862 -73173 -32858
rect -72477 -32242 -72173 -32238
rect -72477 -32858 -72473 -32242
rect -72473 -32858 -72177 -32242
rect -72177 -32858 -72173 -32242
rect -72477 -32862 -72173 -32858
rect -71477 -32242 -71173 -32238
rect -71477 -32858 -71473 -32242
rect -71473 -32858 -71177 -32242
rect -71177 -32858 -71173 -32242
rect -71477 -32862 -71173 -32858
rect -70477 -32242 -70173 -32238
rect -70477 -32858 -70473 -32242
rect -70473 -32858 -70177 -32242
rect -70177 -32858 -70173 -32242
rect -70477 -32862 -70173 -32858
rect -69477 -32242 -69173 -32238
rect -69477 -32858 -69473 -32242
rect -69473 -32858 -69177 -32242
rect -69177 -32858 -69173 -32242
rect -69477 -32862 -69173 -32858
rect -68477 -32242 -68173 -32238
rect -68477 -32858 -68473 -32242
rect -68473 -32858 -68177 -32242
rect -68177 -32858 -68173 -32242
rect -68477 -32862 -68173 -32858
rect -67477 -32242 -67173 -32238
rect -67477 -32858 -67473 -32242
rect -67473 -32858 -67177 -32242
rect -67177 -32858 -67173 -32242
rect -67477 -32862 -67173 -32858
rect -66477 -32242 -66173 -32238
rect -66477 -32858 -66473 -32242
rect -66473 -32858 -66177 -32242
rect -66177 -32858 -66173 -32242
rect -66477 -32862 -66173 -32858
rect -65477 -32242 -65173 -32238
rect -65477 -32858 -65473 -32242
rect -65473 -32858 -65177 -32242
rect -65177 -32858 -65173 -32242
rect -65477 -32862 -65173 -32858
rect -64477 -32242 -64173 -32238
rect -64477 -32858 -64473 -32242
rect -64473 -32858 -64177 -32242
rect -64177 -32858 -64173 -32242
rect -64477 -32862 -64173 -32858
rect -63477 -32242 -63173 -32238
rect -63477 -32858 -63473 -32242
rect -63473 -32858 -63177 -32242
rect -63177 -32858 -63173 -32242
rect -63477 -32862 -63173 -32858
rect -62477 -32242 -62173 -32238
rect -62477 -32858 -62473 -32242
rect -62473 -32858 -62177 -32242
rect -62177 -32858 -62173 -32242
rect -62477 -32862 -62173 -32858
rect -61477 -32242 -61173 -32238
rect -61477 -32858 -61473 -32242
rect -61473 -32858 -61177 -32242
rect -61177 -32858 -61173 -32242
rect -61477 -32862 -61173 -32858
rect -60477 -32242 -60173 -32238
rect -60477 -32858 -60473 -32242
rect -60473 -32858 -60177 -32242
rect -60177 -32858 -60173 -32242
rect -60477 -32862 -60173 -32858
rect -59477 -32242 -59173 -32238
rect -59477 -32858 -59473 -32242
rect -59473 -32858 -59177 -32242
rect -59177 -32858 -59173 -32242
rect -59477 -32862 -59173 -32858
rect -58477 -32242 -58173 -32238
rect -58477 -32858 -58473 -32242
rect -58473 -32858 -58177 -32242
rect -58177 -32858 -58173 -32242
rect -58477 -32862 -58173 -32858
rect -57477 -32242 -57173 -32238
rect -57477 -32858 -57473 -32242
rect -57473 -32858 -57177 -32242
rect -57177 -32858 -57173 -32242
rect -57477 -32862 -57173 -32858
rect -56477 -32242 -56173 -32238
rect -56477 -32858 -56473 -32242
rect -56473 -32858 -56177 -32242
rect -56177 -32858 -56173 -32242
rect -56477 -32862 -56173 -32858
rect -55477 -32242 -55173 -32238
rect -55477 -32858 -55473 -32242
rect -55473 -32858 -55177 -32242
rect -55177 -32858 -55173 -32242
rect -55477 -32862 -55173 -32858
rect -54477 -32242 -54173 -32238
rect -54477 -32858 -54473 -32242
rect -54473 -32858 -54177 -32242
rect -54177 -32858 -54173 -32242
rect -54477 -32862 -54173 -32858
rect -53477 -32242 -53173 -32238
rect -53477 -32858 -53473 -32242
rect -53473 -32858 -53177 -32242
rect -53177 -32858 -53173 -32242
rect -53477 -32862 -53173 -32858
rect -52477 -32242 -52173 -32238
rect -52477 -32858 -52473 -32242
rect -52473 -32858 -52177 -32242
rect -52177 -32858 -52173 -32242
rect -52477 -32862 -52173 -32858
rect -51477 -32242 -51173 -32238
rect -51477 -32858 -51473 -32242
rect -51473 -32858 -51177 -32242
rect -51177 -32858 -51173 -32242
rect -51477 -32862 -51173 -32858
rect -50477 -32242 -50173 -32238
rect -50477 -32858 -50473 -32242
rect -50473 -32858 -50177 -32242
rect -50177 -32858 -50173 -32242
rect -50477 -32862 -50173 -32858
rect -49477 -32242 -49173 -32238
rect -49477 -32858 -49473 -32242
rect -49473 -32858 -49177 -32242
rect -49177 -32858 -49173 -32242
rect -49477 -32862 -49173 -32858
rect -74817 -32902 -74513 -32898
rect -74817 -33198 -74813 -32902
rect -74813 -33198 -74517 -32902
rect -74517 -33198 -74513 -32902
rect -74817 -33202 -74513 -33198
rect -74477 -32902 -74173 -32898
rect -74477 -33198 -74473 -32902
rect -74473 -33198 -74177 -32902
rect -74177 -33198 -74173 -32902
rect -74477 -33202 -74173 -33198
rect -74137 -32902 -73513 -32898
rect -74137 -33198 -74133 -32902
rect -74133 -33198 -73517 -32902
rect -73517 -33198 -73513 -32902
rect -74137 -33202 -73513 -33198
rect -73477 -32902 -73173 -32898
rect -73477 -33198 -73473 -32902
rect -73473 -33198 -73177 -32902
rect -73177 -33198 -73173 -32902
rect -73477 -33202 -73173 -33198
rect -73137 -32902 -72513 -32898
rect -73137 -33198 -73133 -32902
rect -73133 -33198 -72517 -32902
rect -72517 -33198 -72513 -32902
rect -73137 -33202 -72513 -33198
rect -72477 -32902 -72173 -32898
rect -72477 -33198 -72473 -32902
rect -72473 -33198 -72177 -32902
rect -72177 -33198 -72173 -32902
rect -72477 -33202 -72173 -33198
rect -72137 -32902 -71513 -32898
rect -72137 -33198 -72133 -32902
rect -72133 -33198 -71517 -32902
rect -71517 -33198 -71513 -32902
rect -72137 -33202 -71513 -33198
rect -71477 -32902 -71173 -32898
rect -71477 -33198 -71473 -32902
rect -71473 -33198 -71177 -32902
rect -71177 -33198 -71173 -32902
rect -71477 -33202 -71173 -33198
rect -71137 -32902 -70513 -32898
rect -71137 -33198 -71133 -32902
rect -71133 -33198 -70517 -32902
rect -70517 -33198 -70513 -32902
rect -71137 -33202 -70513 -33198
rect -70477 -32902 -70173 -32898
rect -70477 -33198 -70473 -32902
rect -70473 -33198 -70177 -32902
rect -70177 -33198 -70173 -32902
rect -70477 -33202 -70173 -33198
rect -70137 -32902 -69513 -32898
rect -70137 -33198 -70133 -32902
rect -70133 -33198 -69517 -32902
rect -69517 -33198 -69513 -32902
rect -70137 -33202 -69513 -33198
rect -69477 -32902 -69173 -32898
rect -69477 -33198 -69473 -32902
rect -69473 -33198 -69177 -32902
rect -69177 -33198 -69173 -32902
rect -69477 -33202 -69173 -33198
rect -69137 -32902 -68513 -32898
rect -69137 -33198 -69133 -32902
rect -69133 -33198 -68517 -32902
rect -68517 -33198 -68513 -32902
rect -69137 -33202 -68513 -33198
rect -68477 -32902 -68173 -32898
rect -68477 -33198 -68473 -32902
rect -68473 -33198 -68177 -32902
rect -68177 -33198 -68173 -32902
rect -68477 -33202 -68173 -33198
rect -68137 -32902 -67513 -32898
rect -68137 -33198 -68133 -32902
rect -68133 -33198 -67517 -32902
rect -67517 -33198 -67513 -32902
rect -68137 -33202 -67513 -33198
rect -67477 -32902 -67173 -32898
rect -67477 -33198 -67473 -32902
rect -67473 -33198 -67177 -32902
rect -67177 -33198 -67173 -32902
rect -67477 -33202 -67173 -33198
rect -67137 -32902 -66513 -32898
rect -67137 -33198 -67133 -32902
rect -67133 -33198 -66517 -32902
rect -66517 -33198 -66513 -32902
rect -67137 -33202 -66513 -33198
rect -66477 -32902 -66173 -32898
rect -66477 -33198 -66473 -32902
rect -66473 -33198 -66177 -32902
rect -66177 -33198 -66173 -32902
rect -66477 -33202 -66173 -33198
rect -66137 -32902 -65513 -32898
rect -66137 -33198 -66133 -32902
rect -66133 -33198 -65517 -32902
rect -65517 -33198 -65513 -32902
rect -66137 -33202 -65513 -33198
rect -65477 -32902 -65173 -32898
rect -65477 -33198 -65473 -32902
rect -65473 -33198 -65177 -32902
rect -65177 -33198 -65173 -32902
rect -65477 -33202 -65173 -33198
rect -65137 -32902 -64513 -32898
rect -65137 -33198 -65133 -32902
rect -65133 -33198 -64517 -32902
rect -64517 -33198 -64513 -32902
rect -65137 -33202 -64513 -33198
rect -64477 -32902 -64173 -32898
rect -64477 -33198 -64473 -32902
rect -64473 -33198 -64177 -32902
rect -64177 -33198 -64173 -32902
rect -64477 -33202 -64173 -33198
rect -64137 -32902 -63513 -32898
rect -64137 -33198 -64133 -32902
rect -64133 -33198 -63517 -32902
rect -63517 -33198 -63513 -32902
rect -64137 -33202 -63513 -33198
rect -63477 -32902 -63173 -32898
rect -63477 -33198 -63473 -32902
rect -63473 -33198 -63177 -32902
rect -63177 -33198 -63173 -32902
rect -63477 -33202 -63173 -33198
rect -63137 -32902 -62513 -32898
rect -63137 -33198 -63133 -32902
rect -63133 -33198 -62517 -32902
rect -62517 -33198 -62513 -32902
rect -63137 -33202 -62513 -33198
rect -62477 -32902 -62173 -32898
rect -62477 -33198 -62473 -32902
rect -62473 -33198 -62177 -32902
rect -62177 -33198 -62173 -32902
rect -62477 -33202 -62173 -33198
rect -62137 -32902 -61513 -32898
rect -62137 -33198 -62133 -32902
rect -62133 -33198 -61517 -32902
rect -61517 -33198 -61513 -32902
rect -62137 -33202 -61513 -33198
rect -61477 -32902 -61173 -32898
rect -61477 -33198 -61473 -32902
rect -61473 -33198 -61177 -32902
rect -61177 -33198 -61173 -32902
rect -61477 -33202 -61173 -33198
rect -61137 -32902 -60513 -32898
rect -61137 -33198 -61133 -32902
rect -61133 -33198 -60517 -32902
rect -60517 -33198 -60513 -32902
rect -61137 -33202 -60513 -33198
rect -60477 -32902 -60173 -32898
rect -60477 -33198 -60473 -32902
rect -60473 -33198 -60177 -32902
rect -60177 -33198 -60173 -32902
rect -60477 -33202 -60173 -33198
rect -60137 -32902 -59513 -32898
rect -60137 -33198 -60133 -32902
rect -60133 -33198 -59517 -32902
rect -59517 -33198 -59513 -32902
rect -60137 -33202 -59513 -33198
rect -59477 -32902 -59173 -32898
rect -59477 -33198 -59473 -32902
rect -59473 -33198 -59177 -32902
rect -59177 -33198 -59173 -32902
rect -59477 -33202 -59173 -33198
rect -59137 -32902 -58513 -32898
rect -59137 -33198 -59133 -32902
rect -59133 -33198 -58517 -32902
rect -58517 -33198 -58513 -32902
rect -59137 -33202 -58513 -33198
rect -58477 -32902 -58173 -32898
rect -58477 -33198 -58473 -32902
rect -58473 -33198 -58177 -32902
rect -58177 -33198 -58173 -32902
rect -58477 -33202 -58173 -33198
rect -58137 -32902 -57513 -32898
rect -58137 -33198 -58133 -32902
rect -58133 -33198 -57517 -32902
rect -57517 -33198 -57513 -32902
rect -58137 -33202 -57513 -33198
rect -57477 -32902 -57173 -32898
rect -57477 -33198 -57473 -32902
rect -57473 -33198 -57177 -32902
rect -57177 -33198 -57173 -32902
rect -57477 -33202 -57173 -33198
rect -57137 -32902 -56513 -32898
rect -57137 -33198 -57133 -32902
rect -57133 -33198 -56517 -32902
rect -56517 -33198 -56513 -32902
rect -57137 -33202 -56513 -33198
rect -56477 -32902 -56173 -32898
rect -56477 -33198 -56473 -32902
rect -56473 -33198 -56177 -32902
rect -56177 -33198 -56173 -32902
rect -56477 -33202 -56173 -33198
rect -56137 -32902 -55513 -32898
rect -56137 -33198 -56133 -32902
rect -56133 -33198 -55517 -32902
rect -55517 -33198 -55513 -32902
rect -56137 -33202 -55513 -33198
rect -55477 -32902 -55173 -32898
rect -55477 -33198 -55473 -32902
rect -55473 -33198 -55177 -32902
rect -55177 -33198 -55173 -32902
rect -55477 -33202 -55173 -33198
rect -55137 -32902 -54513 -32898
rect -55137 -33198 -55133 -32902
rect -55133 -33198 -54517 -32902
rect -54517 -33198 -54513 -32902
rect -55137 -33202 -54513 -33198
rect -54477 -32902 -54173 -32898
rect -54477 -33198 -54473 -32902
rect -54473 -33198 -54177 -32902
rect -54177 -33198 -54173 -32902
rect -54477 -33202 -54173 -33198
rect -54137 -32902 -53513 -32898
rect -54137 -33198 -54133 -32902
rect -54133 -33198 -53517 -32902
rect -53517 -33198 -53513 -32902
rect -54137 -33202 -53513 -33198
rect -53477 -32902 -53173 -32898
rect -53477 -33198 -53473 -32902
rect -53473 -33198 -53177 -32902
rect -53177 -33198 -53173 -32902
rect -53477 -33202 -53173 -33198
rect -53137 -32902 -52513 -32898
rect -53137 -33198 -53133 -32902
rect -53133 -33198 -52517 -32902
rect -52517 -33198 -52513 -32902
rect -53137 -33202 -52513 -33198
rect -52477 -32902 -52173 -32898
rect -52477 -33198 -52473 -32902
rect -52473 -33198 -52177 -32902
rect -52177 -33198 -52173 -32902
rect -52477 -33202 -52173 -33198
rect -52137 -32902 -51513 -32898
rect -52137 -33198 -52133 -32902
rect -52133 -33198 -51517 -32902
rect -51517 -33198 -51513 -32902
rect -52137 -33202 -51513 -33198
rect -51477 -32902 -51173 -32898
rect -51477 -33198 -51473 -32902
rect -51473 -33198 -51177 -32902
rect -51177 -33198 -51173 -32902
rect -51477 -33202 -51173 -33198
rect -51137 -32902 -50513 -32898
rect -51137 -33198 -51133 -32902
rect -51133 -33198 -50517 -32902
rect -50517 -33198 -50513 -32902
rect -51137 -33202 -50513 -33198
rect -50477 -32902 -50173 -32898
rect -50477 -33198 -50473 -32902
rect -50473 -33198 -50177 -32902
rect -50177 -33198 -50173 -32902
rect -50477 -33202 -50173 -33198
rect -50137 -32902 -49513 -32898
rect -50137 -33198 -50133 -32902
rect -50133 -33198 -49517 -32902
rect -49517 -33198 -49513 -32902
rect -50137 -33202 -49513 -33198
rect -49477 -32902 -49173 -32898
rect -49477 -33198 -49473 -32902
rect -49473 -33198 -49177 -32902
rect -49177 -33198 -49173 -32902
rect -49477 -33202 -49173 -33198
rect -49137 -32902 -48833 -32898
rect -49137 -33198 -49133 -32902
rect -49133 -33198 -48837 -32902
rect -48837 -33198 -48833 -32902
rect -49137 -33202 -48833 -33198
rect -74477 -33242 -74173 -33238
rect -74477 -33858 -74473 -33242
rect -74473 -33858 -74177 -33242
rect -74177 -33858 -74173 -33242
rect -74477 -33862 -74173 -33858
rect -73477 -33242 -73173 -33238
rect -73477 -33858 -73473 -33242
rect -73473 -33858 -73177 -33242
rect -73177 -33858 -73173 -33242
rect -73477 -33862 -73173 -33858
rect -72477 -33242 -72173 -33238
rect -72477 -33858 -72473 -33242
rect -72473 -33858 -72177 -33242
rect -72177 -33858 -72173 -33242
rect -72477 -33862 -72173 -33858
rect -71477 -33242 -71173 -33238
rect -71477 -33858 -71473 -33242
rect -71473 -33858 -71177 -33242
rect -71177 -33858 -71173 -33242
rect -71477 -33862 -71173 -33858
rect -70477 -33242 -70173 -33238
rect -70477 -33858 -70473 -33242
rect -70473 -33858 -70177 -33242
rect -70177 -33858 -70173 -33242
rect -70477 -33862 -70173 -33858
rect -69477 -33242 -69173 -33238
rect -69477 -33858 -69473 -33242
rect -69473 -33858 -69177 -33242
rect -69177 -33858 -69173 -33242
rect -69477 -33862 -69173 -33858
rect -68477 -33242 -68173 -33238
rect -68477 -33858 -68473 -33242
rect -68473 -33858 -68177 -33242
rect -68177 -33858 -68173 -33242
rect -68477 -33862 -68173 -33858
rect -67477 -33242 -67173 -33238
rect -67477 -33858 -67473 -33242
rect -67473 -33858 -67177 -33242
rect -67177 -33858 -67173 -33242
rect -67477 -33862 -67173 -33858
rect -66477 -33242 -66173 -33238
rect -66477 -33858 -66473 -33242
rect -66473 -33858 -66177 -33242
rect -66177 -33858 -66173 -33242
rect -66477 -33862 -66173 -33858
rect -65477 -33242 -65173 -33238
rect -65477 -33858 -65473 -33242
rect -65473 -33858 -65177 -33242
rect -65177 -33858 -65173 -33242
rect -65477 -33862 -65173 -33858
rect -64477 -33242 -64173 -33238
rect -64477 -33858 -64473 -33242
rect -64473 -33858 -64177 -33242
rect -64177 -33858 -64173 -33242
rect -64477 -33862 -64173 -33858
rect -63477 -33242 -63173 -33238
rect -63477 -33858 -63473 -33242
rect -63473 -33858 -63177 -33242
rect -63177 -33858 -63173 -33242
rect -63477 -33862 -63173 -33858
rect -62477 -33242 -62173 -33238
rect -62477 -33858 -62473 -33242
rect -62473 -33858 -62177 -33242
rect -62177 -33858 -62173 -33242
rect -62477 -33862 -62173 -33858
rect -61477 -33242 -61173 -33238
rect -61477 -33858 -61473 -33242
rect -61473 -33858 -61177 -33242
rect -61177 -33858 -61173 -33242
rect -61477 -33862 -61173 -33858
rect -60477 -33242 -60173 -33238
rect -60477 -33858 -60473 -33242
rect -60473 -33858 -60177 -33242
rect -60177 -33858 -60173 -33242
rect -60477 -33862 -60173 -33858
rect -59477 -33242 -59173 -33238
rect -59477 -33858 -59473 -33242
rect -59473 -33858 -59177 -33242
rect -59177 -33858 -59173 -33242
rect -59477 -33862 -59173 -33858
rect -58477 -33242 -58173 -33238
rect -58477 -33858 -58473 -33242
rect -58473 -33858 -58177 -33242
rect -58177 -33858 -58173 -33242
rect -58477 -33862 -58173 -33858
rect -57477 -33242 -57173 -33238
rect -57477 -33858 -57473 -33242
rect -57473 -33858 -57177 -33242
rect -57177 -33858 -57173 -33242
rect -57477 -33862 -57173 -33858
rect -56477 -33242 -56173 -33238
rect -56477 -33858 -56473 -33242
rect -56473 -33858 -56177 -33242
rect -56177 -33858 -56173 -33242
rect -56477 -33862 -56173 -33858
rect -55477 -33242 -55173 -33238
rect -55477 -33858 -55473 -33242
rect -55473 -33858 -55177 -33242
rect -55177 -33858 -55173 -33242
rect -55477 -33862 -55173 -33858
rect -54477 -33242 -54173 -33238
rect -54477 -33858 -54473 -33242
rect -54473 -33858 -54177 -33242
rect -54177 -33858 -54173 -33242
rect -54477 -33862 -54173 -33858
rect -53477 -33242 -53173 -33238
rect -53477 -33858 -53473 -33242
rect -53473 -33858 -53177 -33242
rect -53177 -33858 -53173 -33242
rect -53477 -33862 -53173 -33858
rect -52477 -33242 -52173 -33238
rect -52477 -33858 -52473 -33242
rect -52473 -33858 -52177 -33242
rect -52177 -33858 -52173 -33242
rect -52477 -33862 -52173 -33858
rect -51477 -33242 -51173 -33238
rect -51477 -33858 -51473 -33242
rect -51473 -33858 -51177 -33242
rect -51177 -33858 -51173 -33242
rect -51477 -33862 -51173 -33858
rect -50477 -33242 -50173 -33238
rect -50477 -33858 -50473 -33242
rect -50473 -33858 -50177 -33242
rect -50177 -33858 -50173 -33242
rect -50477 -33862 -50173 -33858
rect -49477 -33242 -49173 -33238
rect -49477 -33858 -49473 -33242
rect -49473 -33858 -49177 -33242
rect -49177 -33858 -49173 -33242
rect -49477 -33862 -49173 -33858
rect -74817 -33902 -74513 -33898
rect -74817 -34198 -74813 -33902
rect -74813 -34198 -74517 -33902
rect -74517 -34198 -74513 -33902
rect -74817 -34202 -74513 -34198
rect -74477 -33902 -74173 -33898
rect -74477 -34198 -74473 -33902
rect -74473 -34198 -74177 -33902
rect -74177 -34198 -74173 -33902
rect -74477 -34202 -74173 -34198
rect -74137 -33902 -73513 -33898
rect -74137 -34198 -74133 -33902
rect -74133 -34198 -73517 -33902
rect -73517 -34198 -73513 -33902
rect -74137 -34202 -73513 -34198
rect -73477 -33902 -73173 -33898
rect -73477 -34198 -73473 -33902
rect -73473 -34198 -73177 -33902
rect -73177 -34198 -73173 -33902
rect -73477 -34202 -73173 -34198
rect -73137 -33902 -72513 -33898
rect -73137 -34198 -73133 -33902
rect -73133 -34198 -72517 -33902
rect -72517 -34198 -72513 -33902
rect -73137 -34202 -72513 -34198
rect -72477 -33902 -72173 -33898
rect -72477 -34198 -72473 -33902
rect -72473 -34198 -72177 -33902
rect -72177 -34198 -72173 -33902
rect -72477 -34202 -72173 -34198
rect -72137 -33902 -71513 -33898
rect -72137 -34198 -72133 -33902
rect -72133 -34198 -71517 -33902
rect -71517 -34198 -71513 -33902
rect -72137 -34202 -71513 -34198
rect -71477 -33902 -71173 -33898
rect -71477 -34198 -71473 -33902
rect -71473 -34198 -71177 -33902
rect -71177 -34198 -71173 -33902
rect -71477 -34202 -71173 -34198
rect -71137 -33902 -70513 -33898
rect -71137 -34198 -71133 -33902
rect -71133 -34198 -70517 -33902
rect -70517 -34198 -70513 -33902
rect -71137 -34202 -70513 -34198
rect -70477 -33902 -70173 -33898
rect -70477 -34198 -70473 -33902
rect -70473 -34198 -70177 -33902
rect -70177 -34198 -70173 -33902
rect -70477 -34202 -70173 -34198
rect -70137 -33902 -69513 -33898
rect -70137 -34198 -70133 -33902
rect -70133 -34198 -69517 -33902
rect -69517 -34198 -69513 -33902
rect -70137 -34202 -69513 -34198
rect -69477 -33902 -69173 -33898
rect -69477 -34198 -69473 -33902
rect -69473 -34198 -69177 -33902
rect -69177 -34198 -69173 -33902
rect -69477 -34202 -69173 -34198
rect -69137 -33902 -68513 -33898
rect -69137 -34198 -69133 -33902
rect -69133 -34198 -68517 -33902
rect -68517 -34198 -68513 -33902
rect -69137 -34202 -68513 -34198
rect -68477 -33902 -68173 -33898
rect -68477 -34198 -68473 -33902
rect -68473 -34198 -68177 -33902
rect -68177 -34198 -68173 -33902
rect -68477 -34202 -68173 -34198
rect -68137 -33902 -67513 -33898
rect -68137 -34198 -68133 -33902
rect -68133 -34198 -67517 -33902
rect -67517 -34198 -67513 -33902
rect -68137 -34202 -67513 -34198
rect -67477 -33902 -67173 -33898
rect -67477 -34198 -67473 -33902
rect -67473 -34198 -67177 -33902
rect -67177 -34198 -67173 -33902
rect -67477 -34202 -67173 -34198
rect -67137 -33902 -66513 -33898
rect -67137 -34198 -67133 -33902
rect -67133 -34198 -66517 -33902
rect -66517 -34198 -66513 -33902
rect -67137 -34202 -66513 -34198
rect -66477 -33902 -66173 -33898
rect -66477 -34198 -66473 -33902
rect -66473 -34198 -66177 -33902
rect -66177 -34198 -66173 -33902
rect -66477 -34202 -66173 -34198
rect -66137 -33902 -65513 -33898
rect -66137 -34198 -66133 -33902
rect -66133 -34198 -65517 -33902
rect -65517 -34198 -65513 -33902
rect -66137 -34202 -65513 -34198
rect -65477 -33902 -65173 -33898
rect -65477 -34198 -65473 -33902
rect -65473 -34198 -65177 -33902
rect -65177 -34198 -65173 -33902
rect -65477 -34202 -65173 -34198
rect -65137 -33902 -64513 -33898
rect -65137 -34198 -65133 -33902
rect -65133 -34198 -64517 -33902
rect -64517 -34198 -64513 -33902
rect -65137 -34202 -64513 -34198
rect -64477 -33902 -64173 -33898
rect -64477 -34198 -64473 -33902
rect -64473 -34198 -64177 -33902
rect -64177 -34198 -64173 -33902
rect -64477 -34202 -64173 -34198
rect -64137 -33902 -63513 -33898
rect -64137 -34198 -64133 -33902
rect -64133 -34198 -63517 -33902
rect -63517 -34198 -63513 -33902
rect -64137 -34202 -63513 -34198
rect -63477 -33902 -63173 -33898
rect -63477 -34198 -63473 -33902
rect -63473 -34198 -63177 -33902
rect -63177 -34198 -63173 -33902
rect -63477 -34202 -63173 -34198
rect -63137 -33902 -62513 -33898
rect -63137 -34198 -63133 -33902
rect -63133 -34198 -62517 -33902
rect -62517 -34198 -62513 -33902
rect -63137 -34202 -62513 -34198
rect -62477 -33902 -62173 -33898
rect -62477 -34198 -62473 -33902
rect -62473 -34198 -62177 -33902
rect -62177 -34198 -62173 -33902
rect -62477 -34202 -62173 -34198
rect -62137 -33902 -61513 -33898
rect -62137 -34198 -62133 -33902
rect -62133 -34198 -61517 -33902
rect -61517 -34198 -61513 -33902
rect -62137 -34202 -61513 -34198
rect -61477 -33902 -61173 -33898
rect -61477 -34198 -61473 -33902
rect -61473 -34198 -61177 -33902
rect -61177 -34198 -61173 -33902
rect -61477 -34202 -61173 -34198
rect -61137 -33902 -60513 -33898
rect -61137 -34198 -61133 -33902
rect -61133 -34198 -60517 -33902
rect -60517 -34198 -60513 -33902
rect -61137 -34202 -60513 -34198
rect -60477 -33902 -60173 -33898
rect -60477 -34198 -60473 -33902
rect -60473 -34198 -60177 -33902
rect -60177 -34198 -60173 -33902
rect -60477 -34202 -60173 -34198
rect -60137 -33902 -59513 -33898
rect -60137 -34198 -60133 -33902
rect -60133 -34198 -59517 -33902
rect -59517 -34198 -59513 -33902
rect -60137 -34202 -59513 -34198
rect -59477 -33902 -59173 -33898
rect -59477 -34198 -59473 -33902
rect -59473 -34198 -59177 -33902
rect -59177 -34198 -59173 -33902
rect -59477 -34202 -59173 -34198
rect -59137 -33902 -58513 -33898
rect -59137 -34198 -59133 -33902
rect -59133 -34198 -58517 -33902
rect -58517 -34198 -58513 -33902
rect -59137 -34202 -58513 -34198
rect -58477 -33902 -58173 -33898
rect -58477 -34198 -58473 -33902
rect -58473 -34198 -58177 -33902
rect -58177 -34198 -58173 -33902
rect -58477 -34202 -58173 -34198
rect -58137 -33902 -57513 -33898
rect -58137 -34198 -58133 -33902
rect -58133 -34198 -57517 -33902
rect -57517 -34198 -57513 -33902
rect -58137 -34202 -57513 -34198
rect -57477 -33902 -57173 -33898
rect -57477 -34198 -57473 -33902
rect -57473 -34198 -57177 -33902
rect -57177 -34198 -57173 -33902
rect -57477 -34202 -57173 -34198
rect -57137 -33902 -56513 -33898
rect -57137 -34198 -57133 -33902
rect -57133 -34198 -56517 -33902
rect -56517 -34198 -56513 -33902
rect -57137 -34202 -56513 -34198
rect -56477 -33902 -56173 -33898
rect -56477 -34198 -56473 -33902
rect -56473 -34198 -56177 -33902
rect -56177 -34198 -56173 -33902
rect -56477 -34202 -56173 -34198
rect -56137 -33902 -55513 -33898
rect -56137 -34198 -56133 -33902
rect -56133 -34198 -55517 -33902
rect -55517 -34198 -55513 -33902
rect -56137 -34202 -55513 -34198
rect -55477 -33902 -55173 -33898
rect -55477 -34198 -55473 -33902
rect -55473 -34198 -55177 -33902
rect -55177 -34198 -55173 -33902
rect -55477 -34202 -55173 -34198
rect -55137 -33902 -54513 -33898
rect -55137 -34198 -55133 -33902
rect -55133 -34198 -54517 -33902
rect -54517 -34198 -54513 -33902
rect -55137 -34202 -54513 -34198
rect -54477 -33902 -54173 -33898
rect -54477 -34198 -54473 -33902
rect -54473 -34198 -54177 -33902
rect -54177 -34198 -54173 -33902
rect -54477 -34202 -54173 -34198
rect -54137 -33902 -53513 -33898
rect -54137 -34198 -54133 -33902
rect -54133 -34198 -53517 -33902
rect -53517 -34198 -53513 -33902
rect -54137 -34202 -53513 -34198
rect -53477 -33902 -53173 -33898
rect -53477 -34198 -53473 -33902
rect -53473 -34198 -53177 -33902
rect -53177 -34198 -53173 -33902
rect -53477 -34202 -53173 -34198
rect -53137 -33902 -52513 -33898
rect -53137 -34198 -53133 -33902
rect -53133 -34198 -52517 -33902
rect -52517 -34198 -52513 -33902
rect -53137 -34202 -52513 -34198
rect -52477 -33902 -52173 -33898
rect -52477 -34198 -52473 -33902
rect -52473 -34198 -52177 -33902
rect -52177 -34198 -52173 -33902
rect -52477 -34202 -52173 -34198
rect -52137 -33902 -51513 -33898
rect -52137 -34198 -52133 -33902
rect -52133 -34198 -51517 -33902
rect -51517 -34198 -51513 -33902
rect -52137 -34202 -51513 -34198
rect -51477 -33902 -51173 -33898
rect -51477 -34198 -51473 -33902
rect -51473 -34198 -51177 -33902
rect -51177 -34198 -51173 -33902
rect -51477 -34202 -51173 -34198
rect -51137 -33902 -50513 -33898
rect -51137 -34198 -51133 -33902
rect -51133 -34198 -50517 -33902
rect -50517 -34198 -50513 -33902
rect -51137 -34202 -50513 -34198
rect -50477 -33902 -50173 -33898
rect -50477 -34198 -50473 -33902
rect -50473 -34198 -50177 -33902
rect -50177 -34198 -50173 -33902
rect -50477 -34202 -50173 -34198
rect -50137 -33902 -49513 -33898
rect -50137 -34198 -50133 -33902
rect -50133 -34198 -49517 -33902
rect -49517 -34198 -49513 -33902
rect -50137 -34202 -49513 -34198
rect -49477 -33902 -49173 -33898
rect -49477 -34198 -49473 -33902
rect -49473 -34198 -49177 -33902
rect -49177 -34198 -49173 -33902
rect -49477 -34202 -49173 -34198
rect -49137 -33902 -48833 -33898
rect -49137 -34198 -49133 -33902
rect -49133 -34198 -48837 -33902
rect -48837 -34198 -48833 -33902
rect -49137 -34202 -48833 -34198
rect -74477 -34242 -74173 -34238
rect -74477 -34858 -74473 -34242
rect -74473 -34858 -74177 -34242
rect -74177 -34858 -74173 -34242
rect -74477 -34862 -74173 -34858
rect -73477 -34242 -73173 -34238
rect -73477 -34858 -73473 -34242
rect -73473 -34858 -73177 -34242
rect -73177 -34858 -73173 -34242
rect -73477 -34862 -73173 -34858
rect -72477 -34242 -72173 -34238
rect -72477 -34858 -72473 -34242
rect -72473 -34858 -72177 -34242
rect -72177 -34858 -72173 -34242
rect -72477 -34862 -72173 -34858
rect -71477 -34242 -71173 -34238
rect -71477 -34858 -71473 -34242
rect -71473 -34858 -71177 -34242
rect -71177 -34858 -71173 -34242
rect -71477 -34862 -71173 -34858
rect -70477 -34242 -70173 -34238
rect -70477 -34858 -70473 -34242
rect -70473 -34858 -70177 -34242
rect -70177 -34858 -70173 -34242
rect -70477 -34862 -70173 -34858
rect -69477 -34242 -69173 -34238
rect -69477 -34858 -69473 -34242
rect -69473 -34858 -69177 -34242
rect -69177 -34858 -69173 -34242
rect -69477 -34862 -69173 -34858
rect -68477 -34242 -68173 -34238
rect -68477 -34858 -68473 -34242
rect -68473 -34858 -68177 -34242
rect -68177 -34858 -68173 -34242
rect -68477 -34862 -68173 -34858
rect -67477 -34242 -67173 -34238
rect -67477 -34858 -67473 -34242
rect -67473 -34858 -67177 -34242
rect -67177 -34858 -67173 -34242
rect -67477 -34862 -67173 -34858
rect -66477 -34242 -66173 -34238
rect -66477 -34858 -66473 -34242
rect -66473 -34858 -66177 -34242
rect -66177 -34858 -66173 -34242
rect -66477 -34862 -66173 -34858
rect -65477 -34242 -65173 -34238
rect -65477 -34858 -65473 -34242
rect -65473 -34858 -65177 -34242
rect -65177 -34858 -65173 -34242
rect -65477 -34862 -65173 -34858
rect -64477 -34242 -64173 -34238
rect -64477 -34858 -64473 -34242
rect -64473 -34858 -64177 -34242
rect -64177 -34858 -64173 -34242
rect -64477 -34862 -64173 -34858
rect -63477 -34242 -63173 -34238
rect -63477 -34858 -63473 -34242
rect -63473 -34858 -63177 -34242
rect -63177 -34858 -63173 -34242
rect -63477 -34862 -63173 -34858
rect -62477 -34242 -62173 -34238
rect -62477 -34858 -62473 -34242
rect -62473 -34858 -62177 -34242
rect -62177 -34858 -62173 -34242
rect -62477 -34862 -62173 -34858
rect -61477 -34242 -61173 -34238
rect -61477 -34858 -61473 -34242
rect -61473 -34858 -61177 -34242
rect -61177 -34858 -61173 -34242
rect -61477 -34862 -61173 -34858
rect -60477 -34242 -60173 -34238
rect -60477 -34858 -60473 -34242
rect -60473 -34858 -60177 -34242
rect -60177 -34858 -60173 -34242
rect -60477 -34862 -60173 -34858
rect -59477 -34242 -59173 -34238
rect -59477 -34858 -59473 -34242
rect -59473 -34858 -59177 -34242
rect -59177 -34858 -59173 -34242
rect -59477 -34862 -59173 -34858
rect -58477 -34242 -58173 -34238
rect -58477 -34858 -58473 -34242
rect -58473 -34858 -58177 -34242
rect -58177 -34858 -58173 -34242
rect -58477 -34862 -58173 -34858
rect -57477 -34242 -57173 -34238
rect -57477 -34858 -57473 -34242
rect -57473 -34858 -57177 -34242
rect -57177 -34858 -57173 -34242
rect -57477 -34862 -57173 -34858
rect -56477 -34242 -56173 -34238
rect -56477 -34858 -56473 -34242
rect -56473 -34858 -56177 -34242
rect -56177 -34858 -56173 -34242
rect -56477 -34862 -56173 -34858
rect -55477 -34242 -55173 -34238
rect -55477 -34858 -55473 -34242
rect -55473 -34858 -55177 -34242
rect -55177 -34858 -55173 -34242
rect -55477 -34862 -55173 -34858
rect -54477 -34242 -54173 -34238
rect -54477 -34858 -54473 -34242
rect -54473 -34858 -54177 -34242
rect -54177 -34858 -54173 -34242
rect -54477 -34862 -54173 -34858
rect -53477 -34242 -53173 -34238
rect -53477 -34858 -53473 -34242
rect -53473 -34858 -53177 -34242
rect -53177 -34858 -53173 -34242
rect -53477 -34862 -53173 -34858
rect -52477 -34242 -52173 -34238
rect -52477 -34858 -52473 -34242
rect -52473 -34858 -52177 -34242
rect -52177 -34858 -52173 -34242
rect -52477 -34862 -52173 -34858
rect -51477 -34242 -51173 -34238
rect -51477 -34858 -51473 -34242
rect -51473 -34858 -51177 -34242
rect -51177 -34858 -51173 -34242
rect -51477 -34862 -51173 -34858
rect -50477 -34242 -50173 -34238
rect -50477 -34858 -50473 -34242
rect -50473 -34858 -50177 -34242
rect -50177 -34858 -50173 -34242
rect -50477 -34862 -50173 -34858
rect -49477 -34242 -49173 -34238
rect -49477 -34858 -49473 -34242
rect -49473 -34858 -49177 -34242
rect -49177 -34858 -49173 -34242
rect -49477 -34862 -49173 -34858
rect -74817 -34902 -74513 -34898
rect -74817 -35198 -74813 -34902
rect -74813 -35198 -74517 -34902
rect -74517 -35198 -74513 -34902
rect -74817 -35202 -74513 -35198
rect -74477 -34902 -74173 -34898
rect -74477 -35198 -74473 -34902
rect -74473 -35198 -74177 -34902
rect -74177 -35198 -74173 -34902
rect -74477 -35202 -74173 -35198
rect -74137 -34902 -73513 -34898
rect -74137 -35198 -74133 -34902
rect -74133 -35198 -73517 -34902
rect -73517 -35198 -73513 -34902
rect -74137 -35202 -73513 -35198
rect -73477 -34902 -73173 -34898
rect -73477 -35198 -73473 -34902
rect -73473 -35198 -73177 -34902
rect -73177 -35198 -73173 -34902
rect -73477 -35202 -73173 -35198
rect -73137 -34902 -72513 -34898
rect -73137 -35198 -73133 -34902
rect -73133 -35198 -72517 -34902
rect -72517 -35198 -72513 -34902
rect -73137 -35202 -72513 -35198
rect -72477 -34902 -72173 -34898
rect -72477 -35198 -72473 -34902
rect -72473 -35198 -72177 -34902
rect -72177 -35198 -72173 -34902
rect -72477 -35202 -72173 -35198
rect -72137 -34902 -71513 -34898
rect -72137 -35198 -72133 -34902
rect -72133 -35198 -71517 -34902
rect -71517 -35198 -71513 -34902
rect -72137 -35202 -71513 -35198
rect -71477 -34902 -71173 -34898
rect -71477 -35198 -71473 -34902
rect -71473 -35198 -71177 -34902
rect -71177 -35198 -71173 -34902
rect -71477 -35202 -71173 -35198
rect -71137 -34902 -70513 -34898
rect -71137 -35198 -71133 -34902
rect -71133 -35198 -70517 -34902
rect -70517 -35198 -70513 -34902
rect -71137 -35202 -70513 -35198
rect -70477 -34902 -70173 -34898
rect -70477 -35198 -70473 -34902
rect -70473 -35198 -70177 -34902
rect -70177 -35198 -70173 -34902
rect -70477 -35202 -70173 -35198
rect -70137 -34902 -69513 -34898
rect -70137 -35198 -70133 -34902
rect -70133 -35198 -69517 -34902
rect -69517 -35198 -69513 -34902
rect -70137 -35202 -69513 -35198
rect -69477 -34902 -69173 -34898
rect -69477 -35198 -69473 -34902
rect -69473 -35198 -69177 -34902
rect -69177 -35198 -69173 -34902
rect -69477 -35202 -69173 -35198
rect -69137 -34902 -68513 -34898
rect -69137 -35198 -69133 -34902
rect -69133 -35198 -68517 -34902
rect -68517 -35198 -68513 -34902
rect -69137 -35202 -68513 -35198
rect -68477 -34902 -68173 -34898
rect -68477 -35198 -68473 -34902
rect -68473 -35198 -68177 -34902
rect -68177 -35198 -68173 -34902
rect -68477 -35202 -68173 -35198
rect -68137 -34902 -67513 -34898
rect -68137 -35198 -68133 -34902
rect -68133 -35198 -67517 -34902
rect -67517 -35198 -67513 -34902
rect -68137 -35202 -67513 -35198
rect -67477 -34902 -67173 -34898
rect -67477 -35198 -67473 -34902
rect -67473 -35198 -67177 -34902
rect -67177 -35198 -67173 -34902
rect -67477 -35202 -67173 -35198
rect -67137 -34902 -66513 -34898
rect -67137 -35198 -67133 -34902
rect -67133 -35198 -66517 -34902
rect -66517 -35198 -66513 -34902
rect -67137 -35202 -66513 -35198
rect -66477 -34902 -66173 -34898
rect -66477 -35198 -66473 -34902
rect -66473 -35198 -66177 -34902
rect -66177 -35198 -66173 -34902
rect -66477 -35202 -66173 -35198
rect -66137 -34902 -65513 -34898
rect -66137 -35198 -66133 -34902
rect -66133 -35198 -65517 -34902
rect -65517 -35198 -65513 -34902
rect -66137 -35202 -65513 -35198
rect -65477 -34902 -65173 -34898
rect -65477 -35198 -65473 -34902
rect -65473 -35198 -65177 -34902
rect -65177 -35198 -65173 -34902
rect -65477 -35202 -65173 -35198
rect -65137 -34902 -64513 -34898
rect -65137 -35198 -65133 -34902
rect -65133 -35198 -64517 -34902
rect -64517 -35198 -64513 -34902
rect -65137 -35202 -64513 -35198
rect -64477 -34902 -64173 -34898
rect -64477 -35198 -64473 -34902
rect -64473 -35198 -64177 -34902
rect -64177 -35198 -64173 -34902
rect -64477 -35202 -64173 -35198
rect -64137 -34902 -63513 -34898
rect -64137 -35198 -64133 -34902
rect -64133 -35198 -63517 -34902
rect -63517 -35198 -63513 -34902
rect -64137 -35202 -63513 -35198
rect -63477 -34902 -63173 -34898
rect -63477 -35198 -63473 -34902
rect -63473 -35198 -63177 -34902
rect -63177 -35198 -63173 -34902
rect -63477 -35202 -63173 -35198
rect -63137 -34902 -62513 -34898
rect -63137 -35198 -63133 -34902
rect -63133 -35198 -62517 -34902
rect -62517 -35198 -62513 -34902
rect -63137 -35202 -62513 -35198
rect -62477 -34902 -62173 -34898
rect -62477 -35198 -62473 -34902
rect -62473 -35198 -62177 -34902
rect -62177 -35198 -62173 -34902
rect -62477 -35202 -62173 -35198
rect -62137 -34902 -61513 -34898
rect -62137 -35198 -62133 -34902
rect -62133 -35198 -61517 -34902
rect -61517 -35198 -61513 -34902
rect -62137 -35202 -61513 -35198
rect -61477 -34902 -61173 -34898
rect -61477 -35198 -61473 -34902
rect -61473 -35198 -61177 -34902
rect -61177 -35198 -61173 -34902
rect -61477 -35202 -61173 -35198
rect -61137 -34902 -60513 -34898
rect -61137 -35198 -61133 -34902
rect -61133 -35198 -60517 -34902
rect -60517 -35198 -60513 -34902
rect -61137 -35202 -60513 -35198
rect -60477 -34902 -60173 -34898
rect -60477 -35198 -60473 -34902
rect -60473 -35198 -60177 -34902
rect -60177 -35198 -60173 -34902
rect -60477 -35202 -60173 -35198
rect -60137 -34902 -59513 -34898
rect -60137 -35198 -60133 -34902
rect -60133 -35198 -59517 -34902
rect -59517 -35198 -59513 -34902
rect -60137 -35202 -59513 -35198
rect -59477 -34902 -59173 -34898
rect -59477 -35198 -59473 -34902
rect -59473 -35198 -59177 -34902
rect -59177 -35198 -59173 -34902
rect -59477 -35202 -59173 -35198
rect -59137 -34902 -58513 -34898
rect -59137 -35198 -59133 -34902
rect -59133 -35198 -58517 -34902
rect -58517 -35198 -58513 -34902
rect -59137 -35202 -58513 -35198
rect -58477 -34902 -58173 -34898
rect -58477 -35198 -58473 -34902
rect -58473 -35198 -58177 -34902
rect -58177 -35198 -58173 -34902
rect -58477 -35202 -58173 -35198
rect -58137 -34902 -57513 -34898
rect -58137 -35198 -58133 -34902
rect -58133 -35198 -57517 -34902
rect -57517 -35198 -57513 -34902
rect -58137 -35202 -57513 -35198
rect -57477 -34902 -57173 -34898
rect -57477 -35198 -57473 -34902
rect -57473 -35198 -57177 -34902
rect -57177 -35198 -57173 -34902
rect -57477 -35202 -57173 -35198
rect -57137 -34902 -56513 -34898
rect -57137 -35198 -57133 -34902
rect -57133 -35198 -56517 -34902
rect -56517 -35198 -56513 -34902
rect -57137 -35202 -56513 -35198
rect -56477 -34902 -56173 -34898
rect -56477 -35198 -56473 -34902
rect -56473 -35198 -56177 -34902
rect -56177 -35198 -56173 -34902
rect -56477 -35202 -56173 -35198
rect -56137 -34902 -55513 -34898
rect -56137 -35198 -56133 -34902
rect -56133 -35198 -55517 -34902
rect -55517 -35198 -55513 -34902
rect -56137 -35202 -55513 -35198
rect -55477 -34902 -55173 -34898
rect -55477 -35198 -55473 -34902
rect -55473 -35198 -55177 -34902
rect -55177 -35198 -55173 -34902
rect -55477 -35202 -55173 -35198
rect -55137 -34902 -54513 -34898
rect -55137 -35198 -55133 -34902
rect -55133 -35198 -54517 -34902
rect -54517 -35198 -54513 -34902
rect -55137 -35202 -54513 -35198
rect -54477 -34902 -54173 -34898
rect -54477 -35198 -54473 -34902
rect -54473 -35198 -54177 -34902
rect -54177 -35198 -54173 -34902
rect -54477 -35202 -54173 -35198
rect -54137 -34902 -53513 -34898
rect -54137 -35198 -54133 -34902
rect -54133 -35198 -53517 -34902
rect -53517 -35198 -53513 -34902
rect -54137 -35202 -53513 -35198
rect -53477 -34902 -53173 -34898
rect -53477 -35198 -53473 -34902
rect -53473 -35198 -53177 -34902
rect -53177 -35198 -53173 -34902
rect -53477 -35202 -53173 -35198
rect -53137 -34902 -52513 -34898
rect -53137 -35198 -53133 -34902
rect -53133 -35198 -52517 -34902
rect -52517 -35198 -52513 -34902
rect -53137 -35202 -52513 -35198
rect -52477 -34902 -52173 -34898
rect -52477 -35198 -52473 -34902
rect -52473 -35198 -52177 -34902
rect -52177 -35198 -52173 -34902
rect -52477 -35202 -52173 -35198
rect -52137 -34902 -51513 -34898
rect -52137 -35198 -52133 -34902
rect -52133 -35198 -51517 -34902
rect -51517 -35198 -51513 -34902
rect -52137 -35202 -51513 -35198
rect -51477 -34902 -51173 -34898
rect -51477 -35198 -51473 -34902
rect -51473 -35198 -51177 -34902
rect -51177 -35198 -51173 -34902
rect -51477 -35202 -51173 -35198
rect -51137 -34902 -50513 -34898
rect -51137 -35198 -51133 -34902
rect -51133 -35198 -50517 -34902
rect -50517 -35198 -50513 -34902
rect -51137 -35202 -50513 -35198
rect -50477 -34902 -50173 -34898
rect -50477 -35198 -50473 -34902
rect -50473 -35198 -50177 -34902
rect -50177 -35198 -50173 -34902
rect -50477 -35202 -50173 -35198
rect -50137 -34902 -49513 -34898
rect -50137 -35198 -50133 -34902
rect -50133 -35198 -49517 -34902
rect -49517 -35198 -49513 -34902
rect -50137 -35202 -49513 -35198
rect -49477 -34902 -49173 -34898
rect -49477 -35198 -49473 -34902
rect -49473 -35198 -49177 -34902
rect -49177 -35198 -49173 -34902
rect -49477 -35202 -49173 -35198
rect -49137 -34902 -48833 -34898
rect -49137 -35198 -49133 -34902
rect -49133 -35198 -48837 -34902
rect -48837 -35198 -48833 -34902
rect -49137 -35202 -48833 -35198
rect -74477 -35242 -74173 -35238
rect -74477 -35858 -74473 -35242
rect -74473 -35858 -74177 -35242
rect -74177 -35858 -74173 -35242
rect -74477 -35862 -74173 -35858
rect -73477 -35242 -73173 -35238
rect -73477 -35858 -73473 -35242
rect -73473 -35858 -73177 -35242
rect -73177 -35858 -73173 -35242
rect -73477 -35862 -73173 -35858
rect -72477 -35242 -72173 -35238
rect -72477 -35858 -72473 -35242
rect -72473 -35858 -72177 -35242
rect -72177 -35858 -72173 -35242
rect -72477 -35862 -72173 -35858
rect -71477 -35242 -71173 -35238
rect -71477 -35858 -71473 -35242
rect -71473 -35858 -71177 -35242
rect -71177 -35858 -71173 -35242
rect -71477 -35862 -71173 -35858
rect -70477 -35242 -70173 -35238
rect -70477 -35858 -70473 -35242
rect -70473 -35858 -70177 -35242
rect -70177 -35858 -70173 -35242
rect -70477 -35862 -70173 -35858
rect -69477 -35242 -69173 -35238
rect -69477 -35858 -69473 -35242
rect -69473 -35858 -69177 -35242
rect -69177 -35858 -69173 -35242
rect -69477 -35862 -69173 -35858
rect -68477 -35242 -68173 -35238
rect -68477 -35858 -68473 -35242
rect -68473 -35858 -68177 -35242
rect -68177 -35858 -68173 -35242
rect -68477 -35862 -68173 -35858
rect -67477 -35242 -67173 -35238
rect -67477 -35858 -67473 -35242
rect -67473 -35858 -67177 -35242
rect -67177 -35858 -67173 -35242
rect -67477 -35862 -67173 -35858
rect -66477 -35242 -66173 -35238
rect -66477 -35858 -66473 -35242
rect -66473 -35858 -66177 -35242
rect -66177 -35858 -66173 -35242
rect -66477 -35862 -66173 -35858
rect -65477 -35242 -65173 -35238
rect -65477 -35858 -65473 -35242
rect -65473 -35858 -65177 -35242
rect -65177 -35858 -65173 -35242
rect -65477 -35862 -65173 -35858
rect -64477 -35242 -64173 -35238
rect -64477 -35858 -64473 -35242
rect -64473 -35858 -64177 -35242
rect -64177 -35858 -64173 -35242
rect -64477 -35862 -64173 -35858
rect -63477 -35242 -63173 -35238
rect -63477 -35858 -63473 -35242
rect -63473 -35858 -63177 -35242
rect -63177 -35858 -63173 -35242
rect -63477 -35862 -63173 -35858
rect -62477 -35242 -62173 -35238
rect -62477 -35858 -62473 -35242
rect -62473 -35858 -62177 -35242
rect -62177 -35858 -62173 -35242
rect -62477 -35862 -62173 -35858
rect -61477 -35242 -61173 -35238
rect -61477 -35858 -61473 -35242
rect -61473 -35858 -61177 -35242
rect -61177 -35858 -61173 -35242
rect -61477 -35862 -61173 -35858
rect -60477 -35242 -60173 -35238
rect -60477 -35858 -60473 -35242
rect -60473 -35858 -60177 -35242
rect -60177 -35858 -60173 -35242
rect -60477 -35862 -60173 -35858
rect -59477 -35242 -59173 -35238
rect -59477 -35858 -59473 -35242
rect -59473 -35858 -59177 -35242
rect -59177 -35858 -59173 -35242
rect -59477 -35862 -59173 -35858
rect -58477 -35242 -58173 -35238
rect -58477 -35858 -58473 -35242
rect -58473 -35858 -58177 -35242
rect -58177 -35858 -58173 -35242
rect -58477 -35862 -58173 -35858
rect -57477 -35242 -57173 -35238
rect -57477 -35858 -57473 -35242
rect -57473 -35858 -57177 -35242
rect -57177 -35858 -57173 -35242
rect -57477 -35862 -57173 -35858
rect -56477 -35242 -56173 -35238
rect -56477 -35858 -56473 -35242
rect -56473 -35858 -56177 -35242
rect -56177 -35858 -56173 -35242
rect -56477 -35862 -56173 -35858
rect -55477 -35242 -55173 -35238
rect -55477 -35858 -55473 -35242
rect -55473 -35858 -55177 -35242
rect -55177 -35858 -55173 -35242
rect -55477 -35862 -55173 -35858
rect -54477 -35242 -54173 -35238
rect -54477 -35858 -54473 -35242
rect -54473 -35858 -54177 -35242
rect -54177 -35858 -54173 -35242
rect -54477 -35862 -54173 -35858
rect -53477 -35242 -53173 -35238
rect -53477 -35858 -53473 -35242
rect -53473 -35858 -53177 -35242
rect -53177 -35858 -53173 -35242
rect -53477 -35862 -53173 -35858
rect -52477 -35242 -52173 -35238
rect -52477 -35858 -52473 -35242
rect -52473 -35858 -52177 -35242
rect -52177 -35858 -52173 -35242
rect -52477 -35862 -52173 -35858
rect -51477 -35242 -51173 -35238
rect -51477 -35858 -51473 -35242
rect -51473 -35858 -51177 -35242
rect -51177 -35858 -51173 -35242
rect -51477 -35862 -51173 -35858
rect -50477 -35242 -50173 -35238
rect -50477 -35858 -50473 -35242
rect -50473 -35858 -50177 -35242
rect -50177 -35858 -50173 -35242
rect -50477 -35862 -50173 -35858
rect -49477 -35242 -49173 -35238
rect -49477 -35858 -49473 -35242
rect -49473 -35858 -49177 -35242
rect -49177 -35858 -49173 -35242
rect -49477 -35862 -49173 -35858
rect -74817 -35902 -74513 -35898
rect -74817 -36198 -74813 -35902
rect -74813 -36198 -74517 -35902
rect -74517 -36198 -74513 -35902
rect -74817 -36202 -74513 -36198
rect -74477 -35902 -74173 -35898
rect -74477 -36198 -74473 -35902
rect -74473 -36198 -74177 -35902
rect -74177 -36198 -74173 -35902
rect -74477 -36202 -74173 -36198
rect -74137 -35902 -73513 -35898
rect -74137 -36198 -74133 -35902
rect -74133 -36198 -73517 -35902
rect -73517 -36198 -73513 -35902
rect -74137 -36202 -73513 -36198
rect -73477 -35902 -73173 -35898
rect -73477 -36198 -73473 -35902
rect -73473 -36198 -73177 -35902
rect -73177 -36198 -73173 -35902
rect -73477 -36202 -73173 -36198
rect -73137 -35902 -72513 -35898
rect -73137 -36198 -73133 -35902
rect -73133 -36198 -72517 -35902
rect -72517 -36198 -72513 -35902
rect -73137 -36202 -72513 -36198
rect -72477 -35902 -72173 -35898
rect -72477 -36198 -72473 -35902
rect -72473 -36198 -72177 -35902
rect -72177 -36198 -72173 -35902
rect -72477 -36202 -72173 -36198
rect -72137 -35902 -71513 -35898
rect -72137 -36198 -72133 -35902
rect -72133 -36198 -71517 -35902
rect -71517 -36198 -71513 -35902
rect -72137 -36202 -71513 -36198
rect -71477 -35902 -71173 -35898
rect -71477 -36198 -71473 -35902
rect -71473 -36198 -71177 -35902
rect -71177 -36198 -71173 -35902
rect -71477 -36202 -71173 -36198
rect -71137 -35902 -70513 -35898
rect -71137 -36198 -71133 -35902
rect -71133 -36198 -70517 -35902
rect -70517 -36198 -70513 -35902
rect -71137 -36202 -70513 -36198
rect -70477 -35902 -70173 -35898
rect -70477 -36198 -70473 -35902
rect -70473 -36198 -70177 -35902
rect -70177 -36198 -70173 -35902
rect -70477 -36202 -70173 -36198
rect -70137 -35902 -69513 -35898
rect -70137 -36198 -70133 -35902
rect -70133 -36198 -69517 -35902
rect -69517 -36198 -69513 -35902
rect -70137 -36202 -69513 -36198
rect -69477 -35902 -69173 -35898
rect -69477 -36198 -69473 -35902
rect -69473 -36198 -69177 -35902
rect -69177 -36198 -69173 -35902
rect -69477 -36202 -69173 -36198
rect -69137 -35902 -68513 -35898
rect -69137 -36198 -69133 -35902
rect -69133 -36198 -68517 -35902
rect -68517 -36198 -68513 -35902
rect -69137 -36202 -68513 -36198
rect -68477 -35902 -68173 -35898
rect -68477 -36198 -68473 -35902
rect -68473 -36198 -68177 -35902
rect -68177 -36198 -68173 -35902
rect -68477 -36202 -68173 -36198
rect -68137 -35902 -67513 -35898
rect -68137 -36198 -68133 -35902
rect -68133 -36198 -67517 -35902
rect -67517 -36198 -67513 -35902
rect -68137 -36202 -67513 -36198
rect -67477 -35902 -67173 -35898
rect -67477 -36198 -67473 -35902
rect -67473 -36198 -67177 -35902
rect -67177 -36198 -67173 -35902
rect -67477 -36202 -67173 -36198
rect -67137 -35902 -66513 -35898
rect -67137 -36198 -67133 -35902
rect -67133 -36198 -66517 -35902
rect -66517 -36198 -66513 -35902
rect -67137 -36202 -66513 -36198
rect -66477 -35902 -66173 -35898
rect -66477 -36198 -66473 -35902
rect -66473 -36198 -66177 -35902
rect -66177 -36198 -66173 -35902
rect -66477 -36202 -66173 -36198
rect -66137 -35902 -65513 -35898
rect -66137 -36198 -66133 -35902
rect -66133 -36198 -65517 -35902
rect -65517 -36198 -65513 -35902
rect -66137 -36202 -65513 -36198
rect -65477 -35902 -65173 -35898
rect -65477 -36198 -65473 -35902
rect -65473 -36198 -65177 -35902
rect -65177 -36198 -65173 -35902
rect -65477 -36202 -65173 -36198
rect -65137 -35902 -64513 -35898
rect -65137 -36198 -65133 -35902
rect -65133 -36198 -64517 -35902
rect -64517 -36198 -64513 -35902
rect -65137 -36202 -64513 -36198
rect -64477 -35902 -64173 -35898
rect -64477 -36198 -64473 -35902
rect -64473 -36198 -64177 -35902
rect -64177 -36198 -64173 -35902
rect -64477 -36202 -64173 -36198
rect -64137 -35902 -63513 -35898
rect -64137 -36198 -64133 -35902
rect -64133 -36198 -63517 -35902
rect -63517 -36198 -63513 -35902
rect -64137 -36202 -63513 -36198
rect -63477 -35902 -63173 -35898
rect -63477 -36198 -63473 -35902
rect -63473 -36198 -63177 -35902
rect -63177 -36198 -63173 -35902
rect -63477 -36202 -63173 -36198
rect -63137 -35902 -62513 -35898
rect -63137 -36198 -63133 -35902
rect -63133 -36198 -62517 -35902
rect -62517 -36198 -62513 -35902
rect -63137 -36202 -62513 -36198
rect -62477 -35902 -62173 -35898
rect -62477 -36198 -62473 -35902
rect -62473 -36198 -62177 -35902
rect -62177 -36198 -62173 -35902
rect -62477 -36202 -62173 -36198
rect -62137 -35902 -61513 -35898
rect -62137 -36198 -62133 -35902
rect -62133 -36198 -61517 -35902
rect -61517 -36198 -61513 -35902
rect -62137 -36202 -61513 -36198
rect -61477 -35902 -61173 -35898
rect -61477 -36198 -61473 -35902
rect -61473 -36198 -61177 -35902
rect -61177 -36198 -61173 -35902
rect -61477 -36202 -61173 -36198
rect -61137 -35902 -60513 -35898
rect -61137 -36198 -61133 -35902
rect -61133 -36198 -60517 -35902
rect -60517 -36198 -60513 -35902
rect -61137 -36202 -60513 -36198
rect -60477 -35902 -60173 -35898
rect -60477 -36198 -60473 -35902
rect -60473 -36198 -60177 -35902
rect -60177 -36198 -60173 -35902
rect -60477 -36202 -60173 -36198
rect -60137 -35902 -59513 -35898
rect -60137 -36198 -60133 -35902
rect -60133 -36198 -59517 -35902
rect -59517 -36198 -59513 -35902
rect -60137 -36202 -59513 -36198
rect -59477 -35902 -59173 -35898
rect -59477 -36198 -59473 -35902
rect -59473 -36198 -59177 -35902
rect -59177 -36198 -59173 -35902
rect -59477 -36202 -59173 -36198
rect -59137 -35902 -58513 -35898
rect -59137 -36198 -59133 -35902
rect -59133 -36198 -58517 -35902
rect -58517 -36198 -58513 -35902
rect -59137 -36202 -58513 -36198
rect -58477 -35902 -58173 -35898
rect -58477 -36198 -58473 -35902
rect -58473 -36198 -58177 -35902
rect -58177 -36198 -58173 -35902
rect -58477 -36202 -58173 -36198
rect -58137 -35902 -57513 -35898
rect -58137 -36198 -58133 -35902
rect -58133 -36198 -57517 -35902
rect -57517 -36198 -57513 -35902
rect -58137 -36202 -57513 -36198
rect -57477 -35902 -57173 -35898
rect -57477 -36198 -57473 -35902
rect -57473 -36198 -57177 -35902
rect -57177 -36198 -57173 -35902
rect -57477 -36202 -57173 -36198
rect -57137 -35902 -56513 -35898
rect -57137 -36198 -57133 -35902
rect -57133 -36198 -56517 -35902
rect -56517 -36198 -56513 -35902
rect -57137 -36202 -56513 -36198
rect -56477 -35902 -56173 -35898
rect -56477 -36198 -56473 -35902
rect -56473 -36198 -56177 -35902
rect -56177 -36198 -56173 -35902
rect -56477 -36202 -56173 -36198
rect -56137 -35902 -55513 -35898
rect -56137 -36198 -56133 -35902
rect -56133 -36198 -55517 -35902
rect -55517 -36198 -55513 -35902
rect -56137 -36202 -55513 -36198
rect -55477 -35902 -55173 -35898
rect -55477 -36198 -55473 -35902
rect -55473 -36198 -55177 -35902
rect -55177 -36198 -55173 -35902
rect -55477 -36202 -55173 -36198
rect -55137 -35902 -54513 -35898
rect -55137 -36198 -55133 -35902
rect -55133 -36198 -54517 -35902
rect -54517 -36198 -54513 -35902
rect -55137 -36202 -54513 -36198
rect -54477 -35902 -54173 -35898
rect -54477 -36198 -54473 -35902
rect -54473 -36198 -54177 -35902
rect -54177 -36198 -54173 -35902
rect -54477 -36202 -54173 -36198
rect -54137 -35902 -53513 -35898
rect -54137 -36198 -54133 -35902
rect -54133 -36198 -53517 -35902
rect -53517 -36198 -53513 -35902
rect -54137 -36202 -53513 -36198
rect -53477 -35902 -53173 -35898
rect -53477 -36198 -53473 -35902
rect -53473 -36198 -53177 -35902
rect -53177 -36198 -53173 -35902
rect -53477 -36202 -53173 -36198
rect -53137 -35902 -52513 -35898
rect -53137 -36198 -53133 -35902
rect -53133 -36198 -52517 -35902
rect -52517 -36198 -52513 -35902
rect -53137 -36202 -52513 -36198
rect -52477 -35902 -52173 -35898
rect -52477 -36198 -52473 -35902
rect -52473 -36198 -52177 -35902
rect -52177 -36198 -52173 -35902
rect -52477 -36202 -52173 -36198
rect -52137 -35902 -51513 -35898
rect -52137 -36198 -52133 -35902
rect -52133 -36198 -51517 -35902
rect -51517 -36198 -51513 -35902
rect -52137 -36202 -51513 -36198
rect -51477 -35902 -51173 -35898
rect -51477 -36198 -51473 -35902
rect -51473 -36198 -51177 -35902
rect -51177 -36198 -51173 -35902
rect -51477 -36202 -51173 -36198
rect -51137 -35902 -50513 -35898
rect -51137 -36198 -51133 -35902
rect -51133 -36198 -50517 -35902
rect -50517 -36198 -50513 -35902
rect -51137 -36202 -50513 -36198
rect -50477 -35902 -50173 -35898
rect -50477 -36198 -50473 -35902
rect -50473 -36198 -50177 -35902
rect -50177 -36198 -50173 -35902
rect -50477 -36202 -50173 -36198
rect -50137 -35902 -49513 -35898
rect -50137 -36198 -50133 -35902
rect -50133 -36198 -49517 -35902
rect -49517 -36198 -49513 -35902
rect -50137 -36202 -49513 -36198
rect -49477 -35902 -49173 -35898
rect -49477 -36198 -49473 -35902
rect -49473 -36198 -49177 -35902
rect -49177 -36198 -49173 -35902
rect -49477 -36202 -49173 -36198
rect -49137 -35902 -48833 -35898
rect -49137 -36198 -49133 -35902
rect -49133 -36198 -48837 -35902
rect -48837 -36198 -48833 -35902
rect -49137 -36202 -48833 -36198
rect -74477 -36242 -74173 -36238
rect -74477 -36858 -74473 -36242
rect -74473 -36858 -74177 -36242
rect -74177 -36858 -74173 -36242
rect -74477 -36862 -74173 -36858
rect -73477 -36242 -73173 -36238
rect -73477 -36858 -73473 -36242
rect -73473 -36858 -73177 -36242
rect -73177 -36858 -73173 -36242
rect -73477 -36862 -73173 -36858
rect -72477 -36242 -72173 -36238
rect -72477 -36858 -72473 -36242
rect -72473 -36858 -72177 -36242
rect -72177 -36858 -72173 -36242
rect -72477 -36862 -72173 -36858
rect -71477 -36242 -71173 -36238
rect -71477 -36858 -71473 -36242
rect -71473 -36858 -71177 -36242
rect -71177 -36858 -71173 -36242
rect -71477 -36862 -71173 -36858
rect -70477 -36242 -70173 -36238
rect -70477 -36858 -70473 -36242
rect -70473 -36858 -70177 -36242
rect -70177 -36858 -70173 -36242
rect -70477 -36862 -70173 -36858
rect -69477 -36242 -69173 -36238
rect -69477 -36858 -69473 -36242
rect -69473 -36858 -69177 -36242
rect -69177 -36858 -69173 -36242
rect -69477 -36862 -69173 -36858
rect -68477 -36242 -68173 -36238
rect -68477 -36858 -68473 -36242
rect -68473 -36858 -68177 -36242
rect -68177 -36858 -68173 -36242
rect -68477 -36862 -68173 -36858
rect -67477 -36242 -67173 -36238
rect -67477 -36858 -67473 -36242
rect -67473 -36858 -67177 -36242
rect -67177 -36858 -67173 -36242
rect -67477 -36862 -67173 -36858
rect -66477 -36242 -66173 -36238
rect -66477 -36858 -66473 -36242
rect -66473 -36858 -66177 -36242
rect -66177 -36858 -66173 -36242
rect -66477 -36862 -66173 -36858
rect -65477 -36242 -65173 -36238
rect -65477 -36858 -65473 -36242
rect -65473 -36858 -65177 -36242
rect -65177 -36858 -65173 -36242
rect -65477 -36862 -65173 -36858
rect -64477 -36242 -64173 -36238
rect -64477 -36858 -64473 -36242
rect -64473 -36858 -64177 -36242
rect -64177 -36858 -64173 -36242
rect -64477 -36862 -64173 -36858
rect -63477 -36242 -63173 -36238
rect -63477 -36858 -63473 -36242
rect -63473 -36858 -63177 -36242
rect -63177 -36858 -63173 -36242
rect -63477 -36862 -63173 -36858
rect -62477 -36242 -62173 -36238
rect -62477 -36858 -62473 -36242
rect -62473 -36858 -62177 -36242
rect -62177 -36858 -62173 -36242
rect -62477 -36862 -62173 -36858
rect -61477 -36242 -61173 -36238
rect -61477 -36858 -61473 -36242
rect -61473 -36858 -61177 -36242
rect -61177 -36858 -61173 -36242
rect -61477 -36862 -61173 -36858
rect -60477 -36242 -60173 -36238
rect -60477 -36858 -60473 -36242
rect -60473 -36858 -60177 -36242
rect -60177 -36858 -60173 -36242
rect -60477 -36862 -60173 -36858
rect -59477 -36242 -59173 -36238
rect -59477 -36858 -59473 -36242
rect -59473 -36858 -59177 -36242
rect -59177 -36858 -59173 -36242
rect -59477 -36862 -59173 -36858
rect -58477 -36242 -58173 -36238
rect -58477 -36858 -58473 -36242
rect -58473 -36858 -58177 -36242
rect -58177 -36858 -58173 -36242
rect -58477 -36862 -58173 -36858
rect -57477 -36242 -57173 -36238
rect -57477 -36858 -57473 -36242
rect -57473 -36858 -57177 -36242
rect -57177 -36858 -57173 -36242
rect -57477 -36862 -57173 -36858
rect -56477 -36242 -56173 -36238
rect -56477 -36858 -56473 -36242
rect -56473 -36858 -56177 -36242
rect -56177 -36858 -56173 -36242
rect -56477 -36862 -56173 -36858
rect -55477 -36242 -55173 -36238
rect -55477 -36858 -55473 -36242
rect -55473 -36858 -55177 -36242
rect -55177 -36858 -55173 -36242
rect -55477 -36862 -55173 -36858
rect -54477 -36242 -54173 -36238
rect -54477 -36858 -54473 -36242
rect -54473 -36858 -54177 -36242
rect -54177 -36858 -54173 -36242
rect -54477 -36862 -54173 -36858
rect -53477 -36242 -53173 -36238
rect -53477 -36858 -53473 -36242
rect -53473 -36858 -53177 -36242
rect -53177 -36858 -53173 -36242
rect -53477 -36862 -53173 -36858
rect -52477 -36242 -52173 -36238
rect -52477 -36858 -52473 -36242
rect -52473 -36858 -52177 -36242
rect -52177 -36858 -52173 -36242
rect -52477 -36862 -52173 -36858
rect -51477 -36242 -51173 -36238
rect -51477 -36858 -51473 -36242
rect -51473 -36858 -51177 -36242
rect -51177 -36858 -51173 -36242
rect -51477 -36862 -51173 -36858
rect -50477 -36242 -50173 -36238
rect -50477 -36858 -50473 -36242
rect -50473 -36858 -50177 -36242
rect -50177 -36858 -50173 -36242
rect -50477 -36862 -50173 -36858
rect -49477 -36242 -49173 -36238
rect -49477 -36858 -49473 -36242
rect -49473 -36858 -49177 -36242
rect -49177 -36858 -49173 -36242
rect -49477 -36862 -49173 -36858
rect -74817 -36902 -74513 -36898
rect -74817 -37198 -74813 -36902
rect -74813 -37198 -74517 -36902
rect -74517 -37198 -74513 -36902
rect -74817 -37202 -74513 -37198
rect -74477 -36902 -74173 -36898
rect -74477 -37198 -74473 -36902
rect -74473 -37198 -74177 -36902
rect -74177 -37198 -74173 -36902
rect -74477 -37202 -74173 -37198
rect -74137 -36902 -73513 -36898
rect -74137 -37198 -74133 -36902
rect -74133 -37198 -73517 -36902
rect -73517 -37198 -73513 -36902
rect -74137 -37202 -73513 -37198
rect -73477 -36902 -73173 -36898
rect -73477 -37198 -73473 -36902
rect -73473 -37198 -73177 -36902
rect -73177 -37198 -73173 -36902
rect -73477 -37202 -73173 -37198
rect -73137 -36902 -72513 -36898
rect -73137 -37198 -73133 -36902
rect -73133 -37198 -72517 -36902
rect -72517 -37198 -72513 -36902
rect -73137 -37202 -72513 -37198
rect -72477 -36902 -72173 -36898
rect -72477 -37198 -72473 -36902
rect -72473 -37198 -72177 -36902
rect -72177 -37198 -72173 -36902
rect -72477 -37202 -72173 -37198
rect -72137 -36902 -71513 -36898
rect -72137 -37198 -72133 -36902
rect -72133 -37198 -71517 -36902
rect -71517 -37198 -71513 -36902
rect -72137 -37202 -71513 -37198
rect -71477 -36902 -71173 -36898
rect -71477 -37198 -71473 -36902
rect -71473 -37198 -71177 -36902
rect -71177 -37198 -71173 -36902
rect -71477 -37202 -71173 -37198
rect -71137 -36902 -70513 -36898
rect -71137 -37198 -71133 -36902
rect -71133 -37198 -70517 -36902
rect -70517 -37198 -70513 -36902
rect -71137 -37202 -70513 -37198
rect -70477 -36902 -70173 -36898
rect -70477 -37198 -70473 -36902
rect -70473 -37198 -70177 -36902
rect -70177 -37198 -70173 -36902
rect -70477 -37202 -70173 -37198
rect -70137 -36902 -69513 -36898
rect -70137 -37198 -70133 -36902
rect -70133 -37198 -69517 -36902
rect -69517 -37198 -69513 -36902
rect -70137 -37202 -69513 -37198
rect -69477 -36902 -69173 -36898
rect -69477 -37198 -69473 -36902
rect -69473 -37198 -69177 -36902
rect -69177 -37198 -69173 -36902
rect -69477 -37202 -69173 -37198
rect -69137 -36902 -68513 -36898
rect -69137 -37198 -69133 -36902
rect -69133 -37198 -68517 -36902
rect -68517 -37198 -68513 -36902
rect -69137 -37202 -68513 -37198
rect -68477 -36902 -68173 -36898
rect -68477 -37198 -68473 -36902
rect -68473 -37198 -68177 -36902
rect -68177 -37198 -68173 -36902
rect -68477 -37202 -68173 -37198
rect -68137 -36902 -67513 -36898
rect -68137 -37198 -68133 -36902
rect -68133 -37198 -67517 -36902
rect -67517 -37198 -67513 -36902
rect -68137 -37202 -67513 -37198
rect -67477 -36902 -67173 -36898
rect -67477 -37198 -67473 -36902
rect -67473 -37198 -67177 -36902
rect -67177 -37198 -67173 -36902
rect -67477 -37202 -67173 -37198
rect -67137 -36902 -66513 -36898
rect -67137 -37198 -67133 -36902
rect -67133 -37198 -66517 -36902
rect -66517 -37198 -66513 -36902
rect -67137 -37202 -66513 -37198
rect -66477 -36902 -66173 -36898
rect -66477 -37198 -66473 -36902
rect -66473 -37198 -66177 -36902
rect -66177 -37198 -66173 -36902
rect -66477 -37202 -66173 -37198
rect -66137 -36902 -65513 -36898
rect -66137 -37198 -66133 -36902
rect -66133 -37198 -65517 -36902
rect -65517 -37198 -65513 -36902
rect -66137 -37202 -65513 -37198
rect -65477 -36902 -65173 -36898
rect -65477 -37198 -65473 -36902
rect -65473 -37198 -65177 -36902
rect -65177 -37198 -65173 -36902
rect -65477 -37202 -65173 -37198
rect -65137 -36902 -64513 -36898
rect -65137 -37198 -65133 -36902
rect -65133 -37198 -64517 -36902
rect -64517 -37198 -64513 -36902
rect -65137 -37202 -64513 -37198
rect -64477 -36902 -64173 -36898
rect -64477 -37198 -64473 -36902
rect -64473 -37198 -64177 -36902
rect -64177 -37198 -64173 -36902
rect -64477 -37202 -64173 -37198
rect -64137 -36902 -63513 -36898
rect -64137 -37198 -64133 -36902
rect -64133 -37198 -63517 -36902
rect -63517 -37198 -63513 -36902
rect -64137 -37202 -63513 -37198
rect -63477 -36902 -63173 -36898
rect -63477 -37198 -63473 -36902
rect -63473 -37198 -63177 -36902
rect -63177 -37198 -63173 -36902
rect -63477 -37202 -63173 -37198
rect -63137 -36902 -62513 -36898
rect -63137 -37198 -63133 -36902
rect -63133 -37198 -62517 -36902
rect -62517 -37198 -62513 -36902
rect -63137 -37202 -62513 -37198
rect -62477 -36902 -62173 -36898
rect -62477 -37198 -62473 -36902
rect -62473 -37198 -62177 -36902
rect -62177 -37198 -62173 -36902
rect -62477 -37202 -62173 -37198
rect -62137 -36902 -61513 -36898
rect -62137 -37198 -62133 -36902
rect -62133 -37198 -61517 -36902
rect -61517 -37198 -61513 -36902
rect -62137 -37202 -61513 -37198
rect -61477 -36902 -61173 -36898
rect -61477 -37198 -61473 -36902
rect -61473 -37198 -61177 -36902
rect -61177 -37198 -61173 -36902
rect -61477 -37202 -61173 -37198
rect -61137 -36902 -60513 -36898
rect -61137 -37198 -61133 -36902
rect -61133 -37198 -60517 -36902
rect -60517 -37198 -60513 -36902
rect -61137 -37202 -60513 -37198
rect -60477 -36902 -60173 -36898
rect -60477 -37198 -60473 -36902
rect -60473 -37198 -60177 -36902
rect -60177 -37198 -60173 -36902
rect -60477 -37202 -60173 -37198
rect -60137 -36902 -59513 -36898
rect -60137 -37198 -60133 -36902
rect -60133 -37198 -59517 -36902
rect -59517 -37198 -59513 -36902
rect -60137 -37202 -59513 -37198
rect -59477 -36902 -59173 -36898
rect -59477 -37198 -59473 -36902
rect -59473 -37198 -59177 -36902
rect -59177 -37198 -59173 -36902
rect -59477 -37202 -59173 -37198
rect -59137 -36902 -58513 -36898
rect -59137 -37198 -59133 -36902
rect -59133 -37198 -58517 -36902
rect -58517 -37198 -58513 -36902
rect -59137 -37202 -58513 -37198
rect -58477 -36902 -58173 -36898
rect -58477 -37198 -58473 -36902
rect -58473 -37198 -58177 -36902
rect -58177 -37198 -58173 -36902
rect -58477 -37202 -58173 -37198
rect -58137 -36902 -57513 -36898
rect -58137 -37198 -58133 -36902
rect -58133 -37198 -57517 -36902
rect -57517 -37198 -57513 -36902
rect -58137 -37202 -57513 -37198
rect -57477 -36902 -57173 -36898
rect -57477 -37198 -57473 -36902
rect -57473 -37198 -57177 -36902
rect -57177 -37198 -57173 -36902
rect -57477 -37202 -57173 -37198
rect -57137 -36902 -56513 -36898
rect -57137 -37198 -57133 -36902
rect -57133 -37198 -56517 -36902
rect -56517 -37198 -56513 -36902
rect -57137 -37202 -56513 -37198
rect -56477 -36902 -56173 -36898
rect -56477 -37198 -56473 -36902
rect -56473 -37198 -56177 -36902
rect -56177 -37198 -56173 -36902
rect -56477 -37202 -56173 -37198
rect -56137 -36902 -55513 -36898
rect -56137 -37198 -56133 -36902
rect -56133 -37198 -55517 -36902
rect -55517 -37198 -55513 -36902
rect -56137 -37202 -55513 -37198
rect -55477 -36902 -55173 -36898
rect -55477 -37198 -55473 -36902
rect -55473 -37198 -55177 -36902
rect -55177 -37198 -55173 -36902
rect -55477 -37202 -55173 -37198
rect -55137 -36902 -54513 -36898
rect -55137 -37198 -55133 -36902
rect -55133 -37198 -54517 -36902
rect -54517 -37198 -54513 -36902
rect -55137 -37202 -54513 -37198
rect -54477 -36902 -54173 -36898
rect -54477 -37198 -54473 -36902
rect -54473 -37198 -54177 -36902
rect -54177 -37198 -54173 -36902
rect -54477 -37202 -54173 -37198
rect -54137 -36902 -53513 -36898
rect -54137 -37198 -54133 -36902
rect -54133 -37198 -53517 -36902
rect -53517 -37198 -53513 -36902
rect -54137 -37202 -53513 -37198
rect -53477 -36902 -53173 -36898
rect -53477 -37198 -53473 -36902
rect -53473 -37198 -53177 -36902
rect -53177 -37198 -53173 -36902
rect -53477 -37202 -53173 -37198
rect -53137 -36902 -52513 -36898
rect -53137 -37198 -53133 -36902
rect -53133 -37198 -52517 -36902
rect -52517 -37198 -52513 -36902
rect -53137 -37202 -52513 -37198
rect -52477 -36902 -52173 -36898
rect -52477 -37198 -52473 -36902
rect -52473 -37198 -52177 -36902
rect -52177 -37198 -52173 -36902
rect -52477 -37202 -52173 -37198
rect -52137 -36902 -51513 -36898
rect -52137 -37198 -52133 -36902
rect -52133 -37198 -51517 -36902
rect -51517 -37198 -51513 -36902
rect -52137 -37202 -51513 -37198
rect -51477 -36902 -51173 -36898
rect -51477 -37198 -51473 -36902
rect -51473 -37198 -51177 -36902
rect -51177 -37198 -51173 -36902
rect -51477 -37202 -51173 -37198
rect -51137 -36902 -50513 -36898
rect -51137 -37198 -51133 -36902
rect -51133 -37198 -50517 -36902
rect -50517 -37198 -50513 -36902
rect -51137 -37202 -50513 -37198
rect -50477 -36902 -50173 -36898
rect -50477 -37198 -50473 -36902
rect -50473 -37198 -50177 -36902
rect -50177 -37198 -50173 -36902
rect -50477 -37202 -50173 -37198
rect -50137 -36902 -49513 -36898
rect -50137 -37198 -50133 -36902
rect -50133 -37198 -49517 -36902
rect -49517 -37198 -49513 -36902
rect -50137 -37202 -49513 -37198
rect -49477 -36902 -49173 -36898
rect -49477 -37198 -49473 -36902
rect -49473 -37198 -49177 -36902
rect -49177 -37198 -49173 -36902
rect -49477 -37202 -49173 -37198
rect -49137 -36902 -48833 -36898
rect -49137 -37198 -49133 -36902
rect -49133 -37198 -48837 -36902
rect -48837 -37198 -48833 -36902
rect -49137 -37202 -48833 -37198
rect -74477 -37242 -74173 -37238
rect -74477 -37858 -74473 -37242
rect -74473 -37858 -74177 -37242
rect -74177 -37858 -74173 -37242
rect -74477 -37862 -74173 -37858
rect -73477 -37242 -73173 -37238
rect -73477 -37858 -73473 -37242
rect -73473 -37858 -73177 -37242
rect -73177 -37858 -73173 -37242
rect -73477 -37862 -73173 -37858
rect -72477 -37242 -72173 -37238
rect -72477 -37858 -72473 -37242
rect -72473 -37858 -72177 -37242
rect -72177 -37858 -72173 -37242
rect -72477 -37862 -72173 -37858
rect -71477 -37242 -71173 -37238
rect -71477 -37858 -71473 -37242
rect -71473 -37858 -71177 -37242
rect -71177 -37858 -71173 -37242
rect -71477 -37862 -71173 -37858
rect -70477 -37242 -70173 -37238
rect -70477 -37858 -70473 -37242
rect -70473 -37858 -70177 -37242
rect -70177 -37858 -70173 -37242
rect -70477 -37862 -70173 -37858
rect -69477 -37242 -69173 -37238
rect -69477 -37858 -69473 -37242
rect -69473 -37858 -69177 -37242
rect -69177 -37858 -69173 -37242
rect -69477 -37862 -69173 -37858
rect -68477 -37242 -68173 -37238
rect -68477 -37858 -68473 -37242
rect -68473 -37858 -68177 -37242
rect -68177 -37858 -68173 -37242
rect -68477 -37862 -68173 -37858
rect -67477 -37242 -67173 -37238
rect -67477 -37858 -67473 -37242
rect -67473 -37858 -67177 -37242
rect -67177 -37858 -67173 -37242
rect -67477 -37862 -67173 -37858
rect -66477 -37242 -66173 -37238
rect -66477 -37858 -66473 -37242
rect -66473 -37858 -66177 -37242
rect -66177 -37858 -66173 -37242
rect -66477 -37862 -66173 -37858
rect -65477 -37242 -65173 -37238
rect -65477 -37858 -65473 -37242
rect -65473 -37858 -65177 -37242
rect -65177 -37858 -65173 -37242
rect -65477 -37862 -65173 -37858
rect -64477 -37242 -64173 -37238
rect -64477 -37858 -64473 -37242
rect -64473 -37858 -64177 -37242
rect -64177 -37858 -64173 -37242
rect -64477 -37862 -64173 -37858
rect -63477 -37242 -63173 -37238
rect -63477 -37858 -63473 -37242
rect -63473 -37858 -63177 -37242
rect -63177 -37858 -63173 -37242
rect -63477 -37862 -63173 -37858
rect -62477 -37242 -62173 -37238
rect -62477 -37858 -62473 -37242
rect -62473 -37858 -62177 -37242
rect -62177 -37858 -62173 -37242
rect -62477 -37862 -62173 -37858
rect -61477 -37242 -61173 -37238
rect -61477 -37858 -61473 -37242
rect -61473 -37858 -61177 -37242
rect -61177 -37858 -61173 -37242
rect -61477 -37862 -61173 -37858
rect -60477 -37242 -60173 -37238
rect -60477 -37858 -60473 -37242
rect -60473 -37858 -60177 -37242
rect -60177 -37858 -60173 -37242
rect -60477 -37862 -60173 -37858
rect -59477 -37242 -59173 -37238
rect -59477 -37858 -59473 -37242
rect -59473 -37858 -59177 -37242
rect -59177 -37858 -59173 -37242
rect -59477 -37862 -59173 -37858
rect -58477 -37242 -58173 -37238
rect -58477 -37858 -58473 -37242
rect -58473 -37858 -58177 -37242
rect -58177 -37858 -58173 -37242
rect -58477 -37862 -58173 -37858
rect -57477 -37242 -57173 -37238
rect -57477 -37858 -57473 -37242
rect -57473 -37858 -57177 -37242
rect -57177 -37858 -57173 -37242
rect -57477 -37862 -57173 -37858
rect -56477 -37242 -56173 -37238
rect -56477 -37858 -56473 -37242
rect -56473 -37858 -56177 -37242
rect -56177 -37858 -56173 -37242
rect -56477 -37862 -56173 -37858
rect -55477 -37242 -55173 -37238
rect -55477 -37858 -55473 -37242
rect -55473 -37858 -55177 -37242
rect -55177 -37858 -55173 -37242
rect -55477 -37862 -55173 -37858
rect -54477 -37242 -54173 -37238
rect -54477 -37858 -54473 -37242
rect -54473 -37858 -54177 -37242
rect -54177 -37858 -54173 -37242
rect -54477 -37862 -54173 -37858
rect -53477 -37242 -53173 -37238
rect -53477 -37858 -53473 -37242
rect -53473 -37858 -53177 -37242
rect -53177 -37858 -53173 -37242
rect -53477 -37862 -53173 -37858
rect -52477 -37242 -52173 -37238
rect -52477 -37858 -52473 -37242
rect -52473 -37858 -52177 -37242
rect -52177 -37858 -52173 -37242
rect -52477 -37862 -52173 -37858
rect -51477 -37242 -51173 -37238
rect -51477 -37858 -51473 -37242
rect -51473 -37858 -51177 -37242
rect -51177 -37858 -51173 -37242
rect -51477 -37862 -51173 -37858
rect -50477 -37242 -50173 -37238
rect -50477 -37858 -50473 -37242
rect -50473 -37858 -50177 -37242
rect -50177 -37858 -50173 -37242
rect -50477 -37862 -50173 -37858
rect -49477 -37242 -49173 -37238
rect -49477 -37858 -49473 -37242
rect -49473 -37858 -49177 -37242
rect -49177 -37858 -49173 -37242
rect -49477 -37862 -49173 -37858
rect -74817 -37902 -74513 -37898
rect -74817 -38198 -74813 -37902
rect -74813 -38198 -74517 -37902
rect -74517 -38198 -74513 -37902
rect -74817 -38202 -74513 -38198
rect -74477 -37902 -74173 -37898
rect -74477 -38198 -74473 -37902
rect -74473 -38198 -74177 -37902
rect -74177 -38198 -74173 -37902
rect -74477 -38202 -74173 -38198
rect -74137 -37902 -73513 -37898
rect -74137 -38198 -74133 -37902
rect -74133 -38198 -73517 -37902
rect -73517 -38198 -73513 -37902
rect -74137 -38202 -73513 -38198
rect -73477 -37902 -73173 -37898
rect -73477 -38198 -73473 -37902
rect -73473 -38198 -73177 -37902
rect -73177 -38198 -73173 -37902
rect -73477 -38202 -73173 -38198
rect -73137 -37902 -72513 -37898
rect -73137 -38198 -73133 -37902
rect -73133 -38198 -72517 -37902
rect -72517 -38198 -72513 -37902
rect -73137 -38202 -72513 -38198
rect -72477 -37902 -72173 -37898
rect -72477 -38198 -72473 -37902
rect -72473 -38198 -72177 -37902
rect -72177 -38198 -72173 -37902
rect -72477 -38202 -72173 -38198
rect -72137 -37902 -71513 -37898
rect -72137 -38198 -72133 -37902
rect -72133 -38198 -71517 -37902
rect -71517 -38198 -71513 -37902
rect -72137 -38202 -71513 -38198
rect -71477 -37902 -71173 -37898
rect -71477 -38198 -71473 -37902
rect -71473 -38198 -71177 -37902
rect -71177 -38198 -71173 -37902
rect -71477 -38202 -71173 -38198
rect -71137 -37902 -70513 -37898
rect -71137 -38198 -71133 -37902
rect -71133 -38198 -70517 -37902
rect -70517 -38198 -70513 -37902
rect -71137 -38202 -70513 -38198
rect -70477 -37902 -70173 -37898
rect -70477 -38198 -70473 -37902
rect -70473 -38198 -70177 -37902
rect -70177 -38198 -70173 -37902
rect -70477 -38202 -70173 -38198
rect -70137 -37902 -69513 -37898
rect -70137 -38198 -70133 -37902
rect -70133 -38198 -69517 -37902
rect -69517 -38198 -69513 -37902
rect -70137 -38202 -69513 -38198
rect -69477 -37902 -69173 -37898
rect -69477 -38198 -69473 -37902
rect -69473 -38198 -69177 -37902
rect -69177 -38198 -69173 -37902
rect -69477 -38202 -69173 -38198
rect -69137 -37902 -68513 -37898
rect -69137 -38198 -69133 -37902
rect -69133 -38198 -68517 -37902
rect -68517 -38198 -68513 -37902
rect -69137 -38202 -68513 -38198
rect -68477 -37902 -68173 -37898
rect -68477 -38198 -68473 -37902
rect -68473 -38198 -68177 -37902
rect -68177 -38198 -68173 -37902
rect -68477 -38202 -68173 -38198
rect -68137 -37902 -67513 -37898
rect -68137 -38198 -68133 -37902
rect -68133 -38198 -67517 -37902
rect -67517 -38198 -67513 -37902
rect -68137 -38202 -67513 -38198
rect -67477 -37902 -67173 -37898
rect -67477 -38198 -67473 -37902
rect -67473 -38198 -67177 -37902
rect -67177 -38198 -67173 -37902
rect -67477 -38202 -67173 -38198
rect -67137 -37902 -66513 -37898
rect -67137 -38198 -67133 -37902
rect -67133 -38198 -66517 -37902
rect -66517 -38198 -66513 -37902
rect -67137 -38202 -66513 -38198
rect -66477 -37902 -66173 -37898
rect -66477 -38198 -66473 -37902
rect -66473 -38198 -66177 -37902
rect -66177 -38198 -66173 -37902
rect -66477 -38202 -66173 -38198
rect -66137 -37902 -65513 -37898
rect -66137 -38198 -66133 -37902
rect -66133 -38198 -65517 -37902
rect -65517 -38198 -65513 -37902
rect -66137 -38202 -65513 -38198
rect -65477 -37902 -65173 -37898
rect -65477 -38198 -65473 -37902
rect -65473 -38198 -65177 -37902
rect -65177 -38198 -65173 -37902
rect -65477 -38202 -65173 -38198
rect -65137 -37902 -64513 -37898
rect -65137 -38198 -65133 -37902
rect -65133 -38198 -64517 -37902
rect -64517 -38198 -64513 -37902
rect -65137 -38202 -64513 -38198
rect -64477 -37902 -64173 -37898
rect -64477 -38198 -64473 -37902
rect -64473 -38198 -64177 -37902
rect -64177 -38198 -64173 -37902
rect -64477 -38202 -64173 -38198
rect -64137 -37902 -63513 -37898
rect -64137 -38198 -64133 -37902
rect -64133 -38198 -63517 -37902
rect -63517 -38198 -63513 -37902
rect -64137 -38202 -63513 -38198
rect -63477 -37902 -63173 -37898
rect -63477 -38198 -63473 -37902
rect -63473 -38198 -63177 -37902
rect -63177 -38198 -63173 -37902
rect -63477 -38202 -63173 -38198
rect -63137 -37902 -62513 -37898
rect -63137 -38198 -63133 -37902
rect -63133 -38198 -62517 -37902
rect -62517 -38198 -62513 -37902
rect -63137 -38202 -62513 -38198
rect -62477 -37902 -62173 -37898
rect -62477 -38198 -62473 -37902
rect -62473 -38198 -62177 -37902
rect -62177 -38198 -62173 -37902
rect -62477 -38202 -62173 -38198
rect -62137 -37902 -61513 -37898
rect -62137 -38198 -62133 -37902
rect -62133 -38198 -61517 -37902
rect -61517 -38198 -61513 -37902
rect -62137 -38202 -61513 -38198
rect -61477 -37902 -61173 -37898
rect -61477 -38198 -61473 -37902
rect -61473 -38198 -61177 -37902
rect -61177 -38198 -61173 -37902
rect -61477 -38202 -61173 -38198
rect -61137 -37902 -60513 -37898
rect -61137 -38198 -61133 -37902
rect -61133 -38198 -60517 -37902
rect -60517 -38198 -60513 -37902
rect -61137 -38202 -60513 -38198
rect -60477 -37902 -60173 -37898
rect -60477 -38198 -60473 -37902
rect -60473 -38198 -60177 -37902
rect -60177 -38198 -60173 -37902
rect -60477 -38202 -60173 -38198
rect -60137 -37902 -59513 -37898
rect -60137 -38198 -60133 -37902
rect -60133 -38198 -59517 -37902
rect -59517 -38198 -59513 -37902
rect -60137 -38202 -59513 -38198
rect -59477 -37902 -59173 -37898
rect -59477 -38198 -59473 -37902
rect -59473 -38198 -59177 -37902
rect -59177 -38198 -59173 -37902
rect -59477 -38202 -59173 -38198
rect -59137 -37902 -58513 -37898
rect -59137 -38198 -59133 -37902
rect -59133 -38198 -58517 -37902
rect -58517 -38198 -58513 -37902
rect -59137 -38202 -58513 -38198
rect -58477 -37902 -58173 -37898
rect -58477 -38198 -58473 -37902
rect -58473 -38198 -58177 -37902
rect -58177 -38198 -58173 -37902
rect -58477 -38202 -58173 -38198
rect -58137 -37902 -57513 -37898
rect -58137 -38198 -58133 -37902
rect -58133 -38198 -57517 -37902
rect -57517 -38198 -57513 -37902
rect -58137 -38202 -57513 -38198
rect -57477 -37902 -57173 -37898
rect -57477 -38198 -57473 -37902
rect -57473 -38198 -57177 -37902
rect -57177 -38198 -57173 -37902
rect -57477 -38202 -57173 -38198
rect -57137 -37902 -56513 -37898
rect -57137 -38198 -57133 -37902
rect -57133 -38198 -56517 -37902
rect -56517 -38198 -56513 -37902
rect -57137 -38202 -56513 -38198
rect -56477 -37902 -56173 -37898
rect -56477 -38198 -56473 -37902
rect -56473 -38198 -56177 -37902
rect -56177 -38198 -56173 -37902
rect -56477 -38202 -56173 -38198
rect -56137 -37902 -55513 -37898
rect -56137 -38198 -56133 -37902
rect -56133 -38198 -55517 -37902
rect -55517 -38198 -55513 -37902
rect -56137 -38202 -55513 -38198
rect -55477 -37902 -55173 -37898
rect -55477 -38198 -55473 -37902
rect -55473 -38198 -55177 -37902
rect -55177 -38198 -55173 -37902
rect -55477 -38202 -55173 -38198
rect -55137 -37902 -54513 -37898
rect -55137 -38198 -55133 -37902
rect -55133 -38198 -54517 -37902
rect -54517 -38198 -54513 -37902
rect -55137 -38202 -54513 -38198
rect -54477 -37902 -54173 -37898
rect -54477 -38198 -54473 -37902
rect -54473 -38198 -54177 -37902
rect -54177 -38198 -54173 -37902
rect -54477 -38202 -54173 -38198
rect -54137 -37902 -53513 -37898
rect -54137 -38198 -54133 -37902
rect -54133 -38198 -53517 -37902
rect -53517 -38198 -53513 -37902
rect -54137 -38202 -53513 -38198
rect -53477 -37902 -53173 -37898
rect -53477 -38198 -53473 -37902
rect -53473 -38198 -53177 -37902
rect -53177 -38198 -53173 -37902
rect -53477 -38202 -53173 -38198
rect -53137 -37902 -52513 -37898
rect -53137 -38198 -53133 -37902
rect -53133 -38198 -52517 -37902
rect -52517 -38198 -52513 -37902
rect -53137 -38202 -52513 -38198
rect -52477 -37902 -52173 -37898
rect -52477 -38198 -52473 -37902
rect -52473 -38198 -52177 -37902
rect -52177 -38198 -52173 -37902
rect -52477 -38202 -52173 -38198
rect -52137 -37902 -51513 -37898
rect -52137 -38198 -52133 -37902
rect -52133 -38198 -51517 -37902
rect -51517 -38198 -51513 -37902
rect -52137 -38202 -51513 -38198
rect -51477 -37902 -51173 -37898
rect -51477 -38198 -51473 -37902
rect -51473 -38198 -51177 -37902
rect -51177 -38198 -51173 -37902
rect -51477 -38202 -51173 -38198
rect -51137 -37902 -50513 -37898
rect -51137 -38198 -51133 -37902
rect -51133 -38198 -50517 -37902
rect -50517 -38198 -50513 -37902
rect -51137 -38202 -50513 -38198
rect -50477 -37902 -50173 -37898
rect -50477 -38198 -50473 -37902
rect -50473 -38198 -50177 -37902
rect -50177 -38198 -50173 -37902
rect -50477 -38202 -50173 -38198
rect -50137 -37902 -49513 -37898
rect -50137 -38198 -50133 -37902
rect -50133 -38198 -49517 -37902
rect -49517 -38198 -49513 -37902
rect -50137 -38202 -49513 -38198
rect -49477 -37902 -49173 -37898
rect -49477 -38198 -49473 -37902
rect -49473 -38198 -49177 -37902
rect -49177 -38198 -49173 -37902
rect -49477 -38202 -49173 -38198
rect -49137 -37902 -48833 -37898
rect -49137 -38198 -49133 -37902
rect -49133 -38198 -48837 -37902
rect -48837 -38198 -48833 -37902
rect -49137 -38202 -48833 -38198
rect -74477 -38242 -74173 -38238
rect -74477 -38858 -74473 -38242
rect -74473 -38858 -74177 -38242
rect -74177 -38858 -74173 -38242
rect -74477 -38862 -74173 -38858
rect -73477 -38242 -73173 -38238
rect -73477 -38858 -73473 -38242
rect -73473 -38858 -73177 -38242
rect -73177 -38858 -73173 -38242
rect -73477 -38862 -73173 -38858
rect -72477 -38242 -72173 -38238
rect -72477 -38858 -72473 -38242
rect -72473 -38858 -72177 -38242
rect -72177 -38858 -72173 -38242
rect -72477 -38862 -72173 -38858
rect -71477 -38242 -71173 -38238
rect -71477 -38858 -71473 -38242
rect -71473 -38858 -71177 -38242
rect -71177 -38858 -71173 -38242
rect -71477 -38862 -71173 -38858
rect -70477 -38242 -70173 -38238
rect -70477 -38858 -70473 -38242
rect -70473 -38858 -70177 -38242
rect -70177 -38858 -70173 -38242
rect -70477 -38862 -70173 -38858
rect -69477 -38242 -69173 -38238
rect -69477 -38858 -69473 -38242
rect -69473 -38858 -69177 -38242
rect -69177 -38858 -69173 -38242
rect -69477 -38862 -69173 -38858
rect -68477 -38242 -68173 -38238
rect -68477 -38858 -68473 -38242
rect -68473 -38858 -68177 -38242
rect -68177 -38858 -68173 -38242
rect -68477 -38862 -68173 -38858
rect -67477 -38242 -67173 -38238
rect -67477 -38858 -67473 -38242
rect -67473 -38858 -67177 -38242
rect -67177 -38858 -67173 -38242
rect -67477 -38862 -67173 -38858
rect -66477 -38242 -66173 -38238
rect -66477 -38858 -66473 -38242
rect -66473 -38858 -66177 -38242
rect -66177 -38858 -66173 -38242
rect -66477 -38862 -66173 -38858
rect -65477 -38242 -65173 -38238
rect -65477 -38858 -65473 -38242
rect -65473 -38858 -65177 -38242
rect -65177 -38858 -65173 -38242
rect -65477 -38862 -65173 -38858
rect -64477 -38242 -64173 -38238
rect -64477 -38858 -64473 -38242
rect -64473 -38858 -64177 -38242
rect -64177 -38858 -64173 -38242
rect -64477 -38862 -64173 -38858
rect -63477 -38242 -63173 -38238
rect -63477 -38858 -63473 -38242
rect -63473 -38858 -63177 -38242
rect -63177 -38858 -63173 -38242
rect -63477 -38862 -63173 -38858
rect -62477 -38242 -62173 -38238
rect -62477 -38858 -62473 -38242
rect -62473 -38858 -62177 -38242
rect -62177 -38858 -62173 -38242
rect -62477 -38862 -62173 -38858
rect -61477 -38242 -61173 -38238
rect -61477 -38858 -61473 -38242
rect -61473 -38858 -61177 -38242
rect -61177 -38858 -61173 -38242
rect -61477 -38862 -61173 -38858
rect -60477 -38242 -60173 -38238
rect -60477 -38858 -60473 -38242
rect -60473 -38858 -60177 -38242
rect -60177 -38858 -60173 -38242
rect -60477 -38862 -60173 -38858
rect -59477 -38242 -59173 -38238
rect -59477 -38858 -59473 -38242
rect -59473 -38858 -59177 -38242
rect -59177 -38858 -59173 -38242
rect -59477 -38862 -59173 -38858
rect -58477 -38242 -58173 -38238
rect -58477 -38858 -58473 -38242
rect -58473 -38858 -58177 -38242
rect -58177 -38858 -58173 -38242
rect -58477 -38862 -58173 -38858
rect -57477 -38242 -57173 -38238
rect -57477 -38858 -57473 -38242
rect -57473 -38858 -57177 -38242
rect -57177 -38858 -57173 -38242
rect -57477 -38862 -57173 -38858
rect -56477 -38242 -56173 -38238
rect -56477 -38858 -56473 -38242
rect -56473 -38858 -56177 -38242
rect -56177 -38858 -56173 -38242
rect -56477 -38862 -56173 -38858
rect -55477 -38242 -55173 -38238
rect -55477 -38858 -55473 -38242
rect -55473 -38858 -55177 -38242
rect -55177 -38858 -55173 -38242
rect -55477 -38862 -55173 -38858
rect -54477 -38242 -54173 -38238
rect -54477 -38858 -54473 -38242
rect -54473 -38858 -54177 -38242
rect -54177 -38858 -54173 -38242
rect -54477 -38862 -54173 -38858
rect -53477 -38242 -53173 -38238
rect -53477 -38858 -53473 -38242
rect -53473 -38858 -53177 -38242
rect -53177 -38858 -53173 -38242
rect -53477 -38862 -53173 -38858
rect -52477 -38242 -52173 -38238
rect -52477 -38858 -52473 -38242
rect -52473 -38858 -52177 -38242
rect -52177 -38858 -52173 -38242
rect -52477 -38862 -52173 -38858
rect -51477 -38242 -51173 -38238
rect -51477 -38858 -51473 -38242
rect -51473 -38858 -51177 -38242
rect -51177 -38858 -51173 -38242
rect -51477 -38862 -51173 -38858
rect -50477 -38242 -50173 -38238
rect -50477 -38858 -50473 -38242
rect -50473 -38858 -50177 -38242
rect -50177 -38858 -50173 -38242
rect -50477 -38862 -50173 -38858
rect -49477 -38242 -49173 -38238
rect -49477 -38858 -49473 -38242
rect -49473 -38858 -49177 -38242
rect -49177 -38858 -49173 -38242
rect -49477 -38862 -49173 -38858
rect -74817 -38902 -74513 -38898
rect -74817 -39198 -74813 -38902
rect -74813 -39198 -74517 -38902
rect -74517 -39198 -74513 -38902
rect -74817 -39202 -74513 -39198
rect -74477 -38902 -74173 -38898
rect -74477 -39198 -74473 -38902
rect -74473 -39198 -74177 -38902
rect -74177 -39198 -74173 -38902
rect -74477 -39202 -74173 -39198
rect -74137 -38902 -73513 -38898
rect -74137 -39198 -74133 -38902
rect -74133 -39198 -73517 -38902
rect -73517 -39198 -73513 -38902
rect -74137 -39202 -73513 -39198
rect -73477 -38902 -73173 -38898
rect -73477 -39198 -73473 -38902
rect -73473 -39198 -73177 -38902
rect -73177 -39198 -73173 -38902
rect -73477 -39202 -73173 -39198
rect -73137 -38902 -72513 -38898
rect -73137 -39198 -73133 -38902
rect -73133 -39198 -72517 -38902
rect -72517 -39198 -72513 -38902
rect -73137 -39202 -72513 -39198
rect -72477 -38902 -72173 -38898
rect -72477 -39198 -72473 -38902
rect -72473 -39198 -72177 -38902
rect -72177 -39198 -72173 -38902
rect -72477 -39202 -72173 -39198
rect -72137 -38902 -71513 -38898
rect -72137 -39198 -72133 -38902
rect -72133 -39198 -71517 -38902
rect -71517 -39198 -71513 -38902
rect -72137 -39202 -71513 -39198
rect -71477 -38902 -71173 -38898
rect -71477 -39198 -71473 -38902
rect -71473 -39198 -71177 -38902
rect -71177 -39198 -71173 -38902
rect -71477 -39202 -71173 -39198
rect -71137 -38902 -70513 -38898
rect -71137 -39198 -71133 -38902
rect -71133 -39198 -70517 -38902
rect -70517 -39198 -70513 -38902
rect -71137 -39202 -70513 -39198
rect -70477 -38902 -70173 -38898
rect -70477 -39198 -70473 -38902
rect -70473 -39198 -70177 -38902
rect -70177 -39198 -70173 -38902
rect -70477 -39202 -70173 -39198
rect -70137 -38902 -69513 -38898
rect -70137 -39198 -70133 -38902
rect -70133 -39198 -69517 -38902
rect -69517 -39198 -69513 -38902
rect -70137 -39202 -69513 -39198
rect -69477 -38902 -69173 -38898
rect -69477 -39198 -69473 -38902
rect -69473 -39198 -69177 -38902
rect -69177 -39198 -69173 -38902
rect -69477 -39202 -69173 -39198
rect -69137 -38902 -68513 -38898
rect -69137 -39198 -69133 -38902
rect -69133 -39198 -68517 -38902
rect -68517 -39198 -68513 -38902
rect -69137 -39202 -68513 -39198
rect -68477 -38902 -68173 -38898
rect -68477 -39198 -68473 -38902
rect -68473 -39198 -68177 -38902
rect -68177 -39198 -68173 -38902
rect -68477 -39202 -68173 -39198
rect -68137 -38902 -67513 -38898
rect -68137 -39198 -68133 -38902
rect -68133 -39198 -67517 -38902
rect -67517 -39198 -67513 -38902
rect -68137 -39202 -67513 -39198
rect -67477 -38902 -67173 -38898
rect -67477 -39198 -67473 -38902
rect -67473 -39198 -67177 -38902
rect -67177 -39198 -67173 -38902
rect -67477 -39202 -67173 -39198
rect -67137 -38902 -66513 -38898
rect -67137 -39198 -67133 -38902
rect -67133 -39198 -66517 -38902
rect -66517 -39198 -66513 -38902
rect -67137 -39202 -66513 -39198
rect -66477 -38902 -66173 -38898
rect -66477 -39198 -66473 -38902
rect -66473 -39198 -66177 -38902
rect -66177 -39198 -66173 -38902
rect -66477 -39202 -66173 -39198
rect -66137 -38902 -65513 -38898
rect -66137 -39198 -66133 -38902
rect -66133 -39198 -65517 -38902
rect -65517 -39198 -65513 -38902
rect -66137 -39202 -65513 -39198
rect -65477 -38902 -65173 -38898
rect -65477 -39198 -65473 -38902
rect -65473 -39198 -65177 -38902
rect -65177 -39198 -65173 -38902
rect -65477 -39202 -65173 -39198
rect -65137 -38902 -64513 -38898
rect -65137 -39198 -65133 -38902
rect -65133 -39198 -64517 -38902
rect -64517 -39198 -64513 -38902
rect -65137 -39202 -64513 -39198
rect -64477 -38902 -64173 -38898
rect -64477 -39198 -64473 -38902
rect -64473 -39198 -64177 -38902
rect -64177 -39198 -64173 -38902
rect -64477 -39202 -64173 -39198
rect -64137 -38902 -63513 -38898
rect -64137 -39198 -64133 -38902
rect -64133 -39198 -63517 -38902
rect -63517 -39198 -63513 -38902
rect -64137 -39202 -63513 -39198
rect -63477 -38902 -63173 -38898
rect -63477 -39198 -63473 -38902
rect -63473 -39198 -63177 -38902
rect -63177 -39198 -63173 -38902
rect -63477 -39202 -63173 -39198
rect -63137 -38902 -62513 -38898
rect -63137 -39198 -63133 -38902
rect -63133 -39198 -62517 -38902
rect -62517 -39198 -62513 -38902
rect -63137 -39202 -62513 -39198
rect -62477 -38902 -62173 -38898
rect -62477 -39198 -62473 -38902
rect -62473 -39198 -62177 -38902
rect -62177 -39198 -62173 -38902
rect -62477 -39202 -62173 -39198
rect -62137 -38902 -61513 -38898
rect -62137 -39198 -62133 -38902
rect -62133 -39198 -61517 -38902
rect -61517 -39198 -61513 -38902
rect -62137 -39202 -61513 -39198
rect -61477 -38902 -61173 -38898
rect -61477 -39198 -61473 -38902
rect -61473 -39198 -61177 -38902
rect -61177 -39198 -61173 -38902
rect -61477 -39202 -61173 -39198
rect -61137 -38902 -60513 -38898
rect -61137 -39198 -61133 -38902
rect -61133 -39198 -60517 -38902
rect -60517 -39198 -60513 -38902
rect -61137 -39202 -60513 -39198
rect -60477 -38902 -60173 -38898
rect -60477 -39198 -60473 -38902
rect -60473 -39198 -60177 -38902
rect -60177 -39198 -60173 -38902
rect -60477 -39202 -60173 -39198
rect -60137 -38902 -59513 -38898
rect -60137 -39198 -60133 -38902
rect -60133 -39198 -59517 -38902
rect -59517 -39198 -59513 -38902
rect -60137 -39202 -59513 -39198
rect -59477 -38902 -59173 -38898
rect -59477 -39198 -59473 -38902
rect -59473 -39198 -59177 -38902
rect -59177 -39198 -59173 -38902
rect -59477 -39202 -59173 -39198
rect -59137 -38902 -58513 -38898
rect -59137 -39198 -59133 -38902
rect -59133 -39198 -58517 -38902
rect -58517 -39198 -58513 -38902
rect -59137 -39202 -58513 -39198
rect -58477 -38902 -58173 -38898
rect -58477 -39198 -58473 -38902
rect -58473 -39198 -58177 -38902
rect -58177 -39198 -58173 -38902
rect -58477 -39202 -58173 -39198
rect -58137 -38902 -57513 -38898
rect -58137 -39198 -58133 -38902
rect -58133 -39198 -57517 -38902
rect -57517 -39198 -57513 -38902
rect -58137 -39202 -57513 -39198
rect -57477 -38902 -57173 -38898
rect -57477 -39198 -57473 -38902
rect -57473 -39198 -57177 -38902
rect -57177 -39198 -57173 -38902
rect -57477 -39202 -57173 -39198
rect -57137 -38902 -56513 -38898
rect -57137 -39198 -57133 -38902
rect -57133 -39198 -56517 -38902
rect -56517 -39198 -56513 -38902
rect -57137 -39202 -56513 -39198
rect -56477 -38902 -56173 -38898
rect -56477 -39198 -56473 -38902
rect -56473 -39198 -56177 -38902
rect -56177 -39198 -56173 -38902
rect -56477 -39202 -56173 -39198
rect -56137 -38902 -55513 -38898
rect -56137 -39198 -56133 -38902
rect -56133 -39198 -55517 -38902
rect -55517 -39198 -55513 -38902
rect -56137 -39202 -55513 -39198
rect -55477 -38902 -55173 -38898
rect -55477 -39198 -55473 -38902
rect -55473 -39198 -55177 -38902
rect -55177 -39198 -55173 -38902
rect -55477 -39202 -55173 -39198
rect -55137 -38902 -54513 -38898
rect -55137 -39198 -55133 -38902
rect -55133 -39198 -54517 -38902
rect -54517 -39198 -54513 -38902
rect -55137 -39202 -54513 -39198
rect -54477 -38902 -54173 -38898
rect -54477 -39198 -54473 -38902
rect -54473 -39198 -54177 -38902
rect -54177 -39198 -54173 -38902
rect -54477 -39202 -54173 -39198
rect -54137 -38902 -53513 -38898
rect -54137 -39198 -54133 -38902
rect -54133 -39198 -53517 -38902
rect -53517 -39198 -53513 -38902
rect -54137 -39202 -53513 -39198
rect -53477 -38902 -53173 -38898
rect -53477 -39198 -53473 -38902
rect -53473 -39198 -53177 -38902
rect -53177 -39198 -53173 -38902
rect -53477 -39202 -53173 -39198
rect -53137 -38902 -52513 -38898
rect -53137 -39198 -53133 -38902
rect -53133 -39198 -52517 -38902
rect -52517 -39198 -52513 -38902
rect -53137 -39202 -52513 -39198
rect -52477 -38902 -52173 -38898
rect -52477 -39198 -52473 -38902
rect -52473 -39198 -52177 -38902
rect -52177 -39198 -52173 -38902
rect -52477 -39202 -52173 -39198
rect -52137 -38902 -51513 -38898
rect -52137 -39198 -52133 -38902
rect -52133 -39198 -51517 -38902
rect -51517 -39198 -51513 -38902
rect -52137 -39202 -51513 -39198
rect -51477 -38902 -51173 -38898
rect -51477 -39198 -51473 -38902
rect -51473 -39198 -51177 -38902
rect -51177 -39198 -51173 -38902
rect -51477 -39202 -51173 -39198
rect -51137 -38902 -50513 -38898
rect -51137 -39198 -51133 -38902
rect -51133 -39198 -50517 -38902
rect -50517 -39198 -50513 -38902
rect -51137 -39202 -50513 -39198
rect -50477 -38902 -50173 -38898
rect -50477 -39198 -50473 -38902
rect -50473 -39198 -50177 -38902
rect -50177 -39198 -50173 -38902
rect -50477 -39202 -50173 -39198
rect -50137 -38902 -49513 -38898
rect -50137 -39198 -50133 -38902
rect -50133 -39198 -49517 -38902
rect -49517 -39198 -49513 -38902
rect -50137 -39202 -49513 -39198
rect -49477 -38902 -49173 -38898
rect -49477 -39198 -49473 -38902
rect -49473 -39198 -49177 -38902
rect -49177 -39198 -49173 -38902
rect -49477 -39202 -49173 -39198
rect -49137 -38902 -48833 -38898
rect -49137 -39198 -49133 -38902
rect -49133 -39198 -48837 -38902
rect -48837 -39198 -48833 -38902
rect -49137 -39202 -48833 -39198
rect -74477 -39242 -74173 -39238
rect -74477 -39858 -74473 -39242
rect -74473 -39858 -74177 -39242
rect -74177 -39858 -74173 -39242
rect -74477 -39862 -74173 -39858
rect -73477 -39242 -73173 -39238
rect -73477 -39858 -73473 -39242
rect -73473 -39858 -73177 -39242
rect -73177 -39858 -73173 -39242
rect -73477 -39862 -73173 -39858
rect -72477 -39242 -72173 -39238
rect -72477 -39858 -72473 -39242
rect -72473 -39858 -72177 -39242
rect -72177 -39858 -72173 -39242
rect -72477 -39862 -72173 -39858
rect -71477 -39242 -71173 -39238
rect -71477 -39858 -71473 -39242
rect -71473 -39858 -71177 -39242
rect -71177 -39858 -71173 -39242
rect -71477 -39862 -71173 -39858
rect -70477 -39242 -70173 -39238
rect -70477 -39858 -70473 -39242
rect -70473 -39858 -70177 -39242
rect -70177 -39858 -70173 -39242
rect -70477 -39862 -70173 -39858
rect -69477 -39242 -69173 -39238
rect -69477 -39858 -69473 -39242
rect -69473 -39858 -69177 -39242
rect -69177 -39858 -69173 -39242
rect -69477 -39862 -69173 -39858
rect -68477 -39242 -68173 -39238
rect -68477 -39858 -68473 -39242
rect -68473 -39858 -68177 -39242
rect -68177 -39858 -68173 -39242
rect -68477 -39862 -68173 -39858
rect -67477 -39242 -67173 -39238
rect -67477 -39858 -67473 -39242
rect -67473 -39858 -67177 -39242
rect -67177 -39858 -67173 -39242
rect -67477 -39862 -67173 -39858
rect -66477 -39242 -66173 -39238
rect -66477 -39858 -66473 -39242
rect -66473 -39858 -66177 -39242
rect -66177 -39858 -66173 -39242
rect -66477 -39862 -66173 -39858
rect -65477 -39242 -65173 -39238
rect -65477 -39858 -65473 -39242
rect -65473 -39858 -65177 -39242
rect -65177 -39858 -65173 -39242
rect -65477 -39862 -65173 -39858
rect -64477 -39242 -64173 -39238
rect -64477 -39858 -64473 -39242
rect -64473 -39858 -64177 -39242
rect -64177 -39858 -64173 -39242
rect -64477 -39862 -64173 -39858
rect -63477 -39242 -63173 -39238
rect -63477 -39858 -63473 -39242
rect -63473 -39858 -63177 -39242
rect -63177 -39858 -63173 -39242
rect -63477 -39862 -63173 -39858
rect -62477 -39242 -62173 -39238
rect -62477 -39858 -62473 -39242
rect -62473 -39858 -62177 -39242
rect -62177 -39858 -62173 -39242
rect -62477 -39862 -62173 -39858
rect -61477 -39242 -61173 -39238
rect -61477 -39858 -61473 -39242
rect -61473 -39858 -61177 -39242
rect -61177 -39858 -61173 -39242
rect -61477 -39862 -61173 -39858
rect -60477 -39242 -60173 -39238
rect -60477 -39858 -60473 -39242
rect -60473 -39858 -60177 -39242
rect -60177 -39858 -60173 -39242
rect -60477 -39862 -60173 -39858
rect -59477 -39242 -59173 -39238
rect -59477 -39858 -59473 -39242
rect -59473 -39858 -59177 -39242
rect -59177 -39858 -59173 -39242
rect -59477 -39862 -59173 -39858
rect -58477 -39242 -58173 -39238
rect -58477 -39858 -58473 -39242
rect -58473 -39858 -58177 -39242
rect -58177 -39858 -58173 -39242
rect -58477 -39862 -58173 -39858
rect -57477 -39242 -57173 -39238
rect -57477 -39858 -57473 -39242
rect -57473 -39858 -57177 -39242
rect -57177 -39858 -57173 -39242
rect -57477 -39862 -57173 -39858
rect -56477 -39242 -56173 -39238
rect -56477 -39858 -56473 -39242
rect -56473 -39858 -56177 -39242
rect -56177 -39858 -56173 -39242
rect -56477 -39862 -56173 -39858
rect -55477 -39242 -55173 -39238
rect -55477 -39858 -55473 -39242
rect -55473 -39858 -55177 -39242
rect -55177 -39858 -55173 -39242
rect -55477 -39862 -55173 -39858
rect -54477 -39242 -54173 -39238
rect -54477 -39858 -54473 -39242
rect -54473 -39858 -54177 -39242
rect -54177 -39858 -54173 -39242
rect -54477 -39862 -54173 -39858
rect -53477 -39242 -53173 -39238
rect -53477 -39858 -53473 -39242
rect -53473 -39858 -53177 -39242
rect -53177 -39858 -53173 -39242
rect -53477 -39862 -53173 -39858
rect -52477 -39242 -52173 -39238
rect -52477 -39858 -52473 -39242
rect -52473 -39858 -52177 -39242
rect -52177 -39858 -52173 -39242
rect -52477 -39862 -52173 -39858
rect -51477 -39242 -51173 -39238
rect -51477 -39858 -51473 -39242
rect -51473 -39858 -51177 -39242
rect -51177 -39858 -51173 -39242
rect -51477 -39862 -51173 -39858
rect -50477 -39242 -50173 -39238
rect -50477 -39858 -50473 -39242
rect -50473 -39858 -50177 -39242
rect -50177 -39858 -50173 -39242
rect -50477 -39862 -50173 -39858
rect -49477 -39242 -49173 -39238
rect -49477 -39858 -49473 -39242
rect -49473 -39858 -49177 -39242
rect -49177 -39858 -49173 -39242
rect -49477 -39862 -49173 -39858
rect -74817 -39902 -74513 -39898
rect -74817 -40198 -74813 -39902
rect -74813 -40198 -74517 -39902
rect -74517 -40198 -74513 -39902
rect -74817 -40202 -74513 -40198
rect -74477 -39902 -74173 -39898
rect -74477 -40198 -74473 -39902
rect -74473 -40198 -74177 -39902
rect -74177 -40198 -74173 -39902
rect -74477 -40202 -74173 -40198
rect -74137 -39902 -73513 -39898
rect -74137 -40198 -74133 -39902
rect -74133 -40198 -73517 -39902
rect -73517 -40198 -73513 -39902
rect -74137 -40202 -73513 -40198
rect -73477 -39902 -73173 -39898
rect -73477 -40198 -73473 -39902
rect -73473 -40198 -73177 -39902
rect -73177 -40198 -73173 -39902
rect -73477 -40202 -73173 -40198
rect -73137 -39902 -72513 -39898
rect -73137 -40198 -73133 -39902
rect -73133 -40198 -72517 -39902
rect -72517 -40198 -72513 -39902
rect -73137 -40202 -72513 -40198
rect -72477 -39902 -72173 -39898
rect -72477 -40198 -72473 -39902
rect -72473 -40198 -72177 -39902
rect -72177 -40198 -72173 -39902
rect -72477 -40202 -72173 -40198
rect -72137 -39902 -71513 -39898
rect -72137 -40198 -72133 -39902
rect -72133 -40198 -71517 -39902
rect -71517 -40198 -71513 -39902
rect -72137 -40202 -71513 -40198
rect -71477 -39902 -71173 -39898
rect -71477 -40198 -71473 -39902
rect -71473 -40198 -71177 -39902
rect -71177 -40198 -71173 -39902
rect -71477 -40202 -71173 -40198
rect -71137 -39902 -70513 -39898
rect -71137 -40198 -71133 -39902
rect -71133 -40198 -70517 -39902
rect -70517 -40198 -70513 -39902
rect -71137 -40202 -70513 -40198
rect -70477 -39902 -70173 -39898
rect -70477 -40198 -70473 -39902
rect -70473 -40198 -70177 -39902
rect -70177 -40198 -70173 -39902
rect -70477 -40202 -70173 -40198
rect -70137 -39902 -69513 -39898
rect -70137 -40198 -70133 -39902
rect -70133 -40198 -69517 -39902
rect -69517 -40198 -69513 -39902
rect -70137 -40202 -69513 -40198
rect -69477 -39902 -69173 -39898
rect -69477 -40198 -69473 -39902
rect -69473 -40198 -69177 -39902
rect -69177 -40198 -69173 -39902
rect -69477 -40202 -69173 -40198
rect -69137 -39902 -68513 -39898
rect -69137 -40198 -69133 -39902
rect -69133 -40198 -68517 -39902
rect -68517 -40198 -68513 -39902
rect -69137 -40202 -68513 -40198
rect -68477 -39902 -68173 -39898
rect -68477 -40198 -68473 -39902
rect -68473 -40198 -68177 -39902
rect -68177 -40198 -68173 -39902
rect -68477 -40202 -68173 -40198
rect -68137 -39902 -67513 -39898
rect -68137 -40198 -68133 -39902
rect -68133 -40198 -67517 -39902
rect -67517 -40198 -67513 -39902
rect -68137 -40202 -67513 -40198
rect -67477 -39902 -67173 -39898
rect -67477 -40198 -67473 -39902
rect -67473 -40198 -67177 -39902
rect -67177 -40198 -67173 -39902
rect -67477 -40202 -67173 -40198
rect -67137 -39902 -66513 -39898
rect -67137 -40198 -67133 -39902
rect -67133 -40198 -66517 -39902
rect -66517 -40198 -66513 -39902
rect -67137 -40202 -66513 -40198
rect -66477 -39902 -66173 -39898
rect -66477 -40198 -66473 -39902
rect -66473 -40198 -66177 -39902
rect -66177 -40198 -66173 -39902
rect -66477 -40202 -66173 -40198
rect -66137 -39902 -65513 -39898
rect -66137 -40198 -66133 -39902
rect -66133 -40198 -65517 -39902
rect -65517 -40198 -65513 -39902
rect -66137 -40202 -65513 -40198
rect -65477 -39902 -65173 -39898
rect -65477 -40198 -65473 -39902
rect -65473 -40198 -65177 -39902
rect -65177 -40198 -65173 -39902
rect -65477 -40202 -65173 -40198
rect -65137 -39902 -64513 -39898
rect -65137 -40198 -65133 -39902
rect -65133 -40198 -64517 -39902
rect -64517 -40198 -64513 -39902
rect -65137 -40202 -64513 -40198
rect -64477 -39902 -64173 -39898
rect -64477 -40198 -64473 -39902
rect -64473 -40198 -64177 -39902
rect -64177 -40198 -64173 -39902
rect -64477 -40202 -64173 -40198
rect -64137 -39902 -63513 -39898
rect -64137 -40198 -64133 -39902
rect -64133 -40198 -63517 -39902
rect -63517 -40198 -63513 -39902
rect -64137 -40202 -63513 -40198
rect -63477 -39902 -63173 -39898
rect -63477 -40198 -63473 -39902
rect -63473 -40198 -63177 -39902
rect -63177 -40198 -63173 -39902
rect -63477 -40202 -63173 -40198
rect -63137 -39902 -62513 -39898
rect -63137 -40198 -63133 -39902
rect -63133 -40198 -62517 -39902
rect -62517 -40198 -62513 -39902
rect -63137 -40202 -62513 -40198
rect -62477 -39902 -62173 -39898
rect -62477 -40198 -62473 -39902
rect -62473 -40198 -62177 -39902
rect -62177 -40198 -62173 -39902
rect -62477 -40202 -62173 -40198
rect -62137 -39902 -61513 -39898
rect -62137 -40198 -62133 -39902
rect -62133 -40198 -61517 -39902
rect -61517 -40198 -61513 -39902
rect -62137 -40202 -61513 -40198
rect -61477 -39902 -61173 -39898
rect -61477 -40198 -61473 -39902
rect -61473 -40198 -61177 -39902
rect -61177 -40198 -61173 -39902
rect -61477 -40202 -61173 -40198
rect -61137 -39902 -60513 -39898
rect -61137 -40198 -61133 -39902
rect -61133 -40198 -60517 -39902
rect -60517 -40198 -60513 -39902
rect -61137 -40202 -60513 -40198
rect -60477 -39902 -60173 -39898
rect -60477 -40198 -60473 -39902
rect -60473 -40198 -60177 -39902
rect -60177 -40198 -60173 -39902
rect -60477 -40202 -60173 -40198
rect -60137 -39902 -59513 -39898
rect -60137 -40198 -60133 -39902
rect -60133 -40198 -59517 -39902
rect -59517 -40198 -59513 -39902
rect -60137 -40202 -59513 -40198
rect -59477 -39902 -59173 -39898
rect -59477 -40198 -59473 -39902
rect -59473 -40198 -59177 -39902
rect -59177 -40198 -59173 -39902
rect -59477 -40202 -59173 -40198
rect -59137 -39902 -58513 -39898
rect -59137 -40198 -59133 -39902
rect -59133 -40198 -58517 -39902
rect -58517 -40198 -58513 -39902
rect -59137 -40202 -58513 -40198
rect -58477 -39902 -58173 -39898
rect -58477 -40198 -58473 -39902
rect -58473 -40198 -58177 -39902
rect -58177 -40198 -58173 -39902
rect -58477 -40202 -58173 -40198
rect -58137 -39902 -57513 -39898
rect -58137 -40198 -58133 -39902
rect -58133 -40198 -57517 -39902
rect -57517 -40198 -57513 -39902
rect -58137 -40202 -57513 -40198
rect -57477 -39902 -57173 -39898
rect -57477 -40198 -57473 -39902
rect -57473 -40198 -57177 -39902
rect -57177 -40198 -57173 -39902
rect -57477 -40202 -57173 -40198
rect -57137 -39902 -56513 -39898
rect -57137 -40198 -57133 -39902
rect -57133 -40198 -56517 -39902
rect -56517 -40198 -56513 -39902
rect -57137 -40202 -56513 -40198
rect -56477 -39902 -56173 -39898
rect -56477 -40198 -56473 -39902
rect -56473 -40198 -56177 -39902
rect -56177 -40198 -56173 -39902
rect -56477 -40202 -56173 -40198
rect -56137 -39902 -55513 -39898
rect -56137 -40198 -56133 -39902
rect -56133 -40198 -55517 -39902
rect -55517 -40198 -55513 -39902
rect -56137 -40202 -55513 -40198
rect -55477 -39902 -55173 -39898
rect -55477 -40198 -55473 -39902
rect -55473 -40198 -55177 -39902
rect -55177 -40198 -55173 -39902
rect -55477 -40202 -55173 -40198
rect -55137 -39902 -54513 -39898
rect -55137 -40198 -55133 -39902
rect -55133 -40198 -54517 -39902
rect -54517 -40198 -54513 -39902
rect -55137 -40202 -54513 -40198
rect -54477 -39902 -54173 -39898
rect -54477 -40198 -54473 -39902
rect -54473 -40198 -54177 -39902
rect -54177 -40198 -54173 -39902
rect -54477 -40202 -54173 -40198
rect -54137 -39902 -53513 -39898
rect -54137 -40198 -54133 -39902
rect -54133 -40198 -53517 -39902
rect -53517 -40198 -53513 -39902
rect -54137 -40202 -53513 -40198
rect -53477 -39902 -53173 -39898
rect -53477 -40198 -53473 -39902
rect -53473 -40198 -53177 -39902
rect -53177 -40198 -53173 -39902
rect -53477 -40202 -53173 -40198
rect -53137 -39902 -52513 -39898
rect -53137 -40198 -53133 -39902
rect -53133 -40198 -52517 -39902
rect -52517 -40198 -52513 -39902
rect -53137 -40202 -52513 -40198
rect -52477 -39902 -52173 -39898
rect -52477 -40198 -52473 -39902
rect -52473 -40198 -52177 -39902
rect -52177 -40198 -52173 -39902
rect -52477 -40202 -52173 -40198
rect -52137 -39902 -51513 -39898
rect -52137 -40198 -52133 -39902
rect -52133 -40198 -51517 -39902
rect -51517 -40198 -51513 -39902
rect -52137 -40202 -51513 -40198
rect -51477 -39902 -51173 -39898
rect -51477 -40198 -51473 -39902
rect -51473 -40198 -51177 -39902
rect -51177 -40198 -51173 -39902
rect -51477 -40202 -51173 -40198
rect -51137 -39902 -50513 -39898
rect -51137 -40198 -51133 -39902
rect -51133 -40198 -50517 -39902
rect -50517 -40198 -50513 -39902
rect -51137 -40202 -50513 -40198
rect -50477 -39902 -50173 -39898
rect -50477 -40198 -50473 -39902
rect -50473 -40198 -50177 -39902
rect -50177 -40198 -50173 -39902
rect -50477 -40202 -50173 -40198
rect -50137 -39902 -49513 -39898
rect -50137 -40198 -50133 -39902
rect -50133 -40198 -49517 -39902
rect -49517 -40198 -49513 -39902
rect -50137 -40202 -49513 -40198
rect -49477 -39902 -49173 -39898
rect -49477 -40198 -49473 -39902
rect -49473 -40198 -49177 -39902
rect -49177 -40198 -49173 -39902
rect -49477 -40202 -49173 -40198
rect -49137 -39902 -48833 -39898
rect -49137 -40198 -49133 -39902
rect -49133 -40198 -48837 -39902
rect -48837 -40198 -48833 -39902
rect -49137 -40202 -48833 -40198
rect -74477 -40242 -74173 -40238
rect -74477 -40858 -74473 -40242
rect -74473 -40858 -74177 -40242
rect -74177 -40858 -74173 -40242
rect -74477 -40862 -74173 -40858
rect -73477 -40242 -73173 -40238
rect -73477 -40858 -73473 -40242
rect -73473 -40858 -73177 -40242
rect -73177 -40858 -73173 -40242
rect -73477 -40862 -73173 -40858
rect -72477 -40242 -72173 -40238
rect -72477 -40858 -72473 -40242
rect -72473 -40858 -72177 -40242
rect -72177 -40858 -72173 -40242
rect -72477 -40862 -72173 -40858
rect -71477 -40242 -71173 -40238
rect -71477 -40858 -71473 -40242
rect -71473 -40858 -71177 -40242
rect -71177 -40858 -71173 -40242
rect -71477 -40862 -71173 -40858
rect -70477 -40242 -70173 -40238
rect -70477 -40858 -70473 -40242
rect -70473 -40858 -70177 -40242
rect -70177 -40858 -70173 -40242
rect -70477 -40862 -70173 -40858
rect -69477 -40242 -69173 -40238
rect -69477 -40858 -69473 -40242
rect -69473 -40858 -69177 -40242
rect -69177 -40858 -69173 -40242
rect -69477 -40862 -69173 -40858
rect -68477 -40242 -68173 -40238
rect -68477 -40858 -68473 -40242
rect -68473 -40858 -68177 -40242
rect -68177 -40858 -68173 -40242
rect -68477 -40862 -68173 -40858
rect -67477 -40242 -67173 -40238
rect -67477 -40858 -67473 -40242
rect -67473 -40858 -67177 -40242
rect -67177 -40858 -67173 -40242
rect -67477 -40862 -67173 -40858
rect -66477 -40242 -66173 -40238
rect -66477 -40858 -66473 -40242
rect -66473 -40858 -66177 -40242
rect -66177 -40858 -66173 -40242
rect -66477 -40862 -66173 -40858
rect -65477 -40242 -65173 -40238
rect -65477 -40858 -65473 -40242
rect -65473 -40858 -65177 -40242
rect -65177 -40858 -65173 -40242
rect -65477 -40862 -65173 -40858
rect -64477 -40242 -64173 -40238
rect -64477 -40858 -64473 -40242
rect -64473 -40858 -64177 -40242
rect -64177 -40858 -64173 -40242
rect -64477 -40862 -64173 -40858
rect -63477 -40242 -63173 -40238
rect -63477 -40858 -63473 -40242
rect -63473 -40858 -63177 -40242
rect -63177 -40858 -63173 -40242
rect -63477 -40862 -63173 -40858
rect -62477 -40242 -62173 -40238
rect -62477 -40858 -62473 -40242
rect -62473 -40858 -62177 -40242
rect -62177 -40858 -62173 -40242
rect -62477 -40862 -62173 -40858
rect -61477 -40242 -61173 -40238
rect -61477 -40858 -61473 -40242
rect -61473 -40858 -61177 -40242
rect -61177 -40858 -61173 -40242
rect -61477 -40862 -61173 -40858
rect -60477 -40242 -60173 -40238
rect -60477 -40858 -60473 -40242
rect -60473 -40858 -60177 -40242
rect -60177 -40858 -60173 -40242
rect -60477 -40862 -60173 -40858
rect -59477 -40242 -59173 -40238
rect -59477 -40858 -59473 -40242
rect -59473 -40858 -59177 -40242
rect -59177 -40858 -59173 -40242
rect -59477 -40862 -59173 -40858
rect -58477 -40242 -58173 -40238
rect -58477 -40858 -58473 -40242
rect -58473 -40858 -58177 -40242
rect -58177 -40858 -58173 -40242
rect -58477 -40862 -58173 -40858
rect -57477 -40242 -57173 -40238
rect -57477 -40858 -57473 -40242
rect -57473 -40858 -57177 -40242
rect -57177 -40858 -57173 -40242
rect -57477 -40862 -57173 -40858
rect -56477 -40242 -56173 -40238
rect -56477 -40858 -56473 -40242
rect -56473 -40858 -56177 -40242
rect -56177 -40858 -56173 -40242
rect -56477 -40862 -56173 -40858
rect -55477 -40242 -55173 -40238
rect -55477 -40858 -55473 -40242
rect -55473 -40858 -55177 -40242
rect -55177 -40858 -55173 -40242
rect -55477 -40862 -55173 -40858
rect -54477 -40242 -54173 -40238
rect -54477 -40858 -54473 -40242
rect -54473 -40858 -54177 -40242
rect -54177 -40858 -54173 -40242
rect -54477 -40862 -54173 -40858
rect -53477 -40242 -53173 -40238
rect -53477 -40858 -53473 -40242
rect -53473 -40858 -53177 -40242
rect -53177 -40858 -53173 -40242
rect -53477 -40862 -53173 -40858
rect -52477 -40242 -52173 -40238
rect -52477 -40858 -52473 -40242
rect -52473 -40858 -52177 -40242
rect -52177 -40858 -52173 -40242
rect -52477 -40862 -52173 -40858
rect -51477 -40242 -51173 -40238
rect -51477 -40858 -51473 -40242
rect -51473 -40858 -51177 -40242
rect -51177 -40858 -51173 -40242
rect -51477 -40862 -51173 -40858
rect -50477 -40242 -50173 -40238
rect -50477 -40858 -50473 -40242
rect -50473 -40858 -50177 -40242
rect -50177 -40858 -50173 -40242
rect -50477 -40862 -50173 -40858
rect -49477 -40242 -49173 -40238
rect -49477 -40858 -49473 -40242
rect -49473 -40858 -49177 -40242
rect -49177 -40858 -49173 -40242
rect -49477 -40862 -49173 -40858
rect -74817 -40902 -74513 -40898
rect -74817 -41198 -74813 -40902
rect -74813 -41198 -74517 -40902
rect -74517 -41198 -74513 -40902
rect -74817 -41202 -74513 -41198
rect -74477 -40902 -74173 -40898
rect -74477 -41198 -74473 -40902
rect -74473 -41198 -74177 -40902
rect -74177 -41198 -74173 -40902
rect -74477 -41202 -74173 -41198
rect -74137 -40902 -73513 -40898
rect -74137 -41198 -74133 -40902
rect -74133 -41198 -73517 -40902
rect -73517 -41198 -73513 -40902
rect -74137 -41202 -73513 -41198
rect -73477 -40902 -73173 -40898
rect -73477 -41198 -73473 -40902
rect -73473 -41198 -73177 -40902
rect -73177 -41198 -73173 -40902
rect -73477 -41202 -73173 -41198
rect -73137 -40902 -72513 -40898
rect -73137 -41198 -73133 -40902
rect -73133 -41198 -72517 -40902
rect -72517 -41198 -72513 -40902
rect -73137 -41202 -72513 -41198
rect -72477 -40902 -72173 -40898
rect -72477 -41198 -72473 -40902
rect -72473 -41198 -72177 -40902
rect -72177 -41198 -72173 -40902
rect -72477 -41202 -72173 -41198
rect -72137 -40902 -71513 -40898
rect -72137 -41198 -72133 -40902
rect -72133 -41198 -71517 -40902
rect -71517 -41198 -71513 -40902
rect -72137 -41202 -71513 -41198
rect -71477 -40902 -71173 -40898
rect -71477 -41198 -71473 -40902
rect -71473 -41198 -71177 -40902
rect -71177 -41198 -71173 -40902
rect -71477 -41202 -71173 -41198
rect -71137 -40902 -70513 -40898
rect -71137 -41198 -71133 -40902
rect -71133 -41198 -70517 -40902
rect -70517 -41198 -70513 -40902
rect -71137 -41202 -70513 -41198
rect -70477 -40902 -70173 -40898
rect -70477 -41198 -70473 -40902
rect -70473 -41198 -70177 -40902
rect -70177 -41198 -70173 -40902
rect -70477 -41202 -70173 -41198
rect -70137 -40902 -69513 -40898
rect -70137 -41198 -70133 -40902
rect -70133 -41198 -69517 -40902
rect -69517 -41198 -69513 -40902
rect -70137 -41202 -69513 -41198
rect -69477 -40902 -69173 -40898
rect -69477 -41198 -69473 -40902
rect -69473 -41198 -69177 -40902
rect -69177 -41198 -69173 -40902
rect -69477 -41202 -69173 -41198
rect -69137 -40902 -68513 -40898
rect -69137 -41198 -69133 -40902
rect -69133 -41198 -68517 -40902
rect -68517 -41198 -68513 -40902
rect -69137 -41202 -68513 -41198
rect -68477 -40902 -68173 -40898
rect -68477 -41198 -68473 -40902
rect -68473 -41198 -68177 -40902
rect -68177 -41198 -68173 -40902
rect -68477 -41202 -68173 -41198
rect -68137 -40902 -67513 -40898
rect -68137 -41198 -68133 -40902
rect -68133 -41198 -67517 -40902
rect -67517 -41198 -67513 -40902
rect -68137 -41202 -67513 -41198
rect -67477 -40902 -67173 -40898
rect -67477 -41198 -67473 -40902
rect -67473 -41198 -67177 -40902
rect -67177 -41198 -67173 -40902
rect -67477 -41202 -67173 -41198
rect -67137 -40902 -66513 -40898
rect -67137 -41198 -67133 -40902
rect -67133 -41198 -66517 -40902
rect -66517 -41198 -66513 -40902
rect -67137 -41202 -66513 -41198
rect -66477 -40902 -66173 -40898
rect -66477 -41198 -66473 -40902
rect -66473 -41198 -66177 -40902
rect -66177 -41198 -66173 -40902
rect -66477 -41202 -66173 -41198
rect -66137 -40902 -65513 -40898
rect -66137 -41198 -66133 -40902
rect -66133 -41198 -65517 -40902
rect -65517 -41198 -65513 -40902
rect -66137 -41202 -65513 -41198
rect -65477 -40902 -65173 -40898
rect -65477 -41198 -65473 -40902
rect -65473 -41198 -65177 -40902
rect -65177 -41198 -65173 -40902
rect -65477 -41202 -65173 -41198
rect -65137 -40902 -64513 -40898
rect -65137 -41198 -65133 -40902
rect -65133 -41198 -64517 -40902
rect -64517 -41198 -64513 -40902
rect -65137 -41202 -64513 -41198
rect -64477 -40902 -64173 -40898
rect -64477 -41198 -64473 -40902
rect -64473 -41198 -64177 -40902
rect -64177 -41198 -64173 -40902
rect -64477 -41202 -64173 -41198
rect -64137 -40902 -63513 -40898
rect -64137 -41198 -64133 -40902
rect -64133 -41198 -63517 -40902
rect -63517 -41198 -63513 -40902
rect -64137 -41202 -63513 -41198
rect -63477 -40902 -63173 -40898
rect -63477 -41198 -63473 -40902
rect -63473 -41198 -63177 -40902
rect -63177 -41198 -63173 -40902
rect -63477 -41202 -63173 -41198
rect -63137 -40902 -62513 -40898
rect -63137 -41198 -63133 -40902
rect -63133 -41198 -62517 -40902
rect -62517 -41198 -62513 -40902
rect -63137 -41202 -62513 -41198
rect -62477 -40902 -62173 -40898
rect -62477 -41198 -62473 -40902
rect -62473 -41198 -62177 -40902
rect -62177 -41198 -62173 -40902
rect -62477 -41202 -62173 -41198
rect -62137 -40902 -61513 -40898
rect -62137 -41198 -62133 -40902
rect -62133 -41198 -61517 -40902
rect -61517 -41198 -61513 -40902
rect -62137 -41202 -61513 -41198
rect -61477 -40902 -61173 -40898
rect -61477 -41198 -61473 -40902
rect -61473 -41198 -61177 -40902
rect -61177 -41198 -61173 -40902
rect -61477 -41202 -61173 -41198
rect -61137 -40902 -60513 -40898
rect -61137 -41198 -61133 -40902
rect -61133 -41198 -60517 -40902
rect -60517 -41198 -60513 -40902
rect -61137 -41202 -60513 -41198
rect -60477 -40902 -60173 -40898
rect -60477 -41198 -60473 -40902
rect -60473 -41198 -60177 -40902
rect -60177 -41198 -60173 -40902
rect -60477 -41202 -60173 -41198
rect -60137 -40902 -59513 -40898
rect -60137 -41198 -60133 -40902
rect -60133 -41198 -59517 -40902
rect -59517 -41198 -59513 -40902
rect -60137 -41202 -59513 -41198
rect -59477 -40902 -59173 -40898
rect -59477 -41198 -59473 -40902
rect -59473 -41198 -59177 -40902
rect -59177 -41198 -59173 -40902
rect -59477 -41202 -59173 -41198
rect -59137 -40902 -58513 -40898
rect -59137 -41198 -59133 -40902
rect -59133 -41198 -58517 -40902
rect -58517 -41198 -58513 -40902
rect -59137 -41202 -58513 -41198
rect -58477 -40902 -58173 -40898
rect -58477 -41198 -58473 -40902
rect -58473 -41198 -58177 -40902
rect -58177 -41198 -58173 -40902
rect -58477 -41202 -58173 -41198
rect -58137 -40902 -57513 -40898
rect -58137 -41198 -58133 -40902
rect -58133 -41198 -57517 -40902
rect -57517 -41198 -57513 -40902
rect -58137 -41202 -57513 -41198
rect -57477 -40902 -57173 -40898
rect -57477 -41198 -57473 -40902
rect -57473 -41198 -57177 -40902
rect -57177 -41198 -57173 -40902
rect -57477 -41202 -57173 -41198
rect -57137 -40902 -56513 -40898
rect -57137 -41198 -57133 -40902
rect -57133 -41198 -56517 -40902
rect -56517 -41198 -56513 -40902
rect -57137 -41202 -56513 -41198
rect -56477 -40902 -56173 -40898
rect -56477 -41198 -56473 -40902
rect -56473 -41198 -56177 -40902
rect -56177 -41198 -56173 -40902
rect -56477 -41202 -56173 -41198
rect -56137 -40902 -55513 -40898
rect -56137 -41198 -56133 -40902
rect -56133 -41198 -55517 -40902
rect -55517 -41198 -55513 -40902
rect -56137 -41202 -55513 -41198
rect -55477 -40902 -55173 -40898
rect -55477 -41198 -55473 -40902
rect -55473 -41198 -55177 -40902
rect -55177 -41198 -55173 -40902
rect -55477 -41202 -55173 -41198
rect -55137 -40902 -54513 -40898
rect -55137 -41198 -55133 -40902
rect -55133 -41198 -54517 -40902
rect -54517 -41198 -54513 -40902
rect -55137 -41202 -54513 -41198
rect -54477 -40902 -54173 -40898
rect -54477 -41198 -54473 -40902
rect -54473 -41198 -54177 -40902
rect -54177 -41198 -54173 -40902
rect -54477 -41202 -54173 -41198
rect -54137 -40902 -53513 -40898
rect -54137 -41198 -54133 -40902
rect -54133 -41198 -53517 -40902
rect -53517 -41198 -53513 -40902
rect -54137 -41202 -53513 -41198
rect -53477 -40902 -53173 -40898
rect -53477 -41198 -53473 -40902
rect -53473 -41198 -53177 -40902
rect -53177 -41198 -53173 -40902
rect -53477 -41202 -53173 -41198
rect -53137 -40902 -52513 -40898
rect -53137 -41198 -53133 -40902
rect -53133 -41198 -52517 -40902
rect -52517 -41198 -52513 -40902
rect -53137 -41202 -52513 -41198
rect -52477 -40902 -52173 -40898
rect -52477 -41198 -52473 -40902
rect -52473 -41198 -52177 -40902
rect -52177 -41198 -52173 -40902
rect -52477 -41202 -52173 -41198
rect -52137 -40902 -51513 -40898
rect -52137 -41198 -52133 -40902
rect -52133 -41198 -51517 -40902
rect -51517 -41198 -51513 -40902
rect -52137 -41202 -51513 -41198
rect -51477 -40902 -51173 -40898
rect -51477 -41198 -51473 -40902
rect -51473 -41198 -51177 -40902
rect -51177 -41198 -51173 -40902
rect -51477 -41202 -51173 -41198
rect -51137 -40902 -50513 -40898
rect -51137 -41198 -51133 -40902
rect -51133 -41198 -50517 -40902
rect -50517 -41198 -50513 -40902
rect -51137 -41202 -50513 -41198
rect -50477 -40902 -50173 -40898
rect -50477 -41198 -50473 -40902
rect -50473 -41198 -50177 -40902
rect -50177 -41198 -50173 -40902
rect -50477 -41202 -50173 -41198
rect -50137 -40902 -49513 -40898
rect -50137 -41198 -50133 -40902
rect -50133 -41198 -49517 -40902
rect -49517 -41198 -49513 -40902
rect -50137 -41202 -49513 -41198
rect -49477 -40902 -49173 -40898
rect -49477 -41198 -49473 -40902
rect -49473 -41198 -49177 -40902
rect -49177 -41198 -49173 -40902
rect -49477 -41202 -49173 -41198
rect -49137 -40902 -48833 -40898
rect -49137 -41198 -49133 -40902
rect -49133 -41198 -48837 -40902
rect -48837 -41198 -48833 -40902
rect -49137 -41202 -48833 -41198
rect -74477 -41242 -74173 -41238
rect -74477 -41858 -74473 -41242
rect -74473 -41858 -74177 -41242
rect -74177 -41858 -74173 -41242
rect -74477 -41862 -74173 -41858
rect -73477 -41242 -73173 -41238
rect -73477 -41858 -73473 -41242
rect -73473 -41858 -73177 -41242
rect -73177 -41858 -73173 -41242
rect -73477 -41862 -73173 -41858
rect -72477 -41242 -72173 -41238
rect -72477 -41858 -72473 -41242
rect -72473 -41858 -72177 -41242
rect -72177 -41858 -72173 -41242
rect -72477 -41862 -72173 -41858
rect -71477 -41242 -71173 -41238
rect -71477 -41858 -71473 -41242
rect -71473 -41858 -71177 -41242
rect -71177 -41858 -71173 -41242
rect -71477 -41862 -71173 -41858
rect -70477 -41242 -70173 -41238
rect -70477 -41858 -70473 -41242
rect -70473 -41858 -70177 -41242
rect -70177 -41858 -70173 -41242
rect -70477 -41862 -70173 -41858
rect -69477 -41242 -69173 -41238
rect -69477 -41858 -69473 -41242
rect -69473 -41858 -69177 -41242
rect -69177 -41858 -69173 -41242
rect -69477 -41862 -69173 -41858
rect -68477 -41242 -68173 -41238
rect -68477 -41858 -68473 -41242
rect -68473 -41858 -68177 -41242
rect -68177 -41858 -68173 -41242
rect -68477 -41862 -68173 -41858
rect -67477 -41242 -67173 -41238
rect -67477 -41858 -67473 -41242
rect -67473 -41858 -67177 -41242
rect -67177 -41858 -67173 -41242
rect -67477 -41862 -67173 -41858
rect -66477 -41242 -66173 -41238
rect -66477 -41858 -66473 -41242
rect -66473 -41858 -66177 -41242
rect -66177 -41858 -66173 -41242
rect -66477 -41862 -66173 -41858
rect -65477 -41242 -65173 -41238
rect -65477 -41858 -65473 -41242
rect -65473 -41858 -65177 -41242
rect -65177 -41858 -65173 -41242
rect -65477 -41862 -65173 -41858
rect -64477 -41242 -64173 -41238
rect -64477 -41858 -64473 -41242
rect -64473 -41858 -64177 -41242
rect -64177 -41858 -64173 -41242
rect -64477 -41862 -64173 -41858
rect -63477 -41242 -63173 -41238
rect -63477 -41858 -63473 -41242
rect -63473 -41858 -63177 -41242
rect -63177 -41858 -63173 -41242
rect -63477 -41862 -63173 -41858
rect -62477 -41242 -62173 -41238
rect -62477 -41858 -62473 -41242
rect -62473 -41858 -62177 -41242
rect -62177 -41858 -62173 -41242
rect -62477 -41862 -62173 -41858
rect -61477 -41242 -61173 -41238
rect -61477 -41858 -61473 -41242
rect -61473 -41858 -61177 -41242
rect -61177 -41858 -61173 -41242
rect -61477 -41862 -61173 -41858
rect -60477 -41242 -60173 -41238
rect -60477 -41858 -60473 -41242
rect -60473 -41858 -60177 -41242
rect -60177 -41858 -60173 -41242
rect -60477 -41862 -60173 -41858
rect -59477 -41242 -59173 -41238
rect -59477 -41858 -59473 -41242
rect -59473 -41858 -59177 -41242
rect -59177 -41858 -59173 -41242
rect -59477 -41862 -59173 -41858
rect -58477 -41242 -58173 -41238
rect -58477 -41858 -58473 -41242
rect -58473 -41858 -58177 -41242
rect -58177 -41858 -58173 -41242
rect -58477 -41862 -58173 -41858
rect -57477 -41242 -57173 -41238
rect -57477 -41858 -57473 -41242
rect -57473 -41858 -57177 -41242
rect -57177 -41858 -57173 -41242
rect -57477 -41862 -57173 -41858
rect -56477 -41242 -56173 -41238
rect -56477 -41858 -56473 -41242
rect -56473 -41858 -56177 -41242
rect -56177 -41858 -56173 -41242
rect -56477 -41862 -56173 -41858
rect -55477 -41242 -55173 -41238
rect -55477 -41858 -55473 -41242
rect -55473 -41858 -55177 -41242
rect -55177 -41858 -55173 -41242
rect -55477 -41862 -55173 -41858
rect -54477 -41242 -54173 -41238
rect -54477 -41858 -54473 -41242
rect -54473 -41858 -54177 -41242
rect -54177 -41858 -54173 -41242
rect -54477 -41862 -54173 -41858
rect -53477 -41242 -53173 -41238
rect -53477 -41858 -53473 -41242
rect -53473 -41858 -53177 -41242
rect -53177 -41858 -53173 -41242
rect -53477 -41862 -53173 -41858
rect -52477 -41242 -52173 -41238
rect -52477 -41858 -52473 -41242
rect -52473 -41858 -52177 -41242
rect -52177 -41858 -52173 -41242
rect -52477 -41862 -52173 -41858
rect -51477 -41242 -51173 -41238
rect -51477 -41858 -51473 -41242
rect -51473 -41858 -51177 -41242
rect -51177 -41858 -51173 -41242
rect -51477 -41862 -51173 -41858
rect -50477 -41242 -50173 -41238
rect -50477 -41858 -50473 -41242
rect -50473 -41858 -50177 -41242
rect -50177 -41858 -50173 -41242
rect -50477 -41862 -50173 -41858
rect -49477 -41242 -49173 -41238
rect -49477 -41858 -49473 -41242
rect -49473 -41858 -49177 -41242
rect -49177 -41858 -49173 -41242
rect -49477 -41862 -49173 -41858
rect -74817 -41902 -74513 -41898
rect -74817 -42198 -74813 -41902
rect -74813 -42198 -74517 -41902
rect -74517 -42198 -74513 -41902
rect -74817 -42202 -74513 -42198
rect -74477 -41902 -74173 -41898
rect -74477 -42198 -74473 -41902
rect -74473 -42198 -74177 -41902
rect -74177 -42198 -74173 -41902
rect -74477 -42202 -74173 -42198
rect -74137 -41902 -73513 -41898
rect -74137 -42198 -74133 -41902
rect -74133 -42198 -73517 -41902
rect -73517 -42198 -73513 -41902
rect -74137 -42202 -73513 -42198
rect -73477 -41902 -73173 -41898
rect -73477 -42198 -73473 -41902
rect -73473 -42198 -73177 -41902
rect -73177 -42198 -73173 -41902
rect -73477 -42202 -73173 -42198
rect -73137 -41902 -72513 -41898
rect -73137 -42198 -73133 -41902
rect -73133 -42198 -72517 -41902
rect -72517 -42198 -72513 -41902
rect -73137 -42202 -72513 -42198
rect -72477 -41902 -72173 -41898
rect -72477 -42198 -72473 -41902
rect -72473 -42198 -72177 -41902
rect -72177 -42198 -72173 -41902
rect -72477 -42202 -72173 -42198
rect -72137 -41902 -71513 -41898
rect -72137 -42198 -72133 -41902
rect -72133 -42198 -71517 -41902
rect -71517 -42198 -71513 -41902
rect -72137 -42202 -71513 -42198
rect -71477 -41902 -71173 -41898
rect -71477 -42198 -71473 -41902
rect -71473 -42198 -71177 -41902
rect -71177 -42198 -71173 -41902
rect -71477 -42202 -71173 -42198
rect -71137 -41902 -70513 -41898
rect -71137 -42198 -71133 -41902
rect -71133 -42198 -70517 -41902
rect -70517 -42198 -70513 -41902
rect -71137 -42202 -70513 -42198
rect -70477 -41902 -70173 -41898
rect -70477 -42198 -70473 -41902
rect -70473 -42198 -70177 -41902
rect -70177 -42198 -70173 -41902
rect -70477 -42202 -70173 -42198
rect -70137 -41902 -69513 -41898
rect -70137 -42198 -70133 -41902
rect -70133 -42198 -69517 -41902
rect -69517 -42198 -69513 -41902
rect -70137 -42202 -69513 -42198
rect -69477 -41902 -69173 -41898
rect -69477 -42198 -69473 -41902
rect -69473 -42198 -69177 -41902
rect -69177 -42198 -69173 -41902
rect -69477 -42202 -69173 -42198
rect -69137 -41902 -68513 -41898
rect -69137 -42198 -69133 -41902
rect -69133 -42198 -68517 -41902
rect -68517 -42198 -68513 -41902
rect -69137 -42202 -68513 -42198
rect -68477 -41902 -68173 -41898
rect -68477 -42198 -68473 -41902
rect -68473 -42198 -68177 -41902
rect -68177 -42198 -68173 -41902
rect -68477 -42202 -68173 -42198
rect -68137 -41902 -67513 -41898
rect -68137 -42198 -68133 -41902
rect -68133 -42198 -67517 -41902
rect -67517 -42198 -67513 -41902
rect -68137 -42202 -67513 -42198
rect -67477 -41902 -67173 -41898
rect -67477 -42198 -67473 -41902
rect -67473 -42198 -67177 -41902
rect -67177 -42198 -67173 -41902
rect -67477 -42202 -67173 -42198
rect -67137 -41902 -66513 -41898
rect -67137 -42198 -67133 -41902
rect -67133 -42198 -66517 -41902
rect -66517 -42198 -66513 -41902
rect -67137 -42202 -66513 -42198
rect -66477 -41902 -66173 -41898
rect -66477 -42198 -66473 -41902
rect -66473 -42198 -66177 -41902
rect -66177 -42198 -66173 -41902
rect -66477 -42202 -66173 -42198
rect -66137 -41902 -65513 -41898
rect -66137 -42198 -66133 -41902
rect -66133 -42198 -65517 -41902
rect -65517 -42198 -65513 -41902
rect -66137 -42202 -65513 -42198
rect -65477 -41902 -65173 -41898
rect -65477 -42198 -65473 -41902
rect -65473 -42198 -65177 -41902
rect -65177 -42198 -65173 -41902
rect -65477 -42202 -65173 -42198
rect -65137 -41902 -64513 -41898
rect -65137 -42198 -65133 -41902
rect -65133 -42198 -64517 -41902
rect -64517 -42198 -64513 -41902
rect -65137 -42202 -64513 -42198
rect -64477 -41902 -64173 -41898
rect -64477 -42198 -64473 -41902
rect -64473 -42198 -64177 -41902
rect -64177 -42198 -64173 -41902
rect -64477 -42202 -64173 -42198
rect -64137 -41902 -63513 -41898
rect -64137 -42198 -64133 -41902
rect -64133 -42198 -63517 -41902
rect -63517 -42198 -63513 -41902
rect -64137 -42202 -63513 -42198
rect -63477 -41902 -63173 -41898
rect -63477 -42198 -63473 -41902
rect -63473 -42198 -63177 -41902
rect -63177 -42198 -63173 -41902
rect -63477 -42202 -63173 -42198
rect -63137 -41902 -62513 -41898
rect -63137 -42198 -63133 -41902
rect -63133 -42198 -62517 -41902
rect -62517 -42198 -62513 -41902
rect -63137 -42202 -62513 -42198
rect -62477 -41902 -62173 -41898
rect -62477 -42198 -62473 -41902
rect -62473 -42198 -62177 -41902
rect -62177 -42198 -62173 -41902
rect -62477 -42202 -62173 -42198
rect -62137 -41902 -61513 -41898
rect -62137 -42198 -62133 -41902
rect -62133 -42198 -61517 -41902
rect -61517 -42198 -61513 -41902
rect -62137 -42202 -61513 -42198
rect -61477 -41902 -61173 -41898
rect -61477 -42198 -61473 -41902
rect -61473 -42198 -61177 -41902
rect -61177 -42198 -61173 -41902
rect -61477 -42202 -61173 -42198
rect -61137 -41902 -60513 -41898
rect -61137 -42198 -61133 -41902
rect -61133 -42198 -60517 -41902
rect -60517 -42198 -60513 -41902
rect -61137 -42202 -60513 -42198
rect -60477 -41902 -60173 -41898
rect -60477 -42198 -60473 -41902
rect -60473 -42198 -60177 -41902
rect -60177 -42198 -60173 -41902
rect -60477 -42202 -60173 -42198
rect -60137 -41902 -59513 -41898
rect -60137 -42198 -60133 -41902
rect -60133 -42198 -59517 -41902
rect -59517 -42198 -59513 -41902
rect -60137 -42202 -59513 -42198
rect -59477 -41902 -59173 -41898
rect -59477 -42198 -59473 -41902
rect -59473 -42198 -59177 -41902
rect -59177 -42198 -59173 -41902
rect -59477 -42202 -59173 -42198
rect -59137 -41902 -58513 -41898
rect -59137 -42198 -59133 -41902
rect -59133 -42198 -58517 -41902
rect -58517 -42198 -58513 -41902
rect -59137 -42202 -58513 -42198
rect -58477 -41902 -58173 -41898
rect -58477 -42198 -58473 -41902
rect -58473 -42198 -58177 -41902
rect -58177 -42198 -58173 -41902
rect -58477 -42202 -58173 -42198
rect -58137 -41902 -57513 -41898
rect -58137 -42198 -58133 -41902
rect -58133 -42198 -57517 -41902
rect -57517 -42198 -57513 -41902
rect -58137 -42202 -57513 -42198
rect -57477 -41902 -57173 -41898
rect -57477 -42198 -57473 -41902
rect -57473 -42198 -57177 -41902
rect -57177 -42198 -57173 -41902
rect -57477 -42202 -57173 -42198
rect -57137 -41902 -56513 -41898
rect -57137 -42198 -57133 -41902
rect -57133 -42198 -56517 -41902
rect -56517 -42198 -56513 -41902
rect -57137 -42202 -56513 -42198
rect -56477 -41902 -56173 -41898
rect -56477 -42198 -56473 -41902
rect -56473 -42198 -56177 -41902
rect -56177 -42198 -56173 -41902
rect -56477 -42202 -56173 -42198
rect -56137 -41902 -55513 -41898
rect -56137 -42198 -56133 -41902
rect -56133 -42198 -55517 -41902
rect -55517 -42198 -55513 -41902
rect -56137 -42202 -55513 -42198
rect -55477 -41902 -55173 -41898
rect -55477 -42198 -55473 -41902
rect -55473 -42198 -55177 -41902
rect -55177 -42198 -55173 -41902
rect -55477 -42202 -55173 -42198
rect -55137 -41902 -54513 -41898
rect -55137 -42198 -55133 -41902
rect -55133 -42198 -54517 -41902
rect -54517 -42198 -54513 -41902
rect -55137 -42202 -54513 -42198
rect -54477 -41902 -54173 -41898
rect -54477 -42198 -54473 -41902
rect -54473 -42198 -54177 -41902
rect -54177 -42198 -54173 -41902
rect -54477 -42202 -54173 -42198
rect -54137 -41902 -53513 -41898
rect -54137 -42198 -54133 -41902
rect -54133 -42198 -53517 -41902
rect -53517 -42198 -53513 -41902
rect -54137 -42202 -53513 -42198
rect -53477 -41902 -53173 -41898
rect -53477 -42198 -53473 -41902
rect -53473 -42198 -53177 -41902
rect -53177 -42198 -53173 -41902
rect -53477 -42202 -53173 -42198
rect -53137 -41902 -52513 -41898
rect -53137 -42198 -53133 -41902
rect -53133 -42198 -52517 -41902
rect -52517 -42198 -52513 -41902
rect -53137 -42202 -52513 -42198
rect -52477 -41902 -52173 -41898
rect -52477 -42198 -52473 -41902
rect -52473 -42198 -52177 -41902
rect -52177 -42198 -52173 -41902
rect -52477 -42202 -52173 -42198
rect -52137 -41902 -51513 -41898
rect -52137 -42198 -52133 -41902
rect -52133 -42198 -51517 -41902
rect -51517 -42198 -51513 -41902
rect -52137 -42202 -51513 -42198
rect -51477 -41902 -51173 -41898
rect -51477 -42198 -51473 -41902
rect -51473 -42198 -51177 -41902
rect -51177 -42198 -51173 -41902
rect -51477 -42202 -51173 -42198
rect -51137 -41902 -50513 -41898
rect -51137 -42198 -51133 -41902
rect -51133 -42198 -50517 -41902
rect -50517 -42198 -50513 -41902
rect -51137 -42202 -50513 -42198
rect -50477 -41902 -50173 -41898
rect -50477 -42198 -50473 -41902
rect -50473 -42198 -50177 -41902
rect -50177 -42198 -50173 -41902
rect -50477 -42202 -50173 -42198
rect -50137 -41902 -49513 -41898
rect -50137 -42198 -50133 -41902
rect -50133 -42198 -49517 -41902
rect -49517 -42198 -49513 -41902
rect -50137 -42202 -49513 -42198
rect -49477 -41902 -49173 -41898
rect -49477 -42198 -49473 -41902
rect -49473 -42198 -49177 -41902
rect -49177 -42198 -49173 -41902
rect -49477 -42202 -49173 -42198
rect -49137 -41902 -48833 -41898
rect -49137 -42198 -49133 -41902
rect -49133 -42198 -48837 -41902
rect -48837 -42198 -48833 -41902
rect -49137 -42202 -48833 -42198
rect -74477 -42242 -74173 -42238
rect -74477 -42858 -74473 -42242
rect -74473 -42858 -74177 -42242
rect -74177 -42858 -74173 -42242
rect -74477 -42862 -74173 -42858
rect -73477 -42242 -73173 -42238
rect -73477 -42858 -73473 -42242
rect -73473 -42858 -73177 -42242
rect -73177 -42858 -73173 -42242
rect -73477 -42862 -73173 -42858
rect -72477 -42242 -72173 -42238
rect -72477 -42858 -72473 -42242
rect -72473 -42858 -72177 -42242
rect -72177 -42858 -72173 -42242
rect -72477 -42862 -72173 -42858
rect -71477 -42242 -71173 -42238
rect -71477 -42858 -71473 -42242
rect -71473 -42858 -71177 -42242
rect -71177 -42858 -71173 -42242
rect -71477 -42862 -71173 -42858
rect -70477 -42242 -70173 -42238
rect -70477 -42858 -70473 -42242
rect -70473 -42858 -70177 -42242
rect -70177 -42858 -70173 -42242
rect -70477 -42862 -70173 -42858
rect -69477 -42242 -69173 -42238
rect -69477 -42858 -69473 -42242
rect -69473 -42858 -69177 -42242
rect -69177 -42858 -69173 -42242
rect -69477 -42862 -69173 -42858
rect -68477 -42242 -68173 -42238
rect -68477 -42858 -68473 -42242
rect -68473 -42858 -68177 -42242
rect -68177 -42858 -68173 -42242
rect -68477 -42862 -68173 -42858
rect -67477 -42242 -67173 -42238
rect -67477 -42858 -67473 -42242
rect -67473 -42858 -67177 -42242
rect -67177 -42858 -67173 -42242
rect -67477 -42862 -67173 -42858
rect -66477 -42242 -66173 -42238
rect -66477 -42858 -66473 -42242
rect -66473 -42858 -66177 -42242
rect -66177 -42858 -66173 -42242
rect -66477 -42862 -66173 -42858
rect -65477 -42242 -65173 -42238
rect -65477 -42858 -65473 -42242
rect -65473 -42858 -65177 -42242
rect -65177 -42858 -65173 -42242
rect -65477 -42862 -65173 -42858
rect -64477 -42242 -64173 -42238
rect -64477 -42858 -64473 -42242
rect -64473 -42858 -64177 -42242
rect -64177 -42858 -64173 -42242
rect -64477 -42862 -64173 -42858
rect -63477 -42242 -63173 -42238
rect -63477 -42858 -63473 -42242
rect -63473 -42858 -63177 -42242
rect -63177 -42858 -63173 -42242
rect -63477 -42862 -63173 -42858
rect -62477 -42242 -62173 -42238
rect -62477 -42858 -62473 -42242
rect -62473 -42858 -62177 -42242
rect -62177 -42858 -62173 -42242
rect -62477 -42862 -62173 -42858
rect -61477 -42242 -61173 -42238
rect -61477 -42858 -61473 -42242
rect -61473 -42858 -61177 -42242
rect -61177 -42858 -61173 -42242
rect -61477 -42862 -61173 -42858
rect -60477 -42242 -60173 -42238
rect -60477 -42858 -60473 -42242
rect -60473 -42858 -60177 -42242
rect -60177 -42858 -60173 -42242
rect -60477 -42862 -60173 -42858
rect -59477 -42242 -59173 -42238
rect -59477 -42858 -59473 -42242
rect -59473 -42858 -59177 -42242
rect -59177 -42858 -59173 -42242
rect -59477 -42862 -59173 -42858
rect -58477 -42242 -58173 -42238
rect -58477 -42858 -58473 -42242
rect -58473 -42858 -58177 -42242
rect -58177 -42858 -58173 -42242
rect -58477 -42862 -58173 -42858
rect -57477 -42242 -57173 -42238
rect -57477 -42858 -57473 -42242
rect -57473 -42858 -57177 -42242
rect -57177 -42858 -57173 -42242
rect -57477 -42862 -57173 -42858
rect -56477 -42242 -56173 -42238
rect -56477 -42858 -56473 -42242
rect -56473 -42858 -56177 -42242
rect -56177 -42858 -56173 -42242
rect -56477 -42862 -56173 -42858
rect -55477 -42242 -55173 -42238
rect -55477 -42858 -55473 -42242
rect -55473 -42858 -55177 -42242
rect -55177 -42858 -55173 -42242
rect -55477 -42862 -55173 -42858
rect -54477 -42242 -54173 -42238
rect -54477 -42858 -54473 -42242
rect -54473 -42858 -54177 -42242
rect -54177 -42858 -54173 -42242
rect -54477 -42862 -54173 -42858
rect -53477 -42242 -53173 -42238
rect -53477 -42858 -53473 -42242
rect -53473 -42858 -53177 -42242
rect -53177 -42858 -53173 -42242
rect -53477 -42862 -53173 -42858
rect -52477 -42242 -52173 -42238
rect -52477 -42858 -52473 -42242
rect -52473 -42858 -52177 -42242
rect -52177 -42858 -52173 -42242
rect -52477 -42862 -52173 -42858
rect -51477 -42242 -51173 -42238
rect -51477 -42858 -51473 -42242
rect -51473 -42858 -51177 -42242
rect -51177 -42858 -51173 -42242
rect -51477 -42862 -51173 -42858
rect -50477 -42242 -50173 -42238
rect -50477 -42858 -50473 -42242
rect -50473 -42858 -50177 -42242
rect -50177 -42858 -50173 -42242
rect -50477 -42862 -50173 -42858
rect -49477 -42242 -49173 -42238
rect -49477 -42858 -49473 -42242
rect -49473 -42858 -49177 -42242
rect -49177 -42858 -49173 -42242
rect -49477 -42862 -49173 -42858
rect -74817 -42902 -74513 -42898
rect -74817 -43198 -74813 -42902
rect -74813 -43198 -74517 -42902
rect -74517 -43198 -74513 -42902
rect -74817 -43202 -74513 -43198
rect -74477 -42902 -74173 -42898
rect -74477 -43198 -74473 -42902
rect -74473 -43198 -74177 -42902
rect -74177 -43198 -74173 -42902
rect -74477 -43202 -74173 -43198
rect -74137 -42902 -73513 -42898
rect -74137 -43198 -74133 -42902
rect -74133 -43198 -73517 -42902
rect -73517 -43198 -73513 -42902
rect -74137 -43202 -73513 -43198
rect -73477 -42902 -73173 -42898
rect -73477 -43198 -73473 -42902
rect -73473 -43198 -73177 -42902
rect -73177 -43198 -73173 -42902
rect -73477 -43202 -73173 -43198
rect -73137 -42902 -72513 -42898
rect -73137 -43198 -73133 -42902
rect -73133 -43198 -72517 -42902
rect -72517 -43198 -72513 -42902
rect -73137 -43202 -72513 -43198
rect -72477 -42902 -72173 -42898
rect -72477 -43198 -72473 -42902
rect -72473 -43198 -72177 -42902
rect -72177 -43198 -72173 -42902
rect -72477 -43202 -72173 -43198
rect -72137 -42902 -71513 -42898
rect -72137 -43198 -72133 -42902
rect -72133 -43198 -71517 -42902
rect -71517 -43198 -71513 -42902
rect -72137 -43202 -71513 -43198
rect -71477 -42902 -71173 -42898
rect -71477 -43198 -71473 -42902
rect -71473 -43198 -71177 -42902
rect -71177 -43198 -71173 -42902
rect -71477 -43202 -71173 -43198
rect -71137 -42902 -70513 -42898
rect -71137 -43198 -71133 -42902
rect -71133 -43198 -70517 -42902
rect -70517 -43198 -70513 -42902
rect -71137 -43202 -70513 -43198
rect -70477 -42902 -70173 -42898
rect -70477 -43198 -70473 -42902
rect -70473 -43198 -70177 -42902
rect -70177 -43198 -70173 -42902
rect -70477 -43202 -70173 -43198
rect -70137 -42902 -69513 -42898
rect -70137 -43198 -70133 -42902
rect -70133 -43198 -69517 -42902
rect -69517 -43198 -69513 -42902
rect -70137 -43202 -69513 -43198
rect -69477 -42902 -69173 -42898
rect -69477 -43198 -69473 -42902
rect -69473 -43198 -69177 -42902
rect -69177 -43198 -69173 -42902
rect -69477 -43202 -69173 -43198
rect -69137 -42902 -68513 -42898
rect -69137 -43198 -69133 -42902
rect -69133 -43198 -68517 -42902
rect -68517 -43198 -68513 -42902
rect -69137 -43202 -68513 -43198
rect -68477 -42902 -68173 -42898
rect -68477 -43198 -68473 -42902
rect -68473 -43198 -68177 -42902
rect -68177 -43198 -68173 -42902
rect -68477 -43202 -68173 -43198
rect -68137 -42902 -67513 -42898
rect -68137 -43198 -68133 -42902
rect -68133 -43198 -67517 -42902
rect -67517 -43198 -67513 -42902
rect -68137 -43202 -67513 -43198
rect -67477 -42902 -67173 -42898
rect -67477 -43198 -67473 -42902
rect -67473 -43198 -67177 -42902
rect -67177 -43198 -67173 -42902
rect -67477 -43202 -67173 -43198
rect -67137 -42902 -66513 -42898
rect -67137 -43198 -67133 -42902
rect -67133 -43198 -66517 -42902
rect -66517 -43198 -66513 -42902
rect -67137 -43202 -66513 -43198
rect -66477 -42902 -66173 -42898
rect -66477 -43198 -66473 -42902
rect -66473 -43198 -66177 -42902
rect -66177 -43198 -66173 -42902
rect -66477 -43202 -66173 -43198
rect -66137 -42902 -65513 -42898
rect -66137 -43198 -66133 -42902
rect -66133 -43198 -65517 -42902
rect -65517 -43198 -65513 -42902
rect -66137 -43202 -65513 -43198
rect -65477 -42902 -65173 -42898
rect -65477 -43198 -65473 -42902
rect -65473 -43198 -65177 -42902
rect -65177 -43198 -65173 -42902
rect -65477 -43202 -65173 -43198
rect -65137 -42902 -64513 -42898
rect -65137 -43198 -65133 -42902
rect -65133 -43198 -64517 -42902
rect -64517 -43198 -64513 -42902
rect -65137 -43202 -64513 -43198
rect -64477 -42902 -64173 -42898
rect -64477 -43198 -64473 -42902
rect -64473 -43198 -64177 -42902
rect -64177 -43198 -64173 -42902
rect -64477 -43202 -64173 -43198
rect -64137 -42902 -63513 -42898
rect -64137 -43198 -64133 -42902
rect -64133 -43198 -63517 -42902
rect -63517 -43198 -63513 -42902
rect -64137 -43202 -63513 -43198
rect -63477 -42902 -63173 -42898
rect -63477 -43198 -63473 -42902
rect -63473 -43198 -63177 -42902
rect -63177 -43198 -63173 -42902
rect -63477 -43202 -63173 -43198
rect -63137 -42902 -62513 -42898
rect -63137 -43198 -63133 -42902
rect -63133 -43198 -62517 -42902
rect -62517 -43198 -62513 -42902
rect -63137 -43202 -62513 -43198
rect -62477 -42902 -62173 -42898
rect -62477 -43198 -62473 -42902
rect -62473 -43198 -62177 -42902
rect -62177 -43198 -62173 -42902
rect -62477 -43202 -62173 -43198
rect -62137 -42902 -61513 -42898
rect -62137 -43198 -62133 -42902
rect -62133 -43198 -61517 -42902
rect -61517 -43198 -61513 -42902
rect -62137 -43202 -61513 -43198
rect -61477 -42902 -61173 -42898
rect -61477 -43198 -61473 -42902
rect -61473 -43198 -61177 -42902
rect -61177 -43198 -61173 -42902
rect -61477 -43202 -61173 -43198
rect -61137 -42902 -60513 -42898
rect -61137 -43198 -61133 -42902
rect -61133 -43198 -60517 -42902
rect -60517 -43198 -60513 -42902
rect -61137 -43202 -60513 -43198
rect -60477 -42902 -60173 -42898
rect -60477 -43198 -60473 -42902
rect -60473 -43198 -60177 -42902
rect -60177 -43198 -60173 -42902
rect -60477 -43202 -60173 -43198
rect -60137 -42902 -59513 -42898
rect -60137 -43198 -60133 -42902
rect -60133 -43198 -59517 -42902
rect -59517 -43198 -59513 -42902
rect -60137 -43202 -59513 -43198
rect -59477 -42902 -59173 -42898
rect -59477 -43198 -59473 -42902
rect -59473 -43198 -59177 -42902
rect -59177 -43198 -59173 -42902
rect -59477 -43202 -59173 -43198
rect -59137 -42902 -58513 -42898
rect -59137 -43198 -59133 -42902
rect -59133 -43198 -58517 -42902
rect -58517 -43198 -58513 -42902
rect -59137 -43202 -58513 -43198
rect -58477 -42902 -58173 -42898
rect -58477 -43198 -58473 -42902
rect -58473 -43198 -58177 -42902
rect -58177 -43198 -58173 -42902
rect -58477 -43202 -58173 -43198
rect -58137 -42902 -57513 -42898
rect -58137 -43198 -58133 -42902
rect -58133 -43198 -57517 -42902
rect -57517 -43198 -57513 -42902
rect -58137 -43202 -57513 -43198
rect -57477 -42902 -57173 -42898
rect -57477 -43198 -57473 -42902
rect -57473 -43198 -57177 -42902
rect -57177 -43198 -57173 -42902
rect -57477 -43202 -57173 -43198
rect -57137 -42902 -56513 -42898
rect -57137 -43198 -57133 -42902
rect -57133 -43198 -56517 -42902
rect -56517 -43198 -56513 -42902
rect -57137 -43202 -56513 -43198
rect -56477 -42902 -56173 -42898
rect -56477 -43198 -56473 -42902
rect -56473 -43198 -56177 -42902
rect -56177 -43198 -56173 -42902
rect -56477 -43202 -56173 -43198
rect -56137 -42902 -55513 -42898
rect -56137 -43198 -56133 -42902
rect -56133 -43198 -55517 -42902
rect -55517 -43198 -55513 -42902
rect -56137 -43202 -55513 -43198
rect -55477 -42902 -55173 -42898
rect -55477 -43198 -55473 -42902
rect -55473 -43198 -55177 -42902
rect -55177 -43198 -55173 -42902
rect -55477 -43202 -55173 -43198
rect -55137 -42902 -54513 -42898
rect -55137 -43198 -55133 -42902
rect -55133 -43198 -54517 -42902
rect -54517 -43198 -54513 -42902
rect -55137 -43202 -54513 -43198
rect -54477 -42902 -54173 -42898
rect -54477 -43198 -54473 -42902
rect -54473 -43198 -54177 -42902
rect -54177 -43198 -54173 -42902
rect -54477 -43202 -54173 -43198
rect -54137 -42902 -53513 -42898
rect -54137 -43198 -54133 -42902
rect -54133 -43198 -53517 -42902
rect -53517 -43198 -53513 -42902
rect -54137 -43202 -53513 -43198
rect -53477 -42902 -53173 -42898
rect -53477 -43198 -53473 -42902
rect -53473 -43198 -53177 -42902
rect -53177 -43198 -53173 -42902
rect -53477 -43202 -53173 -43198
rect -53137 -42902 -52513 -42898
rect -53137 -43198 -53133 -42902
rect -53133 -43198 -52517 -42902
rect -52517 -43198 -52513 -42902
rect -53137 -43202 -52513 -43198
rect -52477 -42902 -52173 -42898
rect -52477 -43198 -52473 -42902
rect -52473 -43198 -52177 -42902
rect -52177 -43198 -52173 -42902
rect -52477 -43202 -52173 -43198
rect -52137 -42902 -51513 -42898
rect -52137 -43198 -52133 -42902
rect -52133 -43198 -51517 -42902
rect -51517 -43198 -51513 -42902
rect -52137 -43202 -51513 -43198
rect -51477 -42902 -51173 -42898
rect -51477 -43198 -51473 -42902
rect -51473 -43198 -51177 -42902
rect -51177 -43198 -51173 -42902
rect -51477 -43202 -51173 -43198
rect -51137 -42902 -50513 -42898
rect -51137 -43198 -51133 -42902
rect -51133 -43198 -50517 -42902
rect -50517 -43198 -50513 -42902
rect -51137 -43202 -50513 -43198
rect -50477 -42902 -50173 -42898
rect -50477 -43198 -50473 -42902
rect -50473 -43198 -50177 -42902
rect -50177 -43198 -50173 -42902
rect -50477 -43202 -50173 -43198
rect -50137 -42902 -49513 -42898
rect -50137 -43198 -50133 -42902
rect -50133 -43198 -49517 -42902
rect -49517 -43198 -49513 -42902
rect -50137 -43202 -49513 -43198
rect -49477 -42902 -49173 -42898
rect -49477 -43198 -49473 -42902
rect -49473 -43198 -49177 -42902
rect -49177 -43198 -49173 -42902
rect -49477 -43202 -49173 -43198
rect -49137 -42902 -48833 -42898
rect -49137 -43198 -49133 -42902
rect -49133 -43198 -48837 -42902
rect -48837 -43198 -48833 -42902
rect -49137 -43202 -48833 -43198
rect -74477 -43242 -74173 -43238
rect -74477 -43858 -74473 -43242
rect -74473 -43858 -74177 -43242
rect -74177 -43858 -74173 -43242
rect -74477 -43862 -74173 -43858
rect -73477 -43242 -73173 -43238
rect -73477 -43858 -73473 -43242
rect -73473 -43858 -73177 -43242
rect -73177 -43858 -73173 -43242
rect -73477 -43862 -73173 -43858
rect -72477 -43242 -72173 -43238
rect -72477 -43858 -72473 -43242
rect -72473 -43858 -72177 -43242
rect -72177 -43858 -72173 -43242
rect -72477 -43862 -72173 -43858
rect -71477 -43242 -71173 -43238
rect -71477 -43858 -71473 -43242
rect -71473 -43858 -71177 -43242
rect -71177 -43858 -71173 -43242
rect -71477 -43862 -71173 -43858
rect -70477 -43242 -70173 -43238
rect -70477 -43858 -70473 -43242
rect -70473 -43858 -70177 -43242
rect -70177 -43858 -70173 -43242
rect -70477 -43862 -70173 -43858
rect -69477 -43242 -69173 -43238
rect -69477 -43858 -69473 -43242
rect -69473 -43858 -69177 -43242
rect -69177 -43858 -69173 -43242
rect -69477 -43862 -69173 -43858
rect -68477 -43242 -68173 -43238
rect -68477 -43858 -68473 -43242
rect -68473 -43858 -68177 -43242
rect -68177 -43858 -68173 -43242
rect -68477 -43862 -68173 -43858
rect -67477 -43242 -67173 -43238
rect -67477 -43858 -67473 -43242
rect -67473 -43858 -67177 -43242
rect -67177 -43858 -67173 -43242
rect -67477 -43862 -67173 -43858
rect -66477 -43242 -66173 -43238
rect -66477 -43858 -66473 -43242
rect -66473 -43858 -66177 -43242
rect -66177 -43858 -66173 -43242
rect -66477 -43862 -66173 -43858
rect -65477 -43242 -65173 -43238
rect -65477 -43858 -65473 -43242
rect -65473 -43858 -65177 -43242
rect -65177 -43858 -65173 -43242
rect -65477 -43862 -65173 -43858
rect -64477 -43242 -64173 -43238
rect -64477 -43858 -64473 -43242
rect -64473 -43858 -64177 -43242
rect -64177 -43858 -64173 -43242
rect -64477 -43862 -64173 -43858
rect -63477 -43242 -63173 -43238
rect -63477 -43858 -63473 -43242
rect -63473 -43858 -63177 -43242
rect -63177 -43858 -63173 -43242
rect -63477 -43862 -63173 -43858
rect -62477 -43242 -62173 -43238
rect -62477 -43858 -62473 -43242
rect -62473 -43858 -62177 -43242
rect -62177 -43858 -62173 -43242
rect -62477 -43862 -62173 -43858
rect -61477 -43242 -61173 -43238
rect -61477 -43858 -61473 -43242
rect -61473 -43858 -61177 -43242
rect -61177 -43858 -61173 -43242
rect -61477 -43862 -61173 -43858
rect -60477 -43242 -60173 -43238
rect -60477 -43858 -60473 -43242
rect -60473 -43858 -60177 -43242
rect -60177 -43858 -60173 -43242
rect -60477 -43862 -60173 -43858
rect -59477 -43242 -59173 -43238
rect -59477 -43858 -59473 -43242
rect -59473 -43858 -59177 -43242
rect -59177 -43858 -59173 -43242
rect -59477 -43862 -59173 -43858
rect -58477 -43242 -58173 -43238
rect -58477 -43858 -58473 -43242
rect -58473 -43858 -58177 -43242
rect -58177 -43858 -58173 -43242
rect -58477 -43862 -58173 -43858
rect -57477 -43242 -57173 -43238
rect -57477 -43858 -57473 -43242
rect -57473 -43858 -57177 -43242
rect -57177 -43858 -57173 -43242
rect -57477 -43862 -57173 -43858
rect -56477 -43242 -56173 -43238
rect -56477 -43858 -56473 -43242
rect -56473 -43858 -56177 -43242
rect -56177 -43858 -56173 -43242
rect -56477 -43862 -56173 -43858
rect -55477 -43242 -55173 -43238
rect -55477 -43858 -55473 -43242
rect -55473 -43858 -55177 -43242
rect -55177 -43858 -55173 -43242
rect -55477 -43862 -55173 -43858
rect -54477 -43242 -54173 -43238
rect -54477 -43858 -54473 -43242
rect -54473 -43858 -54177 -43242
rect -54177 -43858 -54173 -43242
rect -54477 -43862 -54173 -43858
rect -53477 -43242 -53173 -43238
rect -53477 -43858 -53473 -43242
rect -53473 -43858 -53177 -43242
rect -53177 -43858 -53173 -43242
rect -53477 -43862 -53173 -43858
rect -52477 -43242 -52173 -43238
rect -52477 -43858 -52473 -43242
rect -52473 -43858 -52177 -43242
rect -52177 -43858 -52173 -43242
rect -52477 -43862 -52173 -43858
rect -51477 -43242 -51173 -43238
rect -51477 -43858 -51473 -43242
rect -51473 -43858 -51177 -43242
rect -51177 -43858 -51173 -43242
rect -51477 -43862 -51173 -43858
rect -50477 -43242 -50173 -43238
rect -50477 -43858 -50473 -43242
rect -50473 -43858 -50177 -43242
rect -50177 -43858 -50173 -43242
rect -50477 -43862 -50173 -43858
rect -49477 -43242 -49173 -43238
rect -49477 -43858 -49473 -43242
rect -49473 -43858 -49177 -43242
rect -49177 -43858 -49173 -43242
rect -49477 -43862 -49173 -43858
rect -74817 -43902 -74513 -43898
rect -74817 -44198 -74813 -43902
rect -74813 -44198 -74517 -43902
rect -74517 -44198 -74513 -43902
rect -74817 -44202 -74513 -44198
rect -74477 -43902 -74173 -43898
rect -74477 -44198 -74473 -43902
rect -74473 -44198 -74177 -43902
rect -74177 -44198 -74173 -43902
rect -74477 -44202 -74173 -44198
rect -74137 -43902 -73513 -43898
rect -74137 -44198 -74133 -43902
rect -74133 -44198 -73517 -43902
rect -73517 -44198 -73513 -43902
rect -74137 -44202 -73513 -44198
rect -73477 -43902 -73173 -43898
rect -73477 -44198 -73473 -43902
rect -73473 -44198 -73177 -43902
rect -73177 -44198 -73173 -43902
rect -73477 -44202 -73173 -44198
rect -73137 -43902 -72513 -43898
rect -73137 -44198 -73133 -43902
rect -73133 -44198 -72517 -43902
rect -72517 -44198 -72513 -43902
rect -73137 -44202 -72513 -44198
rect -72477 -43902 -72173 -43898
rect -72477 -44198 -72473 -43902
rect -72473 -44198 -72177 -43902
rect -72177 -44198 -72173 -43902
rect -72477 -44202 -72173 -44198
rect -72137 -43902 -71513 -43898
rect -72137 -44198 -72133 -43902
rect -72133 -44198 -71517 -43902
rect -71517 -44198 -71513 -43902
rect -72137 -44202 -71513 -44198
rect -71477 -43902 -71173 -43898
rect -71477 -44198 -71473 -43902
rect -71473 -44198 -71177 -43902
rect -71177 -44198 -71173 -43902
rect -71477 -44202 -71173 -44198
rect -71137 -43902 -70513 -43898
rect -71137 -44198 -71133 -43902
rect -71133 -44198 -70517 -43902
rect -70517 -44198 -70513 -43902
rect -71137 -44202 -70513 -44198
rect -70477 -43902 -70173 -43898
rect -70477 -44198 -70473 -43902
rect -70473 -44198 -70177 -43902
rect -70177 -44198 -70173 -43902
rect -70477 -44202 -70173 -44198
rect -70137 -43902 -69513 -43898
rect -70137 -44198 -70133 -43902
rect -70133 -44198 -69517 -43902
rect -69517 -44198 -69513 -43902
rect -70137 -44202 -69513 -44198
rect -69477 -43902 -69173 -43898
rect -69477 -44198 -69473 -43902
rect -69473 -44198 -69177 -43902
rect -69177 -44198 -69173 -43902
rect -69477 -44202 -69173 -44198
rect -69137 -43902 -68513 -43898
rect -69137 -44198 -69133 -43902
rect -69133 -44198 -68517 -43902
rect -68517 -44198 -68513 -43902
rect -69137 -44202 -68513 -44198
rect -68477 -43902 -68173 -43898
rect -68477 -44198 -68473 -43902
rect -68473 -44198 -68177 -43902
rect -68177 -44198 -68173 -43902
rect -68477 -44202 -68173 -44198
rect -68137 -43902 -67513 -43898
rect -68137 -44198 -68133 -43902
rect -68133 -44198 -67517 -43902
rect -67517 -44198 -67513 -43902
rect -68137 -44202 -67513 -44198
rect -67477 -43902 -67173 -43898
rect -67477 -44198 -67473 -43902
rect -67473 -44198 -67177 -43902
rect -67177 -44198 -67173 -43902
rect -67477 -44202 -67173 -44198
rect -67137 -43902 -66513 -43898
rect -67137 -44198 -67133 -43902
rect -67133 -44198 -66517 -43902
rect -66517 -44198 -66513 -43902
rect -67137 -44202 -66513 -44198
rect -66477 -43902 -66173 -43898
rect -66477 -44198 -66473 -43902
rect -66473 -44198 -66177 -43902
rect -66177 -44198 -66173 -43902
rect -66477 -44202 -66173 -44198
rect -66137 -43902 -65513 -43898
rect -66137 -44198 -66133 -43902
rect -66133 -44198 -65517 -43902
rect -65517 -44198 -65513 -43902
rect -66137 -44202 -65513 -44198
rect -65477 -43902 -65173 -43898
rect -65477 -44198 -65473 -43902
rect -65473 -44198 -65177 -43902
rect -65177 -44198 -65173 -43902
rect -65477 -44202 -65173 -44198
rect -65137 -43902 -64513 -43898
rect -65137 -44198 -65133 -43902
rect -65133 -44198 -64517 -43902
rect -64517 -44198 -64513 -43902
rect -65137 -44202 -64513 -44198
rect -64477 -43902 -64173 -43898
rect -64477 -44198 -64473 -43902
rect -64473 -44198 -64177 -43902
rect -64177 -44198 -64173 -43902
rect -64477 -44202 -64173 -44198
rect -64137 -43902 -63513 -43898
rect -64137 -44198 -64133 -43902
rect -64133 -44198 -63517 -43902
rect -63517 -44198 -63513 -43902
rect -64137 -44202 -63513 -44198
rect -63477 -43902 -63173 -43898
rect -63477 -44198 -63473 -43902
rect -63473 -44198 -63177 -43902
rect -63177 -44198 -63173 -43902
rect -63477 -44202 -63173 -44198
rect -63137 -43902 -62513 -43898
rect -63137 -44198 -63133 -43902
rect -63133 -44198 -62517 -43902
rect -62517 -44198 -62513 -43902
rect -63137 -44202 -62513 -44198
rect -62477 -43902 -62173 -43898
rect -62477 -44198 -62473 -43902
rect -62473 -44198 -62177 -43902
rect -62177 -44198 -62173 -43902
rect -62477 -44202 -62173 -44198
rect -62137 -43902 -61513 -43898
rect -62137 -44198 -62133 -43902
rect -62133 -44198 -61517 -43902
rect -61517 -44198 -61513 -43902
rect -62137 -44202 -61513 -44198
rect -61477 -43902 -61173 -43898
rect -61477 -44198 -61473 -43902
rect -61473 -44198 -61177 -43902
rect -61177 -44198 -61173 -43902
rect -61477 -44202 -61173 -44198
rect -61137 -43902 -60513 -43898
rect -61137 -44198 -61133 -43902
rect -61133 -44198 -60517 -43902
rect -60517 -44198 -60513 -43902
rect -61137 -44202 -60513 -44198
rect -60477 -43902 -60173 -43898
rect -60477 -44198 -60473 -43902
rect -60473 -44198 -60177 -43902
rect -60177 -44198 -60173 -43902
rect -60477 -44202 -60173 -44198
rect -60137 -43902 -59513 -43898
rect -60137 -44198 -60133 -43902
rect -60133 -44198 -59517 -43902
rect -59517 -44198 -59513 -43902
rect -60137 -44202 -59513 -44198
rect -59477 -43902 -59173 -43898
rect -59477 -44198 -59473 -43902
rect -59473 -44198 -59177 -43902
rect -59177 -44198 -59173 -43902
rect -59477 -44202 -59173 -44198
rect -59137 -43902 -58513 -43898
rect -59137 -44198 -59133 -43902
rect -59133 -44198 -58517 -43902
rect -58517 -44198 -58513 -43902
rect -59137 -44202 -58513 -44198
rect -58477 -43902 -58173 -43898
rect -58477 -44198 -58473 -43902
rect -58473 -44198 -58177 -43902
rect -58177 -44198 -58173 -43902
rect -58477 -44202 -58173 -44198
rect -58137 -43902 -57513 -43898
rect -58137 -44198 -58133 -43902
rect -58133 -44198 -57517 -43902
rect -57517 -44198 -57513 -43902
rect -58137 -44202 -57513 -44198
rect -57477 -43902 -57173 -43898
rect -57477 -44198 -57473 -43902
rect -57473 -44198 -57177 -43902
rect -57177 -44198 -57173 -43902
rect -57477 -44202 -57173 -44198
rect -57137 -43902 -56513 -43898
rect -57137 -44198 -57133 -43902
rect -57133 -44198 -56517 -43902
rect -56517 -44198 -56513 -43902
rect -57137 -44202 -56513 -44198
rect -56477 -43902 -56173 -43898
rect -56477 -44198 -56473 -43902
rect -56473 -44198 -56177 -43902
rect -56177 -44198 -56173 -43902
rect -56477 -44202 -56173 -44198
rect -56137 -43902 -55513 -43898
rect -56137 -44198 -56133 -43902
rect -56133 -44198 -55517 -43902
rect -55517 -44198 -55513 -43902
rect -56137 -44202 -55513 -44198
rect -55477 -43902 -55173 -43898
rect -55477 -44198 -55473 -43902
rect -55473 -44198 -55177 -43902
rect -55177 -44198 -55173 -43902
rect -55477 -44202 -55173 -44198
rect -55137 -43902 -54513 -43898
rect -55137 -44198 -55133 -43902
rect -55133 -44198 -54517 -43902
rect -54517 -44198 -54513 -43902
rect -55137 -44202 -54513 -44198
rect -54477 -43902 -54173 -43898
rect -54477 -44198 -54473 -43902
rect -54473 -44198 -54177 -43902
rect -54177 -44198 -54173 -43902
rect -54477 -44202 -54173 -44198
rect -54137 -43902 -53513 -43898
rect -54137 -44198 -54133 -43902
rect -54133 -44198 -53517 -43902
rect -53517 -44198 -53513 -43902
rect -54137 -44202 -53513 -44198
rect -53477 -43902 -53173 -43898
rect -53477 -44198 -53473 -43902
rect -53473 -44198 -53177 -43902
rect -53177 -44198 -53173 -43902
rect -53477 -44202 -53173 -44198
rect -53137 -43902 -52513 -43898
rect -53137 -44198 -53133 -43902
rect -53133 -44198 -52517 -43902
rect -52517 -44198 -52513 -43902
rect -53137 -44202 -52513 -44198
rect -52477 -43902 -52173 -43898
rect -52477 -44198 -52473 -43902
rect -52473 -44198 -52177 -43902
rect -52177 -44198 -52173 -43902
rect -52477 -44202 -52173 -44198
rect -52137 -43902 -51513 -43898
rect -52137 -44198 -52133 -43902
rect -52133 -44198 -51517 -43902
rect -51517 -44198 -51513 -43902
rect -52137 -44202 -51513 -44198
rect -51477 -43902 -51173 -43898
rect -51477 -44198 -51473 -43902
rect -51473 -44198 -51177 -43902
rect -51177 -44198 -51173 -43902
rect -51477 -44202 -51173 -44198
rect -51137 -43902 -50513 -43898
rect -51137 -44198 -51133 -43902
rect -51133 -44198 -50517 -43902
rect -50517 -44198 -50513 -43902
rect -51137 -44202 -50513 -44198
rect -50477 -43902 -50173 -43898
rect -50477 -44198 -50473 -43902
rect -50473 -44198 -50177 -43902
rect -50177 -44198 -50173 -43902
rect -50477 -44202 -50173 -44198
rect -50137 -43902 -49513 -43898
rect -50137 -44198 -50133 -43902
rect -50133 -44198 -49517 -43902
rect -49517 -44198 -49513 -43902
rect -50137 -44202 -49513 -44198
rect -49477 -43902 -49173 -43898
rect -49477 -44198 -49473 -43902
rect -49473 -44198 -49177 -43902
rect -49177 -44198 -49173 -43902
rect -49477 -44202 -49173 -44198
rect -49137 -43902 -48833 -43898
rect -49137 -44198 -49133 -43902
rect -49133 -44198 -48837 -43902
rect -48837 -44198 -48833 -43902
rect -49137 -44202 -48833 -44198
rect -74477 -44242 -74173 -44238
rect -74477 -44858 -74473 -44242
rect -74473 -44858 -74177 -44242
rect -74177 -44858 -74173 -44242
rect -74477 -44862 -74173 -44858
rect -73477 -44242 -73173 -44238
rect -73477 -44858 -73473 -44242
rect -73473 -44858 -73177 -44242
rect -73177 -44858 -73173 -44242
rect -73477 -44862 -73173 -44858
rect -72477 -44242 -72173 -44238
rect -72477 -44858 -72473 -44242
rect -72473 -44858 -72177 -44242
rect -72177 -44858 -72173 -44242
rect -72477 -44862 -72173 -44858
rect -71477 -44242 -71173 -44238
rect -71477 -44858 -71473 -44242
rect -71473 -44858 -71177 -44242
rect -71177 -44858 -71173 -44242
rect -71477 -44862 -71173 -44858
rect -70477 -44242 -70173 -44238
rect -70477 -44858 -70473 -44242
rect -70473 -44858 -70177 -44242
rect -70177 -44858 -70173 -44242
rect -70477 -44862 -70173 -44858
rect -69477 -44242 -69173 -44238
rect -69477 -44858 -69473 -44242
rect -69473 -44858 -69177 -44242
rect -69177 -44858 -69173 -44242
rect -69477 -44862 -69173 -44858
rect -68477 -44242 -68173 -44238
rect -68477 -44858 -68473 -44242
rect -68473 -44858 -68177 -44242
rect -68177 -44858 -68173 -44242
rect -68477 -44862 -68173 -44858
rect -67477 -44242 -67173 -44238
rect -67477 -44858 -67473 -44242
rect -67473 -44858 -67177 -44242
rect -67177 -44858 -67173 -44242
rect -67477 -44862 -67173 -44858
rect -66477 -44242 -66173 -44238
rect -66477 -44858 -66473 -44242
rect -66473 -44858 -66177 -44242
rect -66177 -44858 -66173 -44242
rect -66477 -44862 -66173 -44858
rect -65477 -44242 -65173 -44238
rect -65477 -44858 -65473 -44242
rect -65473 -44858 -65177 -44242
rect -65177 -44858 -65173 -44242
rect -65477 -44862 -65173 -44858
rect -64477 -44242 -64173 -44238
rect -64477 -44858 -64473 -44242
rect -64473 -44858 -64177 -44242
rect -64177 -44858 -64173 -44242
rect -64477 -44862 -64173 -44858
rect -63477 -44242 -63173 -44238
rect -63477 -44858 -63473 -44242
rect -63473 -44858 -63177 -44242
rect -63177 -44858 -63173 -44242
rect -63477 -44862 -63173 -44858
rect -62477 -44242 -62173 -44238
rect -62477 -44858 -62473 -44242
rect -62473 -44858 -62177 -44242
rect -62177 -44858 -62173 -44242
rect -62477 -44862 -62173 -44858
rect -61477 -44242 -61173 -44238
rect -61477 -44858 -61473 -44242
rect -61473 -44858 -61177 -44242
rect -61177 -44858 -61173 -44242
rect -61477 -44862 -61173 -44858
rect -60477 -44242 -60173 -44238
rect -60477 -44858 -60473 -44242
rect -60473 -44858 -60177 -44242
rect -60177 -44858 -60173 -44242
rect -60477 -44862 -60173 -44858
rect -59477 -44242 -59173 -44238
rect -59477 -44858 -59473 -44242
rect -59473 -44858 -59177 -44242
rect -59177 -44858 -59173 -44242
rect -59477 -44862 -59173 -44858
rect -58477 -44242 -58173 -44238
rect -58477 -44858 -58473 -44242
rect -58473 -44858 -58177 -44242
rect -58177 -44858 -58173 -44242
rect -58477 -44862 -58173 -44858
rect -57477 -44242 -57173 -44238
rect -57477 -44858 -57473 -44242
rect -57473 -44858 -57177 -44242
rect -57177 -44858 -57173 -44242
rect -57477 -44862 -57173 -44858
rect -56477 -44242 -56173 -44238
rect -56477 -44858 -56473 -44242
rect -56473 -44858 -56177 -44242
rect -56177 -44858 -56173 -44242
rect -56477 -44862 -56173 -44858
rect -55477 -44242 -55173 -44238
rect -55477 -44858 -55473 -44242
rect -55473 -44858 -55177 -44242
rect -55177 -44858 -55173 -44242
rect -55477 -44862 -55173 -44858
rect -54477 -44242 -54173 -44238
rect -54477 -44858 -54473 -44242
rect -54473 -44858 -54177 -44242
rect -54177 -44858 -54173 -44242
rect -54477 -44862 -54173 -44858
rect -53477 -44242 -53173 -44238
rect -53477 -44858 -53473 -44242
rect -53473 -44858 -53177 -44242
rect -53177 -44858 -53173 -44242
rect -53477 -44862 -53173 -44858
rect -52477 -44242 -52173 -44238
rect -52477 -44858 -52473 -44242
rect -52473 -44858 -52177 -44242
rect -52177 -44858 -52173 -44242
rect -52477 -44862 -52173 -44858
rect -51477 -44242 -51173 -44238
rect -51477 -44858 -51473 -44242
rect -51473 -44858 -51177 -44242
rect -51177 -44858 -51173 -44242
rect -51477 -44862 -51173 -44858
rect -50477 -44242 -50173 -44238
rect -50477 -44858 -50473 -44242
rect -50473 -44858 -50177 -44242
rect -50177 -44858 -50173 -44242
rect -50477 -44862 -50173 -44858
rect -49477 -44242 -49173 -44238
rect -49477 -44858 -49473 -44242
rect -49473 -44858 -49177 -44242
rect -49177 -44858 -49173 -44242
rect -49477 -44862 -49173 -44858
rect -46232 -32602 -36328 -32598
rect -46232 -44498 -46228 -32602
rect -46228 -44498 -36332 -32602
rect -36332 -44498 -36328 -32602
rect -46232 -44502 -36328 -44498
rect -4232 -32602 5672 -32598
rect -4232 -44498 -4228 -32602
rect -4228 -44498 5668 -32602
rect 5668 -44498 5672 -32602
rect -4232 -44502 5672 -44498
rect 8623 -32242 8927 -32238
rect 8623 -32858 8627 -32242
rect 8627 -32858 8923 -32242
rect 8923 -32858 8927 -32242
rect 8623 -32862 8927 -32858
rect 9623 -32242 9927 -32238
rect 9623 -32858 9627 -32242
rect 9627 -32858 9923 -32242
rect 9923 -32858 9927 -32242
rect 9623 -32862 9927 -32858
rect 10623 -32242 10927 -32238
rect 10623 -32858 10627 -32242
rect 10627 -32858 10923 -32242
rect 10923 -32858 10927 -32242
rect 10623 -32862 10927 -32858
rect 11623 -32242 11927 -32238
rect 11623 -32858 11627 -32242
rect 11627 -32858 11923 -32242
rect 11923 -32858 11927 -32242
rect 11623 -32862 11927 -32858
rect 12623 -32242 12927 -32238
rect 12623 -32858 12627 -32242
rect 12627 -32858 12923 -32242
rect 12923 -32858 12927 -32242
rect 12623 -32862 12927 -32858
rect 13623 -32242 13927 -32238
rect 13623 -32858 13627 -32242
rect 13627 -32858 13923 -32242
rect 13923 -32858 13927 -32242
rect 13623 -32862 13927 -32858
rect 14623 -32242 14927 -32238
rect 14623 -32858 14627 -32242
rect 14627 -32858 14923 -32242
rect 14923 -32858 14927 -32242
rect 14623 -32862 14927 -32858
rect 15623 -32242 15927 -32238
rect 15623 -32858 15627 -32242
rect 15627 -32858 15923 -32242
rect 15923 -32858 15927 -32242
rect 15623 -32862 15927 -32858
rect 16623 -32242 16927 -32238
rect 16623 -32858 16627 -32242
rect 16627 -32858 16923 -32242
rect 16923 -32858 16927 -32242
rect 16623 -32862 16927 -32858
rect 17623 -32242 17927 -32238
rect 17623 -32858 17627 -32242
rect 17627 -32858 17923 -32242
rect 17923 -32858 17927 -32242
rect 17623 -32862 17927 -32858
rect 18623 -32242 18927 -32238
rect 18623 -32858 18627 -32242
rect 18627 -32858 18923 -32242
rect 18923 -32858 18927 -32242
rect 18623 -32862 18927 -32858
rect 19623 -32242 19927 -32238
rect 19623 -32858 19627 -32242
rect 19627 -32858 19923 -32242
rect 19923 -32858 19927 -32242
rect 19623 -32862 19927 -32858
rect 20623 -32242 20927 -32238
rect 20623 -32858 20627 -32242
rect 20627 -32858 20923 -32242
rect 20923 -32858 20927 -32242
rect 20623 -32862 20927 -32858
rect 21623 -32242 21927 -32238
rect 21623 -32858 21627 -32242
rect 21627 -32858 21923 -32242
rect 21923 -32858 21927 -32242
rect 21623 -32862 21927 -32858
rect 22623 -32242 22927 -32238
rect 22623 -32858 22627 -32242
rect 22627 -32858 22923 -32242
rect 22923 -32858 22927 -32242
rect 22623 -32862 22927 -32858
rect 23623 -32242 23927 -32238
rect 23623 -32858 23627 -32242
rect 23627 -32858 23923 -32242
rect 23923 -32858 23927 -32242
rect 23623 -32862 23927 -32858
rect 24623 -32242 24927 -32238
rect 24623 -32858 24627 -32242
rect 24627 -32858 24923 -32242
rect 24923 -32858 24927 -32242
rect 24623 -32862 24927 -32858
rect 25623 -32242 25927 -32238
rect 25623 -32858 25627 -32242
rect 25627 -32858 25923 -32242
rect 25923 -32858 25927 -32242
rect 25623 -32862 25927 -32858
rect 26623 -32242 26927 -32238
rect 26623 -32858 26627 -32242
rect 26627 -32858 26923 -32242
rect 26923 -32858 26927 -32242
rect 26623 -32862 26927 -32858
rect 27623 -32242 27927 -32238
rect 27623 -32858 27627 -32242
rect 27627 -32858 27923 -32242
rect 27923 -32858 27927 -32242
rect 27623 -32862 27927 -32858
rect 28623 -32242 28927 -32238
rect 28623 -32858 28627 -32242
rect 28627 -32858 28923 -32242
rect 28923 -32858 28927 -32242
rect 28623 -32862 28927 -32858
rect 29623 -32242 29927 -32238
rect 29623 -32858 29627 -32242
rect 29627 -32858 29923 -32242
rect 29923 -32858 29927 -32242
rect 29623 -32862 29927 -32858
rect 30623 -32242 30927 -32238
rect 30623 -32858 30627 -32242
rect 30627 -32858 30923 -32242
rect 30923 -32858 30927 -32242
rect 30623 -32862 30927 -32858
rect 31623 -32242 31927 -32238
rect 31623 -32858 31627 -32242
rect 31627 -32858 31923 -32242
rect 31923 -32858 31927 -32242
rect 31623 -32862 31927 -32858
rect 32623 -32242 32927 -32238
rect 32623 -32858 32627 -32242
rect 32627 -32858 32923 -32242
rect 32923 -32858 32927 -32242
rect 32623 -32862 32927 -32858
rect 33623 -32242 33927 -32238
rect 33623 -32858 33627 -32242
rect 33627 -32858 33923 -32242
rect 33923 -32858 33927 -32242
rect 33623 -32862 33927 -32858
rect 8283 -32902 8587 -32898
rect 8283 -33198 8287 -32902
rect 8287 -33198 8583 -32902
rect 8583 -33198 8587 -32902
rect 8283 -33202 8587 -33198
rect 8623 -32902 8927 -32898
rect 8623 -33198 8627 -32902
rect 8627 -33198 8923 -32902
rect 8923 -33198 8927 -32902
rect 8623 -33202 8927 -33198
rect 8963 -32902 9587 -32898
rect 8963 -33198 8967 -32902
rect 8967 -33198 9583 -32902
rect 9583 -33198 9587 -32902
rect 8963 -33202 9587 -33198
rect 9623 -32902 9927 -32898
rect 9623 -33198 9627 -32902
rect 9627 -33198 9923 -32902
rect 9923 -33198 9927 -32902
rect 9623 -33202 9927 -33198
rect 9963 -32902 10587 -32898
rect 9963 -33198 9967 -32902
rect 9967 -33198 10583 -32902
rect 10583 -33198 10587 -32902
rect 9963 -33202 10587 -33198
rect 10623 -32902 10927 -32898
rect 10623 -33198 10627 -32902
rect 10627 -33198 10923 -32902
rect 10923 -33198 10927 -32902
rect 10623 -33202 10927 -33198
rect 10963 -32902 11587 -32898
rect 10963 -33198 10967 -32902
rect 10967 -33198 11583 -32902
rect 11583 -33198 11587 -32902
rect 10963 -33202 11587 -33198
rect 11623 -32902 11927 -32898
rect 11623 -33198 11627 -32902
rect 11627 -33198 11923 -32902
rect 11923 -33198 11927 -32902
rect 11623 -33202 11927 -33198
rect 11963 -32902 12587 -32898
rect 11963 -33198 11967 -32902
rect 11967 -33198 12583 -32902
rect 12583 -33198 12587 -32902
rect 11963 -33202 12587 -33198
rect 12623 -32902 12927 -32898
rect 12623 -33198 12627 -32902
rect 12627 -33198 12923 -32902
rect 12923 -33198 12927 -32902
rect 12623 -33202 12927 -33198
rect 12963 -32902 13587 -32898
rect 12963 -33198 12967 -32902
rect 12967 -33198 13583 -32902
rect 13583 -33198 13587 -32902
rect 12963 -33202 13587 -33198
rect 13623 -32902 13927 -32898
rect 13623 -33198 13627 -32902
rect 13627 -33198 13923 -32902
rect 13923 -33198 13927 -32902
rect 13623 -33202 13927 -33198
rect 13963 -32902 14587 -32898
rect 13963 -33198 13967 -32902
rect 13967 -33198 14583 -32902
rect 14583 -33198 14587 -32902
rect 13963 -33202 14587 -33198
rect 14623 -32902 14927 -32898
rect 14623 -33198 14627 -32902
rect 14627 -33198 14923 -32902
rect 14923 -33198 14927 -32902
rect 14623 -33202 14927 -33198
rect 14963 -32902 15587 -32898
rect 14963 -33198 14967 -32902
rect 14967 -33198 15583 -32902
rect 15583 -33198 15587 -32902
rect 14963 -33202 15587 -33198
rect 15623 -32902 15927 -32898
rect 15623 -33198 15627 -32902
rect 15627 -33198 15923 -32902
rect 15923 -33198 15927 -32902
rect 15623 -33202 15927 -33198
rect 15963 -32902 16587 -32898
rect 15963 -33198 15967 -32902
rect 15967 -33198 16583 -32902
rect 16583 -33198 16587 -32902
rect 15963 -33202 16587 -33198
rect 16623 -32902 16927 -32898
rect 16623 -33198 16627 -32902
rect 16627 -33198 16923 -32902
rect 16923 -33198 16927 -32902
rect 16623 -33202 16927 -33198
rect 16963 -32902 17587 -32898
rect 16963 -33198 16967 -32902
rect 16967 -33198 17583 -32902
rect 17583 -33198 17587 -32902
rect 16963 -33202 17587 -33198
rect 17623 -32902 17927 -32898
rect 17623 -33198 17627 -32902
rect 17627 -33198 17923 -32902
rect 17923 -33198 17927 -32902
rect 17623 -33202 17927 -33198
rect 17963 -32902 18587 -32898
rect 17963 -33198 17967 -32902
rect 17967 -33198 18583 -32902
rect 18583 -33198 18587 -32902
rect 17963 -33202 18587 -33198
rect 18623 -32902 18927 -32898
rect 18623 -33198 18627 -32902
rect 18627 -33198 18923 -32902
rect 18923 -33198 18927 -32902
rect 18623 -33202 18927 -33198
rect 18963 -32902 19587 -32898
rect 18963 -33198 18967 -32902
rect 18967 -33198 19583 -32902
rect 19583 -33198 19587 -32902
rect 18963 -33202 19587 -33198
rect 19623 -32902 19927 -32898
rect 19623 -33198 19627 -32902
rect 19627 -33198 19923 -32902
rect 19923 -33198 19927 -32902
rect 19623 -33202 19927 -33198
rect 19963 -32902 20587 -32898
rect 19963 -33198 19967 -32902
rect 19967 -33198 20583 -32902
rect 20583 -33198 20587 -32902
rect 19963 -33202 20587 -33198
rect 20623 -32902 20927 -32898
rect 20623 -33198 20627 -32902
rect 20627 -33198 20923 -32902
rect 20923 -33198 20927 -32902
rect 20623 -33202 20927 -33198
rect 20963 -32902 21587 -32898
rect 20963 -33198 20967 -32902
rect 20967 -33198 21583 -32902
rect 21583 -33198 21587 -32902
rect 20963 -33202 21587 -33198
rect 21623 -32902 21927 -32898
rect 21623 -33198 21627 -32902
rect 21627 -33198 21923 -32902
rect 21923 -33198 21927 -32902
rect 21623 -33202 21927 -33198
rect 21963 -32902 22587 -32898
rect 21963 -33198 21967 -32902
rect 21967 -33198 22583 -32902
rect 22583 -33198 22587 -32902
rect 21963 -33202 22587 -33198
rect 22623 -32902 22927 -32898
rect 22623 -33198 22627 -32902
rect 22627 -33198 22923 -32902
rect 22923 -33198 22927 -32902
rect 22623 -33202 22927 -33198
rect 22963 -32902 23587 -32898
rect 22963 -33198 22967 -32902
rect 22967 -33198 23583 -32902
rect 23583 -33198 23587 -32902
rect 22963 -33202 23587 -33198
rect 23623 -32902 23927 -32898
rect 23623 -33198 23627 -32902
rect 23627 -33198 23923 -32902
rect 23923 -33198 23927 -32902
rect 23623 -33202 23927 -33198
rect 23963 -32902 24587 -32898
rect 23963 -33198 23967 -32902
rect 23967 -33198 24583 -32902
rect 24583 -33198 24587 -32902
rect 23963 -33202 24587 -33198
rect 24623 -32902 24927 -32898
rect 24623 -33198 24627 -32902
rect 24627 -33198 24923 -32902
rect 24923 -33198 24927 -32902
rect 24623 -33202 24927 -33198
rect 24963 -32902 25587 -32898
rect 24963 -33198 24967 -32902
rect 24967 -33198 25583 -32902
rect 25583 -33198 25587 -32902
rect 24963 -33202 25587 -33198
rect 25623 -32902 25927 -32898
rect 25623 -33198 25627 -32902
rect 25627 -33198 25923 -32902
rect 25923 -33198 25927 -32902
rect 25623 -33202 25927 -33198
rect 25963 -32902 26587 -32898
rect 25963 -33198 25967 -32902
rect 25967 -33198 26583 -32902
rect 26583 -33198 26587 -32902
rect 25963 -33202 26587 -33198
rect 26623 -32902 26927 -32898
rect 26623 -33198 26627 -32902
rect 26627 -33198 26923 -32902
rect 26923 -33198 26927 -32902
rect 26623 -33202 26927 -33198
rect 26963 -32902 27587 -32898
rect 26963 -33198 26967 -32902
rect 26967 -33198 27583 -32902
rect 27583 -33198 27587 -32902
rect 26963 -33202 27587 -33198
rect 27623 -32902 27927 -32898
rect 27623 -33198 27627 -32902
rect 27627 -33198 27923 -32902
rect 27923 -33198 27927 -32902
rect 27623 -33202 27927 -33198
rect 27963 -32902 28587 -32898
rect 27963 -33198 27967 -32902
rect 27967 -33198 28583 -32902
rect 28583 -33198 28587 -32902
rect 27963 -33202 28587 -33198
rect 28623 -32902 28927 -32898
rect 28623 -33198 28627 -32902
rect 28627 -33198 28923 -32902
rect 28923 -33198 28927 -32902
rect 28623 -33202 28927 -33198
rect 28963 -32902 29587 -32898
rect 28963 -33198 28967 -32902
rect 28967 -33198 29583 -32902
rect 29583 -33198 29587 -32902
rect 28963 -33202 29587 -33198
rect 29623 -32902 29927 -32898
rect 29623 -33198 29627 -32902
rect 29627 -33198 29923 -32902
rect 29923 -33198 29927 -32902
rect 29623 -33202 29927 -33198
rect 29963 -32902 30587 -32898
rect 29963 -33198 29967 -32902
rect 29967 -33198 30583 -32902
rect 30583 -33198 30587 -32902
rect 29963 -33202 30587 -33198
rect 30623 -32902 30927 -32898
rect 30623 -33198 30627 -32902
rect 30627 -33198 30923 -32902
rect 30923 -33198 30927 -32902
rect 30623 -33202 30927 -33198
rect 30963 -32902 31587 -32898
rect 30963 -33198 30967 -32902
rect 30967 -33198 31583 -32902
rect 31583 -33198 31587 -32902
rect 30963 -33202 31587 -33198
rect 31623 -32902 31927 -32898
rect 31623 -33198 31627 -32902
rect 31627 -33198 31923 -32902
rect 31923 -33198 31927 -32902
rect 31623 -33202 31927 -33198
rect 31963 -32902 32587 -32898
rect 31963 -33198 31967 -32902
rect 31967 -33198 32583 -32902
rect 32583 -33198 32587 -32902
rect 31963 -33202 32587 -33198
rect 32623 -32902 32927 -32898
rect 32623 -33198 32627 -32902
rect 32627 -33198 32923 -32902
rect 32923 -33198 32927 -32902
rect 32623 -33202 32927 -33198
rect 32963 -32902 33587 -32898
rect 32963 -33198 32967 -32902
rect 32967 -33198 33583 -32902
rect 33583 -33198 33587 -32902
rect 32963 -33202 33587 -33198
rect 33623 -32902 33927 -32898
rect 33623 -33198 33627 -32902
rect 33627 -33198 33923 -32902
rect 33923 -33198 33927 -32902
rect 33623 -33202 33927 -33198
rect 33963 -32902 34267 -32898
rect 33963 -33198 33967 -32902
rect 33967 -33198 34263 -32902
rect 34263 -33198 34267 -32902
rect 33963 -33202 34267 -33198
rect 8623 -33242 8927 -33238
rect 8623 -33858 8627 -33242
rect 8627 -33858 8923 -33242
rect 8923 -33858 8927 -33242
rect 8623 -33862 8927 -33858
rect 9623 -33242 9927 -33238
rect 9623 -33858 9627 -33242
rect 9627 -33858 9923 -33242
rect 9923 -33858 9927 -33242
rect 9623 -33862 9927 -33858
rect 10623 -33242 10927 -33238
rect 10623 -33858 10627 -33242
rect 10627 -33858 10923 -33242
rect 10923 -33858 10927 -33242
rect 10623 -33862 10927 -33858
rect 11623 -33242 11927 -33238
rect 11623 -33858 11627 -33242
rect 11627 -33858 11923 -33242
rect 11923 -33858 11927 -33242
rect 11623 -33862 11927 -33858
rect 12623 -33242 12927 -33238
rect 12623 -33858 12627 -33242
rect 12627 -33858 12923 -33242
rect 12923 -33858 12927 -33242
rect 12623 -33862 12927 -33858
rect 13623 -33242 13927 -33238
rect 13623 -33858 13627 -33242
rect 13627 -33858 13923 -33242
rect 13923 -33858 13927 -33242
rect 13623 -33862 13927 -33858
rect 14623 -33242 14927 -33238
rect 14623 -33858 14627 -33242
rect 14627 -33858 14923 -33242
rect 14923 -33858 14927 -33242
rect 14623 -33862 14927 -33858
rect 15623 -33242 15927 -33238
rect 15623 -33858 15627 -33242
rect 15627 -33858 15923 -33242
rect 15923 -33858 15927 -33242
rect 15623 -33862 15927 -33858
rect 16623 -33242 16927 -33238
rect 16623 -33858 16627 -33242
rect 16627 -33858 16923 -33242
rect 16923 -33858 16927 -33242
rect 16623 -33862 16927 -33858
rect 17623 -33242 17927 -33238
rect 17623 -33858 17627 -33242
rect 17627 -33858 17923 -33242
rect 17923 -33858 17927 -33242
rect 17623 -33862 17927 -33858
rect 18623 -33242 18927 -33238
rect 18623 -33858 18627 -33242
rect 18627 -33858 18923 -33242
rect 18923 -33858 18927 -33242
rect 18623 -33862 18927 -33858
rect 19623 -33242 19927 -33238
rect 19623 -33858 19627 -33242
rect 19627 -33858 19923 -33242
rect 19923 -33858 19927 -33242
rect 19623 -33862 19927 -33858
rect 20623 -33242 20927 -33238
rect 20623 -33858 20627 -33242
rect 20627 -33858 20923 -33242
rect 20923 -33858 20927 -33242
rect 20623 -33862 20927 -33858
rect 21623 -33242 21927 -33238
rect 21623 -33858 21627 -33242
rect 21627 -33858 21923 -33242
rect 21923 -33858 21927 -33242
rect 21623 -33862 21927 -33858
rect 22623 -33242 22927 -33238
rect 22623 -33858 22627 -33242
rect 22627 -33858 22923 -33242
rect 22923 -33858 22927 -33242
rect 22623 -33862 22927 -33858
rect 23623 -33242 23927 -33238
rect 23623 -33858 23627 -33242
rect 23627 -33858 23923 -33242
rect 23923 -33858 23927 -33242
rect 23623 -33862 23927 -33858
rect 24623 -33242 24927 -33238
rect 24623 -33858 24627 -33242
rect 24627 -33858 24923 -33242
rect 24923 -33858 24927 -33242
rect 24623 -33862 24927 -33858
rect 25623 -33242 25927 -33238
rect 25623 -33858 25627 -33242
rect 25627 -33858 25923 -33242
rect 25923 -33858 25927 -33242
rect 25623 -33862 25927 -33858
rect 26623 -33242 26927 -33238
rect 26623 -33858 26627 -33242
rect 26627 -33858 26923 -33242
rect 26923 -33858 26927 -33242
rect 26623 -33862 26927 -33858
rect 27623 -33242 27927 -33238
rect 27623 -33858 27627 -33242
rect 27627 -33858 27923 -33242
rect 27923 -33858 27927 -33242
rect 27623 -33862 27927 -33858
rect 28623 -33242 28927 -33238
rect 28623 -33858 28627 -33242
rect 28627 -33858 28923 -33242
rect 28923 -33858 28927 -33242
rect 28623 -33862 28927 -33858
rect 29623 -33242 29927 -33238
rect 29623 -33858 29627 -33242
rect 29627 -33858 29923 -33242
rect 29923 -33858 29927 -33242
rect 29623 -33862 29927 -33858
rect 30623 -33242 30927 -33238
rect 30623 -33858 30627 -33242
rect 30627 -33858 30923 -33242
rect 30923 -33858 30927 -33242
rect 30623 -33862 30927 -33858
rect 31623 -33242 31927 -33238
rect 31623 -33858 31627 -33242
rect 31627 -33858 31923 -33242
rect 31923 -33858 31927 -33242
rect 31623 -33862 31927 -33858
rect 32623 -33242 32927 -33238
rect 32623 -33858 32627 -33242
rect 32627 -33858 32923 -33242
rect 32923 -33858 32927 -33242
rect 32623 -33862 32927 -33858
rect 33623 -33242 33927 -33238
rect 33623 -33858 33627 -33242
rect 33627 -33858 33923 -33242
rect 33923 -33858 33927 -33242
rect 33623 -33862 33927 -33858
rect 8283 -33902 8587 -33898
rect 8283 -34198 8287 -33902
rect 8287 -34198 8583 -33902
rect 8583 -34198 8587 -33902
rect 8283 -34202 8587 -34198
rect 8623 -33902 8927 -33898
rect 8623 -34198 8627 -33902
rect 8627 -34198 8923 -33902
rect 8923 -34198 8927 -33902
rect 8623 -34202 8927 -34198
rect 8963 -33902 9587 -33898
rect 8963 -34198 8967 -33902
rect 8967 -34198 9583 -33902
rect 9583 -34198 9587 -33902
rect 8963 -34202 9587 -34198
rect 9623 -33902 9927 -33898
rect 9623 -34198 9627 -33902
rect 9627 -34198 9923 -33902
rect 9923 -34198 9927 -33902
rect 9623 -34202 9927 -34198
rect 9963 -33902 10587 -33898
rect 9963 -34198 9967 -33902
rect 9967 -34198 10583 -33902
rect 10583 -34198 10587 -33902
rect 9963 -34202 10587 -34198
rect 10623 -33902 10927 -33898
rect 10623 -34198 10627 -33902
rect 10627 -34198 10923 -33902
rect 10923 -34198 10927 -33902
rect 10623 -34202 10927 -34198
rect 10963 -33902 11587 -33898
rect 10963 -34198 10967 -33902
rect 10967 -34198 11583 -33902
rect 11583 -34198 11587 -33902
rect 10963 -34202 11587 -34198
rect 11623 -33902 11927 -33898
rect 11623 -34198 11627 -33902
rect 11627 -34198 11923 -33902
rect 11923 -34198 11927 -33902
rect 11623 -34202 11927 -34198
rect 11963 -33902 12587 -33898
rect 11963 -34198 11967 -33902
rect 11967 -34198 12583 -33902
rect 12583 -34198 12587 -33902
rect 11963 -34202 12587 -34198
rect 12623 -33902 12927 -33898
rect 12623 -34198 12627 -33902
rect 12627 -34198 12923 -33902
rect 12923 -34198 12927 -33902
rect 12623 -34202 12927 -34198
rect 12963 -33902 13587 -33898
rect 12963 -34198 12967 -33902
rect 12967 -34198 13583 -33902
rect 13583 -34198 13587 -33902
rect 12963 -34202 13587 -34198
rect 13623 -33902 13927 -33898
rect 13623 -34198 13627 -33902
rect 13627 -34198 13923 -33902
rect 13923 -34198 13927 -33902
rect 13623 -34202 13927 -34198
rect 13963 -33902 14587 -33898
rect 13963 -34198 13967 -33902
rect 13967 -34198 14583 -33902
rect 14583 -34198 14587 -33902
rect 13963 -34202 14587 -34198
rect 14623 -33902 14927 -33898
rect 14623 -34198 14627 -33902
rect 14627 -34198 14923 -33902
rect 14923 -34198 14927 -33902
rect 14623 -34202 14927 -34198
rect 14963 -33902 15587 -33898
rect 14963 -34198 14967 -33902
rect 14967 -34198 15583 -33902
rect 15583 -34198 15587 -33902
rect 14963 -34202 15587 -34198
rect 15623 -33902 15927 -33898
rect 15623 -34198 15627 -33902
rect 15627 -34198 15923 -33902
rect 15923 -34198 15927 -33902
rect 15623 -34202 15927 -34198
rect 15963 -33902 16587 -33898
rect 15963 -34198 15967 -33902
rect 15967 -34198 16583 -33902
rect 16583 -34198 16587 -33902
rect 15963 -34202 16587 -34198
rect 16623 -33902 16927 -33898
rect 16623 -34198 16627 -33902
rect 16627 -34198 16923 -33902
rect 16923 -34198 16927 -33902
rect 16623 -34202 16927 -34198
rect 16963 -33902 17587 -33898
rect 16963 -34198 16967 -33902
rect 16967 -34198 17583 -33902
rect 17583 -34198 17587 -33902
rect 16963 -34202 17587 -34198
rect 17623 -33902 17927 -33898
rect 17623 -34198 17627 -33902
rect 17627 -34198 17923 -33902
rect 17923 -34198 17927 -33902
rect 17623 -34202 17927 -34198
rect 17963 -33902 18587 -33898
rect 17963 -34198 17967 -33902
rect 17967 -34198 18583 -33902
rect 18583 -34198 18587 -33902
rect 17963 -34202 18587 -34198
rect 18623 -33902 18927 -33898
rect 18623 -34198 18627 -33902
rect 18627 -34198 18923 -33902
rect 18923 -34198 18927 -33902
rect 18623 -34202 18927 -34198
rect 18963 -33902 19587 -33898
rect 18963 -34198 18967 -33902
rect 18967 -34198 19583 -33902
rect 19583 -34198 19587 -33902
rect 18963 -34202 19587 -34198
rect 19623 -33902 19927 -33898
rect 19623 -34198 19627 -33902
rect 19627 -34198 19923 -33902
rect 19923 -34198 19927 -33902
rect 19623 -34202 19927 -34198
rect 19963 -33902 20587 -33898
rect 19963 -34198 19967 -33902
rect 19967 -34198 20583 -33902
rect 20583 -34198 20587 -33902
rect 19963 -34202 20587 -34198
rect 20623 -33902 20927 -33898
rect 20623 -34198 20627 -33902
rect 20627 -34198 20923 -33902
rect 20923 -34198 20927 -33902
rect 20623 -34202 20927 -34198
rect 20963 -33902 21587 -33898
rect 20963 -34198 20967 -33902
rect 20967 -34198 21583 -33902
rect 21583 -34198 21587 -33902
rect 20963 -34202 21587 -34198
rect 21623 -33902 21927 -33898
rect 21623 -34198 21627 -33902
rect 21627 -34198 21923 -33902
rect 21923 -34198 21927 -33902
rect 21623 -34202 21927 -34198
rect 21963 -33902 22587 -33898
rect 21963 -34198 21967 -33902
rect 21967 -34198 22583 -33902
rect 22583 -34198 22587 -33902
rect 21963 -34202 22587 -34198
rect 22623 -33902 22927 -33898
rect 22623 -34198 22627 -33902
rect 22627 -34198 22923 -33902
rect 22923 -34198 22927 -33902
rect 22623 -34202 22927 -34198
rect 22963 -33902 23587 -33898
rect 22963 -34198 22967 -33902
rect 22967 -34198 23583 -33902
rect 23583 -34198 23587 -33902
rect 22963 -34202 23587 -34198
rect 23623 -33902 23927 -33898
rect 23623 -34198 23627 -33902
rect 23627 -34198 23923 -33902
rect 23923 -34198 23927 -33902
rect 23623 -34202 23927 -34198
rect 23963 -33902 24587 -33898
rect 23963 -34198 23967 -33902
rect 23967 -34198 24583 -33902
rect 24583 -34198 24587 -33902
rect 23963 -34202 24587 -34198
rect 24623 -33902 24927 -33898
rect 24623 -34198 24627 -33902
rect 24627 -34198 24923 -33902
rect 24923 -34198 24927 -33902
rect 24623 -34202 24927 -34198
rect 24963 -33902 25587 -33898
rect 24963 -34198 24967 -33902
rect 24967 -34198 25583 -33902
rect 25583 -34198 25587 -33902
rect 24963 -34202 25587 -34198
rect 25623 -33902 25927 -33898
rect 25623 -34198 25627 -33902
rect 25627 -34198 25923 -33902
rect 25923 -34198 25927 -33902
rect 25623 -34202 25927 -34198
rect 25963 -33902 26587 -33898
rect 25963 -34198 25967 -33902
rect 25967 -34198 26583 -33902
rect 26583 -34198 26587 -33902
rect 25963 -34202 26587 -34198
rect 26623 -33902 26927 -33898
rect 26623 -34198 26627 -33902
rect 26627 -34198 26923 -33902
rect 26923 -34198 26927 -33902
rect 26623 -34202 26927 -34198
rect 26963 -33902 27587 -33898
rect 26963 -34198 26967 -33902
rect 26967 -34198 27583 -33902
rect 27583 -34198 27587 -33902
rect 26963 -34202 27587 -34198
rect 27623 -33902 27927 -33898
rect 27623 -34198 27627 -33902
rect 27627 -34198 27923 -33902
rect 27923 -34198 27927 -33902
rect 27623 -34202 27927 -34198
rect 27963 -33902 28587 -33898
rect 27963 -34198 27967 -33902
rect 27967 -34198 28583 -33902
rect 28583 -34198 28587 -33902
rect 27963 -34202 28587 -34198
rect 28623 -33902 28927 -33898
rect 28623 -34198 28627 -33902
rect 28627 -34198 28923 -33902
rect 28923 -34198 28927 -33902
rect 28623 -34202 28927 -34198
rect 28963 -33902 29587 -33898
rect 28963 -34198 28967 -33902
rect 28967 -34198 29583 -33902
rect 29583 -34198 29587 -33902
rect 28963 -34202 29587 -34198
rect 29623 -33902 29927 -33898
rect 29623 -34198 29627 -33902
rect 29627 -34198 29923 -33902
rect 29923 -34198 29927 -33902
rect 29623 -34202 29927 -34198
rect 29963 -33902 30587 -33898
rect 29963 -34198 29967 -33902
rect 29967 -34198 30583 -33902
rect 30583 -34198 30587 -33902
rect 29963 -34202 30587 -34198
rect 30623 -33902 30927 -33898
rect 30623 -34198 30627 -33902
rect 30627 -34198 30923 -33902
rect 30923 -34198 30927 -33902
rect 30623 -34202 30927 -34198
rect 30963 -33902 31587 -33898
rect 30963 -34198 30967 -33902
rect 30967 -34198 31583 -33902
rect 31583 -34198 31587 -33902
rect 30963 -34202 31587 -34198
rect 31623 -33902 31927 -33898
rect 31623 -34198 31627 -33902
rect 31627 -34198 31923 -33902
rect 31923 -34198 31927 -33902
rect 31623 -34202 31927 -34198
rect 31963 -33902 32587 -33898
rect 31963 -34198 31967 -33902
rect 31967 -34198 32583 -33902
rect 32583 -34198 32587 -33902
rect 31963 -34202 32587 -34198
rect 32623 -33902 32927 -33898
rect 32623 -34198 32627 -33902
rect 32627 -34198 32923 -33902
rect 32923 -34198 32927 -33902
rect 32623 -34202 32927 -34198
rect 32963 -33902 33587 -33898
rect 32963 -34198 32967 -33902
rect 32967 -34198 33583 -33902
rect 33583 -34198 33587 -33902
rect 32963 -34202 33587 -34198
rect 33623 -33902 33927 -33898
rect 33623 -34198 33627 -33902
rect 33627 -34198 33923 -33902
rect 33923 -34198 33927 -33902
rect 33623 -34202 33927 -34198
rect 33963 -33902 34267 -33898
rect 33963 -34198 33967 -33902
rect 33967 -34198 34263 -33902
rect 34263 -34198 34267 -33902
rect 33963 -34202 34267 -34198
rect 8623 -34242 8927 -34238
rect 8623 -34858 8627 -34242
rect 8627 -34858 8923 -34242
rect 8923 -34858 8927 -34242
rect 8623 -34862 8927 -34858
rect 9623 -34242 9927 -34238
rect 9623 -34858 9627 -34242
rect 9627 -34858 9923 -34242
rect 9923 -34858 9927 -34242
rect 9623 -34862 9927 -34858
rect 10623 -34242 10927 -34238
rect 10623 -34858 10627 -34242
rect 10627 -34858 10923 -34242
rect 10923 -34858 10927 -34242
rect 10623 -34862 10927 -34858
rect 11623 -34242 11927 -34238
rect 11623 -34858 11627 -34242
rect 11627 -34858 11923 -34242
rect 11923 -34858 11927 -34242
rect 11623 -34862 11927 -34858
rect 12623 -34242 12927 -34238
rect 12623 -34858 12627 -34242
rect 12627 -34858 12923 -34242
rect 12923 -34858 12927 -34242
rect 12623 -34862 12927 -34858
rect 13623 -34242 13927 -34238
rect 13623 -34858 13627 -34242
rect 13627 -34858 13923 -34242
rect 13923 -34858 13927 -34242
rect 13623 -34862 13927 -34858
rect 14623 -34242 14927 -34238
rect 14623 -34858 14627 -34242
rect 14627 -34858 14923 -34242
rect 14923 -34858 14927 -34242
rect 14623 -34862 14927 -34858
rect 15623 -34242 15927 -34238
rect 15623 -34858 15627 -34242
rect 15627 -34858 15923 -34242
rect 15923 -34858 15927 -34242
rect 15623 -34862 15927 -34858
rect 16623 -34242 16927 -34238
rect 16623 -34858 16627 -34242
rect 16627 -34858 16923 -34242
rect 16923 -34858 16927 -34242
rect 16623 -34862 16927 -34858
rect 17623 -34242 17927 -34238
rect 17623 -34858 17627 -34242
rect 17627 -34858 17923 -34242
rect 17923 -34858 17927 -34242
rect 17623 -34862 17927 -34858
rect 18623 -34242 18927 -34238
rect 18623 -34858 18627 -34242
rect 18627 -34858 18923 -34242
rect 18923 -34858 18927 -34242
rect 18623 -34862 18927 -34858
rect 19623 -34242 19927 -34238
rect 19623 -34858 19627 -34242
rect 19627 -34858 19923 -34242
rect 19923 -34858 19927 -34242
rect 19623 -34862 19927 -34858
rect 20623 -34242 20927 -34238
rect 20623 -34858 20627 -34242
rect 20627 -34858 20923 -34242
rect 20923 -34858 20927 -34242
rect 20623 -34862 20927 -34858
rect 21623 -34242 21927 -34238
rect 21623 -34858 21627 -34242
rect 21627 -34858 21923 -34242
rect 21923 -34858 21927 -34242
rect 21623 -34862 21927 -34858
rect 22623 -34242 22927 -34238
rect 22623 -34858 22627 -34242
rect 22627 -34858 22923 -34242
rect 22923 -34858 22927 -34242
rect 22623 -34862 22927 -34858
rect 23623 -34242 23927 -34238
rect 23623 -34858 23627 -34242
rect 23627 -34858 23923 -34242
rect 23923 -34858 23927 -34242
rect 23623 -34862 23927 -34858
rect 24623 -34242 24927 -34238
rect 24623 -34858 24627 -34242
rect 24627 -34858 24923 -34242
rect 24923 -34858 24927 -34242
rect 24623 -34862 24927 -34858
rect 25623 -34242 25927 -34238
rect 25623 -34858 25627 -34242
rect 25627 -34858 25923 -34242
rect 25923 -34858 25927 -34242
rect 25623 -34862 25927 -34858
rect 26623 -34242 26927 -34238
rect 26623 -34858 26627 -34242
rect 26627 -34858 26923 -34242
rect 26923 -34858 26927 -34242
rect 26623 -34862 26927 -34858
rect 27623 -34242 27927 -34238
rect 27623 -34858 27627 -34242
rect 27627 -34858 27923 -34242
rect 27923 -34858 27927 -34242
rect 27623 -34862 27927 -34858
rect 28623 -34242 28927 -34238
rect 28623 -34858 28627 -34242
rect 28627 -34858 28923 -34242
rect 28923 -34858 28927 -34242
rect 28623 -34862 28927 -34858
rect 29623 -34242 29927 -34238
rect 29623 -34858 29627 -34242
rect 29627 -34858 29923 -34242
rect 29923 -34858 29927 -34242
rect 29623 -34862 29927 -34858
rect 30623 -34242 30927 -34238
rect 30623 -34858 30627 -34242
rect 30627 -34858 30923 -34242
rect 30923 -34858 30927 -34242
rect 30623 -34862 30927 -34858
rect 31623 -34242 31927 -34238
rect 31623 -34858 31627 -34242
rect 31627 -34858 31923 -34242
rect 31923 -34858 31927 -34242
rect 31623 -34862 31927 -34858
rect 32623 -34242 32927 -34238
rect 32623 -34858 32627 -34242
rect 32627 -34858 32923 -34242
rect 32923 -34858 32927 -34242
rect 32623 -34862 32927 -34858
rect 33623 -34242 33927 -34238
rect 33623 -34858 33627 -34242
rect 33627 -34858 33923 -34242
rect 33923 -34858 33927 -34242
rect 33623 -34862 33927 -34858
rect 8283 -34902 8587 -34898
rect 8283 -35198 8287 -34902
rect 8287 -35198 8583 -34902
rect 8583 -35198 8587 -34902
rect 8283 -35202 8587 -35198
rect 8623 -34902 8927 -34898
rect 8623 -35198 8627 -34902
rect 8627 -35198 8923 -34902
rect 8923 -35198 8927 -34902
rect 8623 -35202 8927 -35198
rect 8963 -34902 9587 -34898
rect 8963 -35198 8967 -34902
rect 8967 -35198 9583 -34902
rect 9583 -35198 9587 -34902
rect 8963 -35202 9587 -35198
rect 9623 -34902 9927 -34898
rect 9623 -35198 9627 -34902
rect 9627 -35198 9923 -34902
rect 9923 -35198 9927 -34902
rect 9623 -35202 9927 -35198
rect 9963 -34902 10587 -34898
rect 9963 -35198 9967 -34902
rect 9967 -35198 10583 -34902
rect 10583 -35198 10587 -34902
rect 9963 -35202 10587 -35198
rect 10623 -34902 10927 -34898
rect 10623 -35198 10627 -34902
rect 10627 -35198 10923 -34902
rect 10923 -35198 10927 -34902
rect 10623 -35202 10927 -35198
rect 10963 -34902 11587 -34898
rect 10963 -35198 10967 -34902
rect 10967 -35198 11583 -34902
rect 11583 -35198 11587 -34902
rect 10963 -35202 11587 -35198
rect 11623 -34902 11927 -34898
rect 11623 -35198 11627 -34902
rect 11627 -35198 11923 -34902
rect 11923 -35198 11927 -34902
rect 11623 -35202 11927 -35198
rect 11963 -34902 12587 -34898
rect 11963 -35198 11967 -34902
rect 11967 -35198 12583 -34902
rect 12583 -35198 12587 -34902
rect 11963 -35202 12587 -35198
rect 12623 -34902 12927 -34898
rect 12623 -35198 12627 -34902
rect 12627 -35198 12923 -34902
rect 12923 -35198 12927 -34902
rect 12623 -35202 12927 -35198
rect 12963 -34902 13587 -34898
rect 12963 -35198 12967 -34902
rect 12967 -35198 13583 -34902
rect 13583 -35198 13587 -34902
rect 12963 -35202 13587 -35198
rect 13623 -34902 13927 -34898
rect 13623 -35198 13627 -34902
rect 13627 -35198 13923 -34902
rect 13923 -35198 13927 -34902
rect 13623 -35202 13927 -35198
rect 13963 -34902 14587 -34898
rect 13963 -35198 13967 -34902
rect 13967 -35198 14583 -34902
rect 14583 -35198 14587 -34902
rect 13963 -35202 14587 -35198
rect 14623 -34902 14927 -34898
rect 14623 -35198 14627 -34902
rect 14627 -35198 14923 -34902
rect 14923 -35198 14927 -34902
rect 14623 -35202 14927 -35198
rect 14963 -34902 15587 -34898
rect 14963 -35198 14967 -34902
rect 14967 -35198 15583 -34902
rect 15583 -35198 15587 -34902
rect 14963 -35202 15587 -35198
rect 15623 -34902 15927 -34898
rect 15623 -35198 15627 -34902
rect 15627 -35198 15923 -34902
rect 15923 -35198 15927 -34902
rect 15623 -35202 15927 -35198
rect 15963 -34902 16587 -34898
rect 15963 -35198 15967 -34902
rect 15967 -35198 16583 -34902
rect 16583 -35198 16587 -34902
rect 15963 -35202 16587 -35198
rect 16623 -34902 16927 -34898
rect 16623 -35198 16627 -34902
rect 16627 -35198 16923 -34902
rect 16923 -35198 16927 -34902
rect 16623 -35202 16927 -35198
rect 16963 -34902 17587 -34898
rect 16963 -35198 16967 -34902
rect 16967 -35198 17583 -34902
rect 17583 -35198 17587 -34902
rect 16963 -35202 17587 -35198
rect 17623 -34902 17927 -34898
rect 17623 -35198 17627 -34902
rect 17627 -35198 17923 -34902
rect 17923 -35198 17927 -34902
rect 17623 -35202 17927 -35198
rect 17963 -34902 18587 -34898
rect 17963 -35198 17967 -34902
rect 17967 -35198 18583 -34902
rect 18583 -35198 18587 -34902
rect 17963 -35202 18587 -35198
rect 18623 -34902 18927 -34898
rect 18623 -35198 18627 -34902
rect 18627 -35198 18923 -34902
rect 18923 -35198 18927 -34902
rect 18623 -35202 18927 -35198
rect 18963 -34902 19587 -34898
rect 18963 -35198 18967 -34902
rect 18967 -35198 19583 -34902
rect 19583 -35198 19587 -34902
rect 18963 -35202 19587 -35198
rect 19623 -34902 19927 -34898
rect 19623 -35198 19627 -34902
rect 19627 -35198 19923 -34902
rect 19923 -35198 19927 -34902
rect 19623 -35202 19927 -35198
rect 19963 -34902 20587 -34898
rect 19963 -35198 19967 -34902
rect 19967 -35198 20583 -34902
rect 20583 -35198 20587 -34902
rect 19963 -35202 20587 -35198
rect 20623 -34902 20927 -34898
rect 20623 -35198 20627 -34902
rect 20627 -35198 20923 -34902
rect 20923 -35198 20927 -34902
rect 20623 -35202 20927 -35198
rect 20963 -34902 21587 -34898
rect 20963 -35198 20967 -34902
rect 20967 -35198 21583 -34902
rect 21583 -35198 21587 -34902
rect 20963 -35202 21587 -35198
rect 21623 -34902 21927 -34898
rect 21623 -35198 21627 -34902
rect 21627 -35198 21923 -34902
rect 21923 -35198 21927 -34902
rect 21623 -35202 21927 -35198
rect 21963 -34902 22587 -34898
rect 21963 -35198 21967 -34902
rect 21967 -35198 22583 -34902
rect 22583 -35198 22587 -34902
rect 21963 -35202 22587 -35198
rect 22623 -34902 22927 -34898
rect 22623 -35198 22627 -34902
rect 22627 -35198 22923 -34902
rect 22923 -35198 22927 -34902
rect 22623 -35202 22927 -35198
rect 22963 -34902 23587 -34898
rect 22963 -35198 22967 -34902
rect 22967 -35198 23583 -34902
rect 23583 -35198 23587 -34902
rect 22963 -35202 23587 -35198
rect 23623 -34902 23927 -34898
rect 23623 -35198 23627 -34902
rect 23627 -35198 23923 -34902
rect 23923 -35198 23927 -34902
rect 23623 -35202 23927 -35198
rect 23963 -34902 24587 -34898
rect 23963 -35198 23967 -34902
rect 23967 -35198 24583 -34902
rect 24583 -35198 24587 -34902
rect 23963 -35202 24587 -35198
rect 24623 -34902 24927 -34898
rect 24623 -35198 24627 -34902
rect 24627 -35198 24923 -34902
rect 24923 -35198 24927 -34902
rect 24623 -35202 24927 -35198
rect 24963 -34902 25587 -34898
rect 24963 -35198 24967 -34902
rect 24967 -35198 25583 -34902
rect 25583 -35198 25587 -34902
rect 24963 -35202 25587 -35198
rect 25623 -34902 25927 -34898
rect 25623 -35198 25627 -34902
rect 25627 -35198 25923 -34902
rect 25923 -35198 25927 -34902
rect 25623 -35202 25927 -35198
rect 25963 -34902 26587 -34898
rect 25963 -35198 25967 -34902
rect 25967 -35198 26583 -34902
rect 26583 -35198 26587 -34902
rect 25963 -35202 26587 -35198
rect 26623 -34902 26927 -34898
rect 26623 -35198 26627 -34902
rect 26627 -35198 26923 -34902
rect 26923 -35198 26927 -34902
rect 26623 -35202 26927 -35198
rect 26963 -34902 27587 -34898
rect 26963 -35198 26967 -34902
rect 26967 -35198 27583 -34902
rect 27583 -35198 27587 -34902
rect 26963 -35202 27587 -35198
rect 27623 -34902 27927 -34898
rect 27623 -35198 27627 -34902
rect 27627 -35198 27923 -34902
rect 27923 -35198 27927 -34902
rect 27623 -35202 27927 -35198
rect 27963 -34902 28587 -34898
rect 27963 -35198 27967 -34902
rect 27967 -35198 28583 -34902
rect 28583 -35198 28587 -34902
rect 27963 -35202 28587 -35198
rect 28623 -34902 28927 -34898
rect 28623 -35198 28627 -34902
rect 28627 -35198 28923 -34902
rect 28923 -35198 28927 -34902
rect 28623 -35202 28927 -35198
rect 28963 -34902 29587 -34898
rect 28963 -35198 28967 -34902
rect 28967 -35198 29583 -34902
rect 29583 -35198 29587 -34902
rect 28963 -35202 29587 -35198
rect 29623 -34902 29927 -34898
rect 29623 -35198 29627 -34902
rect 29627 -35198 29923 -34902
rect 29923 -35198 29927 -34902
rect 29623 -35202 29927 -35198
rect 29963 -34902 30587 -34898
rect 29963 -35198 29967 -34902
rect 29967 -35198 30583 -34902
rect 30583 -35198 30587 -34902
rect 29963 -35202 30587 -35198
rect 30623 -34902 30927 -34898
rect 30623 -35198 30627 -34902
rect 30627 -35198 30923 -34902
rect 30923 -35198 30927 -34902
rect 30623 -35202 30927 -35198
rect 30963 -34902 31587 -34898
rect 30963 -35198 30967 -34902
rect 30967 -35198 31583 -34902
rect 31583 -35198 31587 -34902
rect 30963 -35202 31587 -35198
rect 31623 -34902 31927 -34898
rect 31623 -35198 31627 -34902
rect 31627 -35198 31923 -34902
rect 31923 -35198 31927 -34902
rect 31623 -35202 31927 -35198
rect 31963 -34902 32587 -34898
rect 31963 -35198 31967 -34902
rect 31967 -35198 32583 -34902
rect 32583 -35198 32587 -34902
rect 31963 -35202 32587 -35198
rect 32623 -34902 32927 -34898
rect 32623 -35198 32627 -34902
rect 32627 -35198 32923 -34902
rect 32923 -35198 32927 -34902
rect 32623 -35202 32927 -35198
rect 32963 -34902 33587 -34898
rect 32963 -35198 32967 -34902
rect 32967 -35198 33583 -34902
rect 33583 -35198 33587 -34902
rect 32963 -35202 33587 -35198
rect 33623 -34902 33927 -34898
rect 33623 -35198 33627 -34902
rect 33627 -35198 33923 -34902
rect 33923 -35198 33927 -34902
rect 33623 -35202 33927 -35198
rect 33963 -34902 34267 -34898
rect 33963 -35198 33967 -34902
rect 33967 -35198 34263 -34902
rect 34263 -35198 34267 -34902
rect 33963 -35202 34267 -35198
rect 8623 -35242 8927 -35238
rect 8623 -35858 8627 -35242
rect 8627 -35858 8923 -35242
rect 8923 -35858 8927 -35242
rect 8623 -35862 8927 -35858
rect 9623 -35242 9927 -35238
rect 9623 -35858 9627 -35242
rect 9627 -35858 9923 -35242
rect 9923 -35858 9927 -35242
rect 9623 -35862 9927 -35858
rect 10623 -35242 10927 -35238
rect 10623 -35858 10627 -35242
rect 10627 -35858 10923 -35242
rect 10923 -35858 10927 -35242
rect 10623 -35862 10927 -35858
rect 11623 -35242 11927 -35238
rect 11623 -35858 11627 -35242
rect 11627 -35858 11923 -35242
rect 11923 -35858 11927 -35242
rect 11623 -35862 11927 -35858
rect 12623 -35242 12927 -35238
rect 12623 -35858 12627 -35242
rect 12627 -35858 12923 -35242
rect 12923 -35858 12927 -35242
rect 12623 -35862 12927 -35858
rect 13623 -35242 13927 -35238
rect 13623 -35858 13627 -35242
rect 13627 -35858 13923 -35242
rect 13923 -35858 13927 -35242
rect 13623 -35862 13927 -35858
rect 14623 -35242 14927 -35238
rect 14623 -35858 14627 -35242
rect 14627 -35858 14923 -35242
rect 14923 -35858 14927 -35242
rect 14623 -35862 14927 -35858
rect 15623 -35242 15927 -35238
rect 15623 -35858 15627 -35242
rect 15627 -35858 15923 -35242
rect 15923 -35858 15927 -35242
rect 15623 -35862 15927 -35858
rect 16623 -35242 16927 -35238
rect 16623 -35858 16627 -35242
rect 16627 -35858 16923 -35242
rect 16923 -35858 16927 -35242
rect 16623 -35862 16927 -35858
rect 17623 -35242 17927 -35238
rect 17623 -35858 17627 -35242
rect 17627 -35858 17923 -35242
rect 17923 -35858 17927 -35242
rect 17623 -35862 17927 -35858
rect 18623 -35242 18927 -35238
rect 18623 -35858 18627 -35242
rect 18627 -35858 18923 -35242
rect 18923 -35858 18927 -35242
rect 18623 -35862 18927 -35858
rect 19623 -35242 19927 -35238
rect 19623 -35858 19627 -35242
rect 19627 -35858 19923 -35242
rect 19923 -35858 19927 -35242
rect 19623 -35862 19927 -35858
rect 20623 -35242 20927 -35238
rect 20623 -35858 20627 -35242
rect 20627 -35858 20923 -35242
rect 20923 -35858 20927 -35242
rect 20623 -35862 20927 -35858
rect 21623 -35242 21927 -35238
rect 21623 -35858 21627 -35242
rect 21627 -35858 21923 -35242
rect 21923 -35858 21927 -35242
rect 21623 -35862 21927 -35858
rect 22623 -35242 22927 -35238
rect 22623 -35858 22627 -35242
rect 22627 -35858 22923 -35242
rect 22923 -35858 22927 -35242
rect 22623 -35862 22927 -35858
rect 23623 -35242 23927 -35238
rect 23623 -35858 23627 -35242
rect 23627 -35858 23923 -35242
rect 23923 -35858 23927 -35242
rect 23623 -35862 23927 -35858
rect 24623 -35242 24927 -35238
rect 24623 -35858 24627 -35242
rect 24627 -35858 24923 -35242
rect 24923 -35858 24927 -35242
rect 24623 -35862 24927 -35858
rect 25623 -35242 25927 -35238
rect 25623 -35858 25627 -35242
rect 25627 -35858 25923 -35242
rect 25923 -35858 25927 -35242
rect 25623 -35862 25927 -35858
rect 26623 -35242 26927 -35238
rect 26623 -35858 26627 -35242
rect 26627 -35858 26923 -35242
rect 26923 -35858 26927 -35242
rect 26623 -35862 26927 -35858
rect 27623 -35242 27927 -35238
rect 27623 -35858 27627 -35242
rect 27627 -35858 27923 -35242
rect 27923 -35858 27927 -35242
rect 27623 -35862 27927 -35858
rect 28623 -35242 28927 -35238
rect 28623 -35858 28627 -35242
rect 28627 -35858 28923 -35242
rect 28923 -35858 28927 -35242
rect 28623 -35862 28927 -35858
rect 29623 -35242 29927 -35238
rect 29623 -35858 29627 -35242
rect 29627 -35858 29923 -35242
rect 29923 -35858 29927 -35242
rect 29623 -35862 29927 -35858
rect 30623 -35242 30927 -35238
rect 30623 -35858 30627 -35242
rect 30627 -35858 30923 -35242
rect 30923 -35858 30927 -35242
rect 30623 -35862 30927 -35858
rect 31623 -35242 31927 -35238
rect 31623 -35858 31627 -35242
rect 31627 -35858 31923 -35242
rect 31923 -35858 31927 -35242
rect 31623 -35862 31927 -35858
rect 32623 -35242 32927 -35238
rect 32623 -35858 32627 -35242
rect 32627 -35858 32923 -35242
rect 32923 -35858 32927 -35242
rect 32623 -35862 32927 -35858
rect 33623 -35242 33927 -35238
rect 33623 -35858 33627 -35242
rect 33627 -35858 33923 -35242
rect 33923 -35858 33927 -35242
rect 33623 -35862 33927 -35858
rect 8283 -35902 8587 -35898
rect 8283 -36198 8287 -35902
rect 8287 -36198 8583 -35902
rect 8583 -36198 8587 -35902
rect 8283 -36202 8587 -36198
rect 8623 -35902 8927 -35898
rect 8623 -36198 8627 -35902
rect 8627 -36198 8923 -35902
rect 8923 -36198 8927 -35902
rect 8623 -36202 8927 -36198
rect 8963 -35902 9587 -35898
rect 8963 -36198 8967 -35902
rect 8967 -36198 9583 -35902
rect 9583 -36198 9587 -35902
rect 8963 -36202 9587 -36198
rect 9623 -35902 9927 -35898
rect 9623 -36198 9627 -35902
rect 9627 -36198 9923 -35902
rect 9923 -36198 9927 -35902
rect 9623 -36202 9927 -36198
rect 9963 -35902 10587 -35898
rect 9963 -36198 9967 -35902
rect 9967 -36198 10583 -35902
rect 10583 -36198 10587 -35902
rect 9963 -36202 10587 -36198
rect 10623 -35902 10927 -35898
rect 10623 -36198 10627 -35902
rect 10627 -36198 10923 -35902
rect 10923 -36198 10927 -35902
rect 10623 -36202 10927 -36198
rect 10963 -35902 11587 -35898
rect 10963 -36198 10967 -35902
rect 10967 -36198 11583 -35902
rect 11583 -36198 11587 -35902
rect 10963 -36202 11587 -36198
rect 11623 -35902 11927 -35898
rect 11623 -36198 11627 -35902
rect 11627 -36198 11923 -35902
rect 11923 -36198 11927 -35902
rect 11623 -36202 11927 -36198
rect 11963 -35902 12587 -35898
rect 11963 -36198 11967 -35902
rect 11967 -36198 12583 -35902
rect 12583 -36198 12587 -35902
rect 11963 -36202 12587 -36198
rect 12623 -35902 12927 -35898
rect 12623 -36198 12627 -35902
rect 12627 -36198 12923 -35902
rect 12923 -36198 12927 -35902
rect 12623 -36202 12927 -36198
rect 12963 -35902 13587 -35898
rect 12963 -36198 12967 -35902
rect 12967 -36198 13583 -35902
rect 13583 -36198 13587 -35902
rect 12963 -36202 13587 -36198
rect 13623 -35902 13927 -35898
rect 13623 -36198 13627 -35902
rect 13627 -36198 13923 -35902
rect 13923 -36198 13927 -35902
rect 13623 -36202 13927 -36198
rect 13963 -35902 14587 -35898
rect 13963 -36198 13967 -35902
rect 13967 -36198 14583 -35902
rect 14583 -36198 14587 -35902
rect 13963 -36202 14587 -36198
rect 14623 -35902 14927 -35898
rect 14623 -36198 14627 -35902
rect 14627 -36198 14923 -35902
rect 14923 -36198 14927 -35902
rect 14623 -36202 14927 -36198
rect 14963 -35902 15587 -35898
rect 14963 -36198 14967 -35902
rect 14967 -36198 15583 -35902
rect 15583 -36198 15587 -35902
rect 14963 -36202 15587 -36198
rect 15623 -35902 15927 -35898
rect 15623 -36198 15627 -35902
rect 15627 -36198 15923 -35902
rect 15923 -36198 15927 -35902
rect 15623 -36202 15927 -36198
rect 15963 -35902 16587 -35898
rect 15963 -36198 15967 -35902
rect 15967 -36198 16583 -35902
rect 16583 -36198 16587 -35902
rect 15963 -36202 16587 -36198
rect 16623 -35902 16927 -35898
rect 16623 -36198 16627 -35902
rect 16627 -36198 16923 -35902
rect 16923 -36198 16927 -35902
rect 16623 -36202 16927 -36198
rect 16963 -35902 17587 -35898
rect 16963 -36198 16967 -35902
rect 16967 -36198 17583 -35902
rect 17583 -36198 17587 -35902
rect 16963 -36202 17587 -36198
rect 17623 -35902 17927 -35898
rect 17623 -36198 17627 -35902
rect 17627 -36198 17923 -35902
rect 17923 -36198 17927 -35902
rect 17623 -36202 17927 -36198
rect 17963 -35902 18587 -35898
rect 17963 -36198 17967 -35902
rect 17967 -36198 18583 -35902
rect 18583 -36198 18587 -35902
rect 17963 -36202 18587 -36198
rect 18623 -35902 18927 -35898
rect 18623 -36198 18627 -35902
rect 18627 -36198 18923 -35902
rect 18923 -36198 18927 -35902
rect 18623 -36202 18927 -36198
rect 18963 -35902 19587 -35898
rect 18963 -36198 18967 -35902
rect 18967 -36198 19583 -35902
rect 19583 -36198 19587 -35902
rect 18963 -36202 19587 -36198
rect 19623 -35902 19927 -35898
rect 19623 -36198 19627 -35902
rect 19627 -36198 19923 -35902
rect 19923 -36198 19927 -35902
rect 19623 -36202 19927 -36198
rect 19963 -35902 20587 -35898
rect 19963 -36198 19967 -35902
rect 19967 -36198 20583 -35902
rect 20583 -36198 20587 -35902
rect 19963 -36202 20587 -36198
rect 20623 -35902 20927 -35898
rect 20623 -36198 20627 -35902
rect 20627 -36198 20923 -35902
rect 20923 -36198 20927 -35902
rect 20623 -36202 20927 -36198
rect 20963 -35902 21587 -35898
rect 20963 -36198 20967 -35902
rect 20967 -36198 21583 -35902
rect 21583 -36198 21587 -35902
rect 20963 -36202 21587 -36198
rect 21623 -35902 21927 -35898
rect 21623 -36198 21627 -35902
rect 21627 -36198 21923 -35902
rect 21923 -36198 21927 -35902
rect 21623 -36202 21927 -36198
rect 21963 -35902 22587 -35898
rect 21963 -36198 21967 -35902
rect 21967 -36198 22583 -35902
rect 22583 -36198 22587 -35902
rect 21963 -36202 22587 -36198
rect 22623 -35902 22927 -35898
rect 22623 -36198 22627 -35902
rect 22627 -36198 22923 -35902
rect 22923 -36198 22927 -35902
rect 22623 -36202 22927 -36198
rect 22963 -35902 23587 -35898
rect 22963 -36198 22967 -35902
rect 22967 -36198 23583 -35902
rect 23583 -36198 23587 -35902
rect 22963 -36202 23587 -36198
rect 23623 -35902 23927 -35898
rect 23623 -36198 23627 -35902
rect 23627 -36198 23923 -35902
rect 23923 -36198 23927 -35902
rect 23623 -36202 23927 -36198
rect 23963 -35902 24587 -35898
rect 23963 -36198 23967 -35902
rect 23967 -36198 24583 -35902
rect 24583 -36198 24587 -35902
rect 23963 -36202 24587 -36198
rect 24623 -35902 24927 -35898
rect 24623 -36198 24627 -35902
rect 24627 -36198 24923 -35902
rect 24923 -36198 24927 -35902
rect 24623 -36202 24927 -36198
rect 24963 -35902 25587 -35898
rect 24963 -36198 24967 -35902
rect 24967 -36198 25583 -35902
rect 25583 -36198 25587 -35902
rect 24963 -36202 25587 -36198
rect 25623 -35902 25927 -35898
rect 25623 -36198 25627 -35902
rect 25627 -36198 25923 -35902
rect 25923 -36198 25927 -35902
rect 25623 -36202 25927 -36198
rect 25963 -35902 26587 -35898
rect 25963 -36198 25967 -35902
rect 25967 -36198 26583 -35902
rect 26583 -36198 26587 -35902
rect 25963 -36202 26587 -36198
rect 26623 -35902 26927 -35898
rect 26623 -36198 26627 -35902
rect 26627 -36198 26923 -35902
rect 26923 -36198 26927 -35902
rect 26623 -36202 26927 -36198
rect 26963 -35902 27587 -35898
rect 26963 -36198 26967 -35902
rect 26967 -36198 27583 -35902
rect 27583 -36198 27587 -35902
rect 26963 -36202 27587 -36198
rect 27623 -35902 27927 -35898
rect 27623 -36198 27627 -35902
rect 27627 -36198 27923 -35902
rect 27923 -36198 27927 -35902
rect 27623 -36202 27927 -36198
rect 27963 -35902 28587 -35898
rect 27963 -36198 27967 -35902
rect 27967 -36198 28583 -35902
rect 28583 -36198 28587 -35902
rect 27963 -36202 28587 -36198
rect 28623 -35902 28927 -35898
rect 28623 -36198 28627 -35902
rect 28627 -36198 28923 -35902
rect 28923 -36198 28927 -35902
rect 28623 -36202 28927 -36198
rect 28963 -35902 29587 -35898
rect 28963 -36198 28967 -35902
rect 28967 -36198 29583 -35902
rect 29583 -36198 29587 -35902
rect 28963 -36202 29587 -36198
rect 29623 -35902 29927 -35898
rect 29623 -36198 29627 -35902
rect 29627 -36198 29923 -35902
rect 29923 -36198 29927 -35902
rect 29623 -36202 29927 -36198
rect 29963 -35902 30587 -35898
rect 29963 -36198 29967 -35902
rect 29967 -36198 30583 -35902
rect 30583 -36198 30587 -35902
rect 29963 -36202 30587 -36198
rect 30623 -35902 30927 -35898
rect 30623 -36198 30627 -35902
rect 30627 -36198 30923 -35902
rect 30923 -36198 30927 -35902
rect 30623 -36202 30927 -36198
rect 30963 -35902 31587 -35898
rect 30963 -36198 30967 -35902
rect 30967 -36198 31583 -35902
rect 31583 -36198 31587 -35902
rect 30963 -36202 31587 -36198
rect 31623 -35902 31927 -35898
rect 31623 -36198 31627 -35902
rect 31627 -36198 31923 -35902
rect 31923 -36198 31927 -35902
rect 31623 -36202 31927 -36198
rect 31963 -35902 32587 -35898
rect 31963 -36198 31967 -35902
rect 31967 -36198 32583 -35902
rect 32583 -36198 32587 -35902
rect 31963 -36202 32587 -36198
rect 32623 -35902 32927 -35898
rect 32623 -36198 32627 -35902
rect 32627 -36198 32923 -35902
rect 32923 -36198 32927 -35902
rect 32623 -36202 32927 -36198
rect 32963 -35902 33587 -35898
rect 32963 -36198 32967 -35902
rect 32967 -36198 33583 -35902
rect 33583 -36198 33587 -35902
rect 32963 -36202 33587 -36198
rect 33623 -35902 33927 -35898
rect 33623 -36198 33627 -35902
rect 33627 -36198 33923 -35902
rect 33923 -36198 33927 -35902
rect 33623 -36202 33927 -36198
rect 33963 -35902 34267 -35898
rect 33963 -36198 33967 -35902
rect 33967 -36198 34263 -35902
rect 34263 -36198 34267 -35902
rect 33963 -36202 34267 -36198
rect 8623 -36242 8927 -36238
rect 8623 -36858 8627 -36242
rect 8627 -36858 8923 -36242
rect 8923 -36858 8927 -36242
rect 8623 -36862 8927 -36858
rect 9623 -36242 9927 -36238
rect 9623 -36858 9627 -36242
rect 9627 -36858 9923 -36242
rect 9923 -36858 9927 -36242
rect 9623 -36862 9927 -36858
rect 10623 -36242 10927 -36238
rect 10623 -36858 10627 -36242
rect 10627 -36858 10923 -36242
rect 10923 -36858 10927 -36242
rect 10623 -36862 10927 -36858
rect 11623 -36242 11927 -36238
rect 11623 -36858 11627 -36242
rect 11627 -36858 11923 -36242
rect 11923 -36858 11927 -36242
rect 11623 -36862 11927 -36858
rect 12623 -36242 12927 -36238
rect 12623 -36858 12627 -36242
rect 12627 -36858 12923 -36242
rect 12923 -36858 12927 -36242
rect 12623 -36862 12927 -36858
rect 13623 -36242 13927 -36238
rect 13623 -36858 13627 -36242
rect 13627 -36858 13923 -36242
rect 13923 -36858 13927 -36242
rect 13623 -36862 13927 -36858
rect 14623 -36242 14927 -36238
rect 14623 -36858 14627 -36242
rect 14627 -36858 14923 -36242
rect 14923 -36858 14927 -36242
rect 14623 -36862 14927 -36858
rect 15623 -36242 15927 -36238
rect 15623 -36858 15627 -36242
rect 15627 -36858 15923 -36242
rect 15923 -36858 15927 -36242
rect 15623 -36862 15927 -36858
rect 16623 -36242 16927 -36238
rect 16623 -36858 16627 -36242
rect 16627 -36858 16923 -36242
rect 16923 -36858 16927 -36242
rect 16623 -36862 16927 -36858
rect 17623 -36242 17927 -36238
rect 17623 -36858 17627 -36242
rect 17627 -36858 17923 -36242
rect 17923 -36858 17927 -36242
rect 17623 -36862 17927 -36858
rect 18623 -36242 18927 -36238
rect 18623 -36858 18627 -36242
rect 18627 -36858 18923 -36242
rect 18923 -36858 18927 -36242
rect 18623 -36862 18927 -36858
rect 19623 -36242 19927 -36238
rect 19623 -36858 19627 -36242
rect 19627 -36858 19923 -36242
rect 19923 -36858 19927 -36242
rect 19623 -36862 19927 -36858
rect 20623 -36242 20927 -36238
rect 20623 -36858 20627 -36242
rect 20627 -36858 20923 -36242
rect 20923 -36858 20927 -36242
rect 20623 -36862 20927 -36858
rect 21623 -36242 21927 -36238
rect 21623 -36858 21627 -36242
rect 21627 -36858 21923 -36242
rect 21923 -36858 21927 -36242
rect 21623 -36862 21927 -36858
rect 22623 -36242 22927 -36238
rect 22623 -36858 22627 -36242
rect 22627 -36858 22923 -36242
rect 22923 -36858 22927 -36242
rect 22623 -36862 22927 -36858
rect 23623 -36242 23927 -36238
rect 23623 -36858 23627 -36242
rect 23627 -36858 23923 -36242
rect 23923 -36858 23927 -36242
rect 23623 -36862 23927 -36858
rect 24623 -36242 24927 -36238
rect 24623 -36858 24627 -36242
rect 24627 -36858 24923 -36242
rect 24923 -36858 24927 -36242
rect 24623 -36862 24927 -36858
rect 25623 -36242 25927 -36238
rect 25623 -36858 25627 -36242
rect 25627 -36858 25923 -36242
rect 25923 -36858 25927 -36242
rect 25623 -36862 25927 -36858
rect 26623 -36242 26927 -36238
rect 26623 -36858 26627 -36242
rect 26627 -36858 26923 -36242
rect 26923 -36858 26927 -36242
rect 26623 -36862 26927 -36858
rect 27623 -36242 27927 -36238
rect 27623 -36858 27627 -36242
rect 27627 -36858 27923 -36242
rect 27923 -36858 27927 -36242
rect 27623 -36862 27927 -36858
rect 28623 -36242 28927 -36238
rect 28623 -36858 28627 -36242
rect 28627 -36858 28923 -36242
rect 28923 -36858 28927 -36242
rect 28623 -36862 28927 -36858
rect 29623 -36242 29927 -36238
rect 29623 -36858 29627 -36242
rect 29627 -36858 29923 -36242
rect 29923 -36858 29927 -36242
rect 29623 -36862 29927 -36858
rect 30623 -36242 30927 -36238
rect 30623 -36858 30627 -36242
rect 30627 -36858 30923 -36242
rect 30923 -36858 30927 -36242
rect 30623 -36862 30927 -36858
rect 31623 -36242 31927 -36238
rect 31623 -36858 31627 -36242
rect 31627 -36858 31923 -36242
rect 31923 -36858 31927 -36242
rect 31623 -36862 31927 -36858
rect 32623 -36242 32927 -36238
rect 32623 -36858 32627 -36242
rect 32627 -36858 32923 -36242
rect 32923 -36858 32927 -36242
rect 32623 -36862 32927 -36858
rect 33623 -36242 33927 -36238
rect 33623 -36858 33627 -36242
rect 33627 -36858 33923 -36242
rect 33923 -36858 33927 -36242
rect 33623 -36862 33927 -36858
rect 8283 -36902 8587 -36898
rect 8283 -37198 8287 -36902
rect 8287 -37198 8583 -36902
rect 8583 -37198 8587 -36902
rect 8283 -37202 8587 -37198
rect 8623 -36902 8927 -36898
rect 8623 -37198 8627 -36902
rect 8627 -37198 8923 -36902
rect 8923 -37198 8927 -36902
rect 8623 -37202 8927 -37198
rect 8963 -36902 9587 -36898
rect 8963 -37198 8967 -36902
rect 8967 -37198 9583 -36902
rect 9583 -37198 9587 -36902
rect 8963 -37202 9587 -37198
rect 9623 -36902 9927 -36898
rect 9623 -37198 9627 -36902
rect 9627 -37198 9923 -36902
rect 9923 -37198 9927 -36902
rect 9623 -37202 9927 -37198
rect 9963 -36902 10587 -36898
rect 9963 -37198 9967 -36902
rect 9967 -37198 10583 -36902
rect 10583 -37198 10587 -36902
rect 9963 -37202 10587 -37198
rect 10623 -36902 10927 -36898
rect 10623 -37198 10627 -36902
rect 10627 -37198 10923 -36902
rect 10923 -37198 10927 -36902
rect 10623 -37202 10927 -37198
rect 10963 -36902 11587 -36898
rect 10963 -37198 10967 -36902
rect 10967 -37198 11583 -36902
rect 11583 -37198 11587 -36902
rect 10963 -37202 11587 -37198
rect 11623 -36902 11927 -36898
rect 11623 -37198 11627 -36902
rect 11627 -37198 11923 -36902
rect 11923 -37198 11927 -36902
rect 11623 -37202 11927 -37198
rect 11963 -36902 12587 -36898
rect 11963 -37198 11967 -36902
rect 11967 -37198 12583 -36902
rect 12583 -37198 12587 -36902
rect 11963 -37202 12587 -37198
rect 12623 -36902 12927 -36898
rect 12623 -37198 12627 -36902
rect 12627 -37198 12923 -36902
rect 12923 -37198 12927 -36902
rect 12623 -37202 12927 -37198
rect 12963 -36902 13587 -36898
rect 12963 -37198 12967 -36902
rect 12967 -37198 13583 -36902
rect 13583 -37198 13587 -36902
rect 12963 -37202 13587 -37198
rect 13623 -36902 13927 -36898
rect 13623 -37198 13627 -36902
rect 13627 -37198 13923 -36902
rect 13923 -37198 13927 -36902
rect 13623 -37202 13927 -37198
rect 13963 -36902 14587 -36898
rect 13963 -37198 13967 -36902
rect 13967 -37198 14583 -36902
rect 14583 -37198 14587 -36902
rect 13963 -37202 14587 -37198
rect 14623 -36902 14927 -36898
rect 14623 -37198 14627 -36902
rect 14627 -37198 14923 -36902
rect 14923 -37198 14927 -36902
rect 14623 -37202 14927 -37198
rect 14963 -36902 15587 -36898
rect 14963 -37198 14967 -36902
rect 14967 -37198 15583 -36902
rect 15583 -37198 15587 -36902
rect 14963 -37202 15587 -37198
rect 15623 -36902 15927 -36898
rect 15623 -37198 15627 -36902
rect 15627 -37198 15923 -36902
rect 15923 -37198 15927 -36902
rect 15623 -37202 15927 -37198
rect 15963 -36902 16587 -36898
rect 15963 -37198 15967 -36902
rect 15967 -37198 16583 -36902
rect 16583 -37198 16587 -36902
rect 15963 -37202 16587 -37198
rect 16623 -36902 16927 -36898
rect 16623 -37198 16627 -36902
rect 16627 -37198 16923 -36902
rect 16923 -37198 16927 -36902
rect 16623 -37202 16927 -37198
rect 16963 -36902 17587 -36898
rect 16963 -37198 16967 -36902
rect 16967 -37198 17583 -36902
rect 17583 -37198 17587 -36902
rect 16963 -37202 17587 -37198
rect 17623 -36902 17927 -36898
rect 17623 -37198 17627 -36902
rect 17627 -37198 17923 -36902
rect 17923 -37198 17927 -36902
rect 17623 -37202 17927 -37198
rect 17963 -36902 18587 -36898
rect 17963 -37198 17967 -36902
rect 17967 -37198 18583 -36902
rect 18583 -37198 18587 -36902
rect 17963 -37202 18587 -37198
rect 18623 -36902 18927 -36898
rect 18623 -37198 18627 -36902
rect 18627 -37198 18923 -36902
rect 18923 -37198 18927 -36902
rect 18623 -37202 18927 -37198
rect 18963 -36902 19587 -36898
rect 18963 -37198 18967 -36902
rect 18967 -37198 19583 -36902
rect 19583 -37198 19587 -36902
rect 18963 -37202 19587 -37198
rect 19623 -36902 19927 -36898
rect 19623 -37198 19627 -36902
rect 19627 -37198 19923 -36902
rect 19923 -37198 19927 -36902
rect 19623 -37202 19927 -37198
rect 19963 -36902 20587 -36898
rect 19963 -37198 19967 -36902
rect 19967 -37198 20583 -36902
rect 20583 -37198 20587 -36902
rect 19963 -37202 20587 -37198
rect 20623 -36902 20927 -36898
rect 20623 -37198 20627 -36902
rect 20627 -37198 20923 -36902
rect 20923 -37198 20927 -36902
rect 20623 -37202 20927 -37198
rect 20963 -36902 21587 -36898
rect 20963 -37198 20967 -36902
rect 20967 -37198 21583 -36902
rect 21583 -37198 21587 -36902
rect 20963 -37202 21587 -37198
rect 21623 -36902 21927 -36898
rect 21623 -37198 21627 -36902
rect 21627 -37198 21923 -36902
rect 21923 -37198 21927 -36902
rect 21623 -37202 21927 -37198
rect 21963 -36902 22587 -36898
rect 21963 -37198 21967 -36902
rect 21967 -37198 22583 -36902
rect 22583 -37198 22587 -36902
rect 21963 -37202 22587 -37198
rect 22623 -36902 22927 -36898
rect 22623 -37198 22627 -36902
rect 22627 -37198 22923 -36902
rect 22923 -37198 22927 -36902
rect 22623 -37202 22927 -37198
rect 22963 -36902 23587 -36898
rect 22963 -37198 22967 -36902
rect 22967 -37198 23583 -36902
rect 23583 -37198 23587 -36902
rect 22963 -37202 23587 -37198
rect 23623 -36902 23927 -36898
rect 23623 -37198 23627 -36902
rect 23627 -37198 23923 -36902
rect 23923 -37198 23927 -36902
rect 23623 -37202 23927 -37198
rect 23963 -36902 24587 -36898
rect 23963 -37198 23967 -36902
rect 23967 -37198 24583 -36902
rect 24583 -37198 24587 -36902
rect 23963 -37202 24587 -37198
rect 24623 -36902 24927 -36898
rect 24623 -37198 24627 -36902
rect 24627 -37198 24923 -36902
rect 24923 -37198 24927 -36902
rect 24623 -37202 24927 -37198
rect 24963 -36902 25587 -36898
rect 24963 -37198 24967 -36902
rect 24967 -37198 25583 -36902
rect 25583 -37198 25587 -36902
rect 24963 -37202 25587 -37198
rect 25623 -36902 25927 -36898
rect 25623 -37198 25627 -36902
rect 25627 -37198 25923 -36902
rect 25923 -37198 25927 -36902
rect 25623 -37202 25927 -37198
rect 25963 -36902 26587 -36898
rect 25963 -37198 25967 -36902
rect 25967 -37198 26583 -36902
rect 26583 -37198 26587 -36902
rect 25963 -37202 26587 -37198
rect 26623 -36902 26927 -36898
rect 26623 -37198 26627 -36902
rect 26627 -37198 26923 -36902
rect 26923 -37198 26927 -36902
rect 26623 -37202 26927 -37198
rect 26963 -36902 27587 -36898
rect 26963 -37198 26967 -36902
rect 26967 -37198 27583 -36902
rect 27583 -37198 27587 -36902
rect 26963 -37202 27587 -37198
rect 27623 -36902 27927 -36898
rect 27623 -37198 27627 -36902
rect 27627 -37198 27923 -36902
rect 27923 -37198 27927 -36902
rect 27623 -37202 27927 -37198
rect 27963 -36902 28587 -36898
rect 27963 -37198 27967 -36902
rect 27967 -37198 28583 -36902
rect 28583 -37198 28587 -36902
rect 27963 -37202 28587 -37198
rect 28623 -36902 28927 -36898
rect 28623 -37198 28627 -36902
rect 28627 -37198 28923 -36902
rect 28923 -37198 28927 -36902
rect 28623 -37202 28927 -37198
rect 28963 -36902 29587 -36898
rect 28963 -37198 28967 -36902
rect 28967 -37198 29583 -36902
rect 29583 -37198 29587 -36902
rect 28963 -37202 29587 -37198
rect 29623 -36902 29927 -36898
rect 29623 -37198 29627 -36902
rect 29627 -37198 29923 -36902
rect 29923 -37198 29927 -36902
rect 29623 -37202 29927 -37198
rect 29963 -36902 30587 -36898
rect 29963 -37198 29967 -36902
rect 29967 -37198 30583 -36902
rect 30583 -37198 30587 -36902
rect 29963 -37202 30587 -37198
rect 30623 -36902 30927 -36898
rect 30623 -37198 30627 -36902
rect 30627 -37198 30923 -36902
rect 30923 -37198 30927 -36902
rect 30623 -37202 30927 -37198
rect 30963 -36902 31587 -36898
rect 30963 -37198 30967 -36902
rect 30967 -37198 31583 -36902
rect 31583 -37198 31587 -36902
rect 30963 -37202 31587 -37198
rect 31623 -36902 31927 -36898
rect 31623 -37198 31627 -36902
rect 31627 -37198 31923 -36902
rect 31923 -37198 31927 -36902
rect 31623 -37202 31927 -37198
rect 31963 -36902 32587 -36898
rect 31963 -37198 31967 -36902
rect 31967 -37198 32583 -36902
rect 32583 -37198 32587 -36902
rect 31963 -37202 32587 -37198
rect 32623 -36902 32927 -36898
rect 32623 -37198 32627 -36902
rect 32627 -37198 32923 -36902
rect 32923 -37198 32927 -36902
rect 32623 -37202 32927 -37198
rect 32963 -36902 33587 -36898
rect 32963 -37198 32967 -36902
rect 32967 -37198 33583 -36902
rect 33583 -37198 33587 -36902
rect 32963 -37202 33587 -37198
rect 33623 -36902 33927 -36898
rect 33623 -37198 33627 -36902
rect 33627 -37198 33923 -36902
rect 33923 -37198 33927 -36902
rect 33623 -37202 33927 -37198
rect 33963 -36902 34267 -36898
rect 33963 -37198 33967 -36902
rect 33967 -37198 34263 -36902
rect 34263 -37198 34267 -36902
rect 33963 -37202 34267 -37198
rect 8623 -37242 8927 -37238
rect 8623 -37858 8627 -37242
rect 8627 -37858 8923 -37242
rect 8923 -37858 8927 -37242
rect 8623 -37862 8927 -37858
rect 9623 -37242 9927 -37238
rect 9623 -37858 9627 -37242
rect 9627 -37858 9923 -37242
rect 9923 -37858 9927 -37242
rect 9623 -37862 9927 -37858
rect 10623 -37242 10927 -37238
rect 10623 -37858 10627 -37242
rect 10627 -37858 10923 -37242
rect 10923 -37858 10927 -37242
rect 10623 -37862 10927 -37858
rect 11623 -37242 11927 -37238
rect 11623 -37858 11627 -37242
rect 11627 -37858 11923 -37242
rect 11923 -37858 11927 -37242
rect 11623 -37862 11927 -37858
rect 12623 -37242 12927 -37238
rect 12623 -37858 12627 -37242
rect 12627 -37858 12923 -37242
rect 12923 -37858 12927 -37242
rect 12623 -37862 12927 -37858
rect 13623 -37242 13927 -37238
rect 13623 -37858 13627 -37242
rect 13627 -37858 13923 -37242
rect 13923 -37858 13927 -37242
rect 13623 -37862 13927 -37858
rect 14623 -37242 14927 -37238
rect 14623 -37858 14627 -37242
rect 14627 -37858 14923 -37242
rect 14923 -37858 14927 -37242
rect 14623 -37862 14927 -37858
rect 15623 -37242 15927 -37238
rect 15623 -37858 15627 -37242
rect 15627 -37858 15923 -37242
rect 15923 -37858 15927 -37242
rect 15623 -37862 15927 -37858
rect 16623 -37242 16927 -37238
rect 16623 -37858 16627 -37242
rect 16627 -37858 16923 -37242
rect 16923 -37858 16927 -37242
rect 16623 -37862 16927 -37858
rect 17623 -37242 17927 -37238
rect 17623 -37858 17627 -37242
rect 17627 -37858 17923 -37242
rect 17923 -37858 17927 -37242
rect 17623 -37862 17927 -37858
rect 18623 -37242 18927 -37238
rect 18623 -37858 18627 -37242
rect 18627 -37858 18923 -37242
rect 18923 -37858 18927 -37242
rect 18623 -37862 18927 -37858
rect 19623 -37242 19927 -37238
rect 19623 -37858 19627 -37242
rect 19627 -37858 19923 -37242
rect 19923 -37858 19927 -37242
rect 19623 -37862 19927 -37858
rect 20623 -37242 20927 -37238
rect 20623 -37858 20627 -37242
rect 20627 -37858 20923 -37242
rect 20923 -37858 20927 -37242
rect 20623 -37862 20927 -37858
rect 21623 -37242 21927 -37238
rect 21623 -37858 21627 -37242
rect 21627 -37858 21923 -37242
rect 21923 -37858 21927 -37242
rect 21623 -37862 21927 -37858
rect 22623 -37242 22927 -37238
rect 22623 -37858 22627 -37242
rect 22627 -37858 22923 -37242
rect 22923 -37858 22927 -37242
rect 22623 -37862 22927 -37858
rect 23623 -37242 23927 -37238
rect 23623 -37858 23627 -37242
rect 23627 -37858 23923 -37242
rect 23923 -37858 23927 -37242
rect 23623 -37862 23927 -37858
rect 24623 -37242 24927 -37238
rect 24623 -37858 24627 -37242
rect 24627 -37858 24923 -37242
rect 24923 -37858 24927 -37242
rect 24623 -37862 24927 -37858
rect 25623 -37242 25927 -37238
rect 25623 -37858 25627 -37242
rect 25627 -37858 25923 -37242
rect 25923 -37858 25927 -37242
rect 25623 -37862 25927 -37858
rect 26623 -37242 26927 -37238
rect 26623 -37858 26627 -37242
rect 26627 -37858 26923 -37242
rect 26923 -37858 26927 -37242
rect 26623 -37862 26927 -37858
rect 27623 -37242 27927 -37238
rect 27623 -37858 27627 -37242
rect 27627 -37858 27923 -37242
rect 27923 -37858 27927 -37242
rect 27623 -37862 27927 -37858
rect 28623 -37242 28927 -37238
rect 28623 -37858 28627 -37242
rect 28627 -37858 28923 -37242
rect 28923 -37858 28927 -37242
rect 28623 -37862 28927 -37858
rect 29623 -37242 29927 -37238
rect 29623 -37858 29627 -37242
rect 29627 -37858 29923 -37242
rect 29923 -37858 29927 -37242
rect 29623 -37862 29927 -37858
rect 30623 -37242 30927 -37238
rect 30623 -37858 30627 -37242
rect 30627 -37858 30923 -37242
rect 30923 -37858 30927 -37242
rect 30623 -37862 30927 -37858
rect 31623 -37242 31927 -37238
rect 31623 -37858 31627 -37242
rect 31627 -37858 31923 -37242
rect 31923 -37858 31927 -37242
rect 31623 -37862 31927 -37858
rect 32623 -37242 32927 -37238
rect 32623 -37858 32627 -37242
rect 32627 -37858 32923 -37242
rect 32923 -37858 32927 -37242
rect 32623 -37862 32927 -37858
rect 33623 -37242 33927 -37238
rect 33623 -37858 33627 -37242
rect 33627 -37858 33923 -37242
rect 33923 -37858 33927 -37242
rect 33623 -37862 33927 -37858
rect 8283 -37902 8587 -37898
rect 8283 -38198 8287 -37902
rect 8287 -38198 8583 -37902
rect 8583 -38198 8587 -37902
rect 8283 -38202 8587 -38198
rect 8623 -37902 8927 -37898
rect 8623 -38198 8627 -37902
rect 8627 -38198 8923 -37902
rect 8923 -38198 8927 -37902
rect 8623 -38202 8927 -38198
rect 8963 -37902 9587 -37898
rect 8963 -38198 8967 -37902
rect 8967 -38198 9583 -37902
rect 9583 -38198 9587 -37902
rect 8963 -38202 9587 -38198
rect 9623 -37902 9927 -37898
rect 9623 -38198 9627 -37902
rect 9627 -38198 9923 -37902
rect 9923 -38198 9927 -37902
rect 9623 -38202 9927 -38198
rect 9963 -37902 10587 -37898
rect 9963 -38198 9967 -37902
rect 9967 -38198 10583 -37902
rect 10583 -38198 10587 -37902
rect 9963 -38202 10587 -38198
rect 10623 -37902 10927 -37898
rect 10623 -38198 10627 -37902
rect 10627 -38198 10923 -37902
rect 10923 -38198 10927 -37902
rect 10623 -38202 10927 -38198
rect 10963 -37902 11587 -37898
rect 10963 -38198 10967 -37902
rect 10967 -38198 11583 -37902
rect 11583 -38198 11587 -37902
rect 10963 -38202 11587 -38198
rect 11623 -37902 11927 -37898
rect 11623 -38198 11627 -37902
rect 11627 -38198 11923 -37902
rect 11923 -38198 11927 -37902
rect 11623 -38202 11927 -38198
rect 11963 -37902 12587 -37898
rect 11963 -38198 11967 -37902
rect 11967 -38198 12583 -37902
rect 12583 -38198 12587 -37902
rect 11963 -38202 12587 -38198
rect 12623 -37902 12927 -37898
rect 12623 -38198 12627 -37902
rect 12627 -38198 12923 -37902
rect 12923 -38198 12927 -37902
rect 12623 -38202 12927 -38198
rect 12963 -37902 13587 -37898
rect 12963 -38198 12967 -37902
rect 12967 -38198 13583 -37902
rect 13583 -38198 13587 -37902
rect 12963 -38202 13587 -38198
rect 13623 -37902 13927 -37898
rect 13623 -38198 13627 -37902
rect 13627 -38198 13923 -37902
rect 13923 -38198 13927 -37902
rect 13623 -38202 13927 -38198
rect 13963 -37902 14587 -37898
rect 13963 -38198 13967 -37902
rect 13967 -38198 14583 -37902
rect 14583 -38198 14587 -37902
rect 13963 -38202 14587 -38198
rect 14623 -37902 14927 -37898
rect 14623 -38198 14627 -37902
rect 14627 -38198 14923 -37902
rect 14923 -38198 14927 -37902
rect 14623 -38202 14927 -38198
rect 14963 -37902 15587 -37898
rect 14963 -38198 14967 -37902
rect 14967 -38198 15583 -37902
rect 15583 -38198 15587 -37902
rect 14963 -38202 15587 -38198
rect 15623 -37902 15927 -37898
rect 15623 -38198 15627 -37902
rect 15627 -38198 15923 -37902
rect 15923 -38198 15927 -37902
rect 15623 -38202 15927 -38198
rect 15963 -37902 16587 -37898
rect 15963 -38198 15967 -37902
rect 15967 -38198 16583 -37902
rect 16583 -38198 16587 -37902
rect 15963 -38202 16587 -38198
rect 16623 -37902 16927 -37898
rect 16623 -38198 16627 -37902
rect 16627 -38198 16923 -37902
rect 16923 -38198 16927 -37902
rect 16623 -38202 16927 -38198
rect 16963 -37902 17587 -37898
rect 16963 -38198 16967 -37902
rect 16967 -38198 17583 -37902
rect 17583 -38198 17587 -37902
rect 16963 -38202 17587 -38198
rect 17623 -37902 17927 -37898
rect 17623 -38198 17627 -37902
rect 17627 -38198 17923 -37902
rect 17923 -38198 17927 -37902
rect 17623 -38202 17927 -38198
rect 17963 -37902 18587 -37898
rect 17963 -38198 17967 -37902
rect 17967 -38198 18583 -37902
rect 18583 -38198 18587 -37902
rect 17963 -38202 18587 -38198
rect 18623 -37902 18927 -37898
rect 18623 -38198 18627 -37902
rect 18627 -38198 18923 -37902
rect 18923 -38198 18927 -37902
rect 18623 -38202 18927 -38198
rect 18963 -37902 19587 -37898
rect 18963 -38198 18967 -37902
rect 18967 -38198 19583 -37902
rect 19583 -38198 19587 -37902
rect 18963 -38202 19587 -38198
rect 19623 -37902 19927 -37898
rect 19623 -38198 19627 -37902
rect 19627 -38198 19923 -37902
rect 19923 -38198 19927 -37902
rect 19623 -38202 19927 -38198
rect 19963 -37902 20587 -37898
rect 19963 -38198 19967 -37902
rect 19967 -38198 20583 -37902
rect 20583 -38198 20587 -37902
rect 19963 -38202 20587 -38198
rect 20623 -37902 20927 -37898
rect 20623 -38198 20627 -37902
rect 20627 -38198 20923 -37902
rect 20923 -38198 20927 -37902
rect 20623 -38202 20927 -38198
rect 20963 -37902 21587 -37898
rect 20963 -38198 20967 -37902
rect 20967 -38198 21583 -37902
rect 21583 -38198 21587 -37902
rect 20963 -38202 21587 -38198
rect 21623 -37902 21927 -37898
rect 21623 -38198 21627 -37902
rect 21627 -38198 21923 -37902
rect 21923 -38198 21927 -37902
rect 21623 -38202 21927 -38198
rect 21963 -37902 22587 -37898
rect 21963 -38198 21967 -37902
rect 21967 -38198 22583 -37902
rect 22583 -38198 22587 -37902
rect 21963 -38202 22587 -38198
rect 22623 -37902 22927 -37898
rect 22623 -38198 22627 -37902
rect 22627 -38198 22923 -37902
rect 22923 -38198 22927 -37902
rect 22623 -38202 22927 -38198
rect 22963 -37902 23587 -37898
rect 22963 -38198 22967 -37902
rect 22967 -38198 23583 -37902
rect 23583 -38198 23587 -37902
rect 22963 -38202 23587 -38198
rect 23623 -37902 23927 -37898
rect 23623 -38198 23627 -37902
rect 23627 -38198 23923 -37902
rect 23923 -38198 23927 -37902
rect 23623 -38202 23927 -38198
rect 23963 -37902 24587 -37898
rect 23963 -38198 23967 -37902
rect 23967 -38198 24583 -37902
rect 24583 -38198 24587 -37902
rect 23963 -38202 24587 -38198
rect 24623 -37902 24927 -37898
rect 24623 -38198 24627 -37902
rect 24627 -38198 24923 -37902
rect 24923 -38198 24927 -37902
rect 24623 -38202 24927 -38198
rect 24963 -37902 25587 -37898
rect 24963 -38198 24967 -37902
rect 24967 -38198 25583 -37902
rect 25583 -38198 25587 -37902
rect 24963 -38202 25587 -38198
rect 25623 -37902 25927 -37898
rect 25623 -38198 25627 -37902
rect 25627 -38198 25923 -37902
rect 25923 -38198 25927 -37902
rect 25623 -38202 25927 -38198
rect 25963 -37902 26587 -37898
rect 25963 -38198 25967 -37902
rect 25967 -38198 26583 -37902
rect 26583 -38198 26587 -37902
rect 25963 -38202 26587 -38198
rect 26623 -37902 26927 -37898
rect 26623 -38198 26627 -37902
rect 26627 -38198 26923 -37902
rect 26923 -38198 26927 -37902
rect 26623 -38202 26927 -38198
rect 26963 -37902 27587 -37898
rect 26963 -38198 26967 -37902
rect 26967 -38198 27583 -37902
rect 27583 -38198 27587 -37902
rect 26963 -38202 27587 -38198
rect 27623 -37902 27927 -37898
rect 27623 -38198 27627 -37902
rect 27627 -38198 27923 -37902
rect 27923 -38198 27927 -37902
rect 27623 -38202 27927 -38198
rect 27963 -37902 28587 -37898
rect 27963 -38198 27967 -37902
rect 27967 -38198 28583 -37902
rect 28583 -38198 28587 -37902
rect 27963 -38202 28587 -38198
rect 28623 -37902 28927 -37898
rect 28623 -38198 28627 -37902
rect 28627 -38198 28923 -37902
rect 28923 -38198 28927 -37902
rect 28623 -38202 28927 -38198
rect 28963 -37902 29587 -37898
rect 28963 -38198 28967 -37902
rect 28967 -38198 29583 -37902
rect 29583 -38198 29587 -37902
rect 28963 -38202 29587 -38198
rect 29623 -37902 29927 -37898
rect 29623 -38198 29627 -37902
rect 29627 -38198 29923 -37902
rect 29923 -38198 29927 -37902
rect 29623 -38202 29927 -38198
rect 29963 -37902 30587 -37898
rect 29963 -38198 29967 -37902
rect 29967 -38198 30583 -37902
rect 30583 -38198 30587 -37902
rect 29963 -38202 30587 -38198
rect 30623 -37902 30927 -37898
rect 30623 -38198 30627 -37902
rect 30627 -38198 30923 -37902
rect 30923 -38198 30927 -37902
rect 30623 -38202 30927 -38198
rect 30963 -37902 31587 -37898
rect 30963 -38198 30967 -37902
rect 30967 -38198 31583 -37902
rect 31583 -38198 31587 -37902
rect 30963 -38202 31587 -38198
rect 31623 -37902 31927 -37898
rect 31623 -38198 31627 -37902
rect 31627 -38198 31923 -37902
rect 31923 -38198 31927 -37902
rect 31623 -38202 31927 -38198
rect 31963 -37902 32587 -37898
rect 31963 -38198 31967 -37902
rect 31967 -38198 32583 -37902
rect 32583 -38198 32587 -37902
rect 31963 -38202 32587 -38198
rect 32623 -37902 32927 -37898
rect 32623 -38198 32627 -37902
rect 32627 -38198 32923 -37902
rect 32923 -38198 32927 -37902
rect 32623 -38202 32927 -38198
rect 32963 -37902 33587 -37898
rect 32963 -38198 32967 -37902
rect 32967 -38198 33583 -37902
rect 33583 -38198 33587 -37902
rect 32963 -38202 33587 -38198
rect 33623 -37902 33927 -37898
rect 33623 -38198 33627 -37902
rect 33627 -38198 33923 -37902
rect 33923 -38198 33927 -37902
rect 33623 -38202 33927 -38198
rect 33963 -37902 34267 -37898
rect 33963 -38198 33967 -37902
rect 33967 -38198 34263 -37902
rect 34263 -38198 34267 -37902
rect 33963 -38202 34267 -38198
rect 8623 -38242 8927 -38238
rect 8623 -38858 8627 -38242
rect 8627 -38858 8923 -38242
rect 8923 -38858 8927 -38242
rect 8623 -38862 8927 -38858
rect 9623 -38242 9927 -38238
rect 9623 -38858 9627 -38242
rect 9627 -38858 9923 -38242
rect 9923 -38858 9927 -38242
rect 9623 -38862 9927 -38858
rect 10623 -38242 10927 -38238
rect 10623 -38858 10627 -38242
rect 10627 -38858 10923 -38242
rect 10923 -38858 10927 -38242
rect 10623 -38862 10927 -38858
rect 11623 -38242 11927 -38238
rect 11623 -38858 11627 -38242
rect 11627 -38858 11923 -38242
rect 11923 -38858 11927 -38242
rect 11623 -38862 11927 -38858
rect 12623 -38242 12927 -38238
rect 12623 -38858 12627 -38242
rect 12627 -38858 12923 -38242
rect 12923 -38858 12927 -38242
rect 12623 -38862 12927 -38858
rect 13623 -38242 13927 -38238
rect 13623 -38858 13627 -38242
rect 13627 -38858 13923 -38242
rect 13923 -38858 13927 -38242
rect 13623 -38862 13927 -38858
rect 14623 -38242 14927 -38238
rect 14623 -38858 14627 -38242
rect 14627 -38858 14923 -38242
rect 14923 -38858 14927 -38242
rect 14623 -38862 14927 -38858
rect 15623 -38242 15927 -38238
rect 15623 -38858 15627 -38242
rect 15627 -38858 15923 -38242
rect 15923 -38858 15927 -38242
rect 15623 -38862 15927 -38858
rect 16623 -38242 16927 -38238
rect 16623 -38858 16627 -38242
rect 16627 -38858 16923 -38242
rect 16923 -38858 16927 -38242
rect 16623 -38862 16927 -38858
rect 17623 -38242 17927 -38238
rect 17623 -38858 17627 -38242
rect 17627 -38858 17923 -38242
rect 17923 -38858 17927 -38242
rect 17623 -38862 17927 -38858
rect 18623 -38242 18927 -38238
rect 18623 -38858 18627 -38242
rect 18627 -38858 18923 -38242
rect 18923 -38858 18927 -38242
rect 18623 -38862 18927 -38858
rect 19623 -38242 19927 -38238
rect 19623 -38858 19627 -38242
rect 19627 -38858 19923 -38242
rect 19923 -38858 19927 -38242
rect 19623 -38862 19927 -38858
rect 20623 -38242 20927 -38238
rect 20623 -38858 20627 -38242
rect 20627 -38858 20923 -38242
rect 20923 -38858 20927 -38242
rect 20623 -38862 20927 -38858
rect 21623 -38242 21927 -38238
rect 21623 -38858 21627 -38242
rect 21627 -38858 21923 -38242
rect 21923 -38858 21927 -38242
rect 21623 -38862 21927 -38858
rect 22623 -38242 22927 -38238
rect 22623 -38858 22627 -38242
rect 22627 -38858 22923 -38242
rect 22923 -38858 22927 -38242
rect 22623 -38862 22927 -38858
rect 23623 -38242 23927 -38238
rect 23623 -38858 23627 -38242
rect 23627 -38858 23923 -38242
rect 23923 -38858 23927 -38242
rect 23623 -38862 23927 -38858
rect 24623 -38242 24927 -38238
rect 24623 -38858 24627 -38242
rect 24627 -38858 24923 -38242
rect 24923 -38858 24927 -38242
rect 24623 -38862 24927 -38858
rect 25623 -38242 25927 -38238
rect 25623 -38858 25627 -38242
rect 25627 -38858 25923 -38242
rect 25923 -38858 25927 -38242
rect 25623 -38862 25927 -38858
rect 26623 -38242 26927 -38238
rect 26623 -38858 26627 -38242
rect 26627 -38858 26923 -38242
rect 26923 -38858 26927 -38242
rect 26623 -38862 26927 -38858
rect 27623 -38242 27927 -38238
rect 27623 -38858 27627 -38242
rect 27627 -38858 27923 -38242
rect 27923 -38858 27927 -38242
rect 27623 -38862 27927 -38858
rect 28623 -38242 28927 -38238
rect 28623 -38858 28627 -38242
rect 28627 -38858 28923 -38242
rect 28923 -38858 28927 -38242
rect 28623 -38862 28927 -38858
rect 29623 -38242 29927 -38238
rect 29623 -38858 29627 -38242
rect 29627 -38858 29923 -38242
rect 29923 -38858 29927 -38242
rect 29623 -38862 29927 -38858
rect 30623 -38242 30927 -38238
rect 30623 -38858 30627 -38242
rect 30627 -38858 30923 -38242
rect 30923 -38858 30927 -38242
rect 30623 -38862 30927 -38858
rect 31623 -38242 31927 -38238
rect 31623 -38858 31627 -38242
rect 31627 -38858 31923 -38242
rect 31923 -38858 31927 -38242
rect 31623 -38862 31927 -38858
rect 32623 -38242 32927 -38238
rect 32623 -38858 32627 -38242
rect 32627 -38858 32923 -38242
rect 32923 -38858 32927 -38242
rect 32623 -38862 32927 -38858
rect 33623 -38242 33927 -38238
rect 33623 -38858 33627 -38242
rect 33627 -38858 33923 -38242
rect 33923 -38858 33927 -38242
rect 33623 -38862 33927 -38858
rect 8283 -38902 8587 -38898
rect 8283 -39198 8287 -38902
rect 8287 -39198 8583 -38902
rect 8583 -39198 8587 -38902
rect 8283 -39202 8587 -39198
rect 8623 -38902 8927 -38898
rect 8623 -39198 8627 -38902
rect 8627 -39198 8923 -38902
rect 8923 -39198 8927 -38902
rect 8623 -39202 8927 -39198
rect 8963 -38902 9587 -38898
rect 8963 -39198 8967 -38902
rect 8967 -39198 9583 -38902
rect 9583 -39198 9587 -38902
rect 8963 -39202 9587 -39198
rect 9623 -38902 9927 -38898
rect 9623 -39198 9627 -38902
rect 9627 -39198 9923 -38902
rect 9923 -39198 9927 -38902
rect 9623 -39202 9927 -39198
rect 9963 -38902 10587 -38898
rect 9963 -39198 9967 -38902
rect 9967 -39198 10583 -38902
rect 10583 -39198 10587 -38902
rect 9963 -39202 10587 -39198
rect 10623 -38902 10927 -38898
rect 10623 -39198 10627 -38902
rect 10627 -39198 10923 -38902
rect 10923 -39198 10927 -38902
rect 10623 -39202 10927 -39198
rect 10963 -38902 11587 -38898
rect 10963 -39198 10967 -38902
rect 10967 -39198 11583 -38902
rect 11583 -39198 11587 -38902
rect 10963 -39202 11587 -39198
rect 11623 -38902 11927 -38898
rect 11623 -39198 11627 -38902
rect 11627 -39198 11923 -38902
rect 11923 -39198 11927 -38902
rect 11623 -39202 11927 -39198
rect 11963 -38902 12587 -38898
rect 11963 -39198 11967 -38902
rect 11967 -39198 12583 -38902
rect 12583 -39198 12587 -38902
rect 11963 -39202 12587 -39198
rect 12623 -38902 12927 -38898
rect 12623 -39198 12627 -38902
rect 12627 -39198 12923 -38902
rect 12923 -39198 12927 -38902
rect 12623 -39202 12927 -39198
rect 12963 -38902 13587 -38898
rect 12963 -39198 12967 -38902
rect 12967 -39198 13583 -38902
rect 13583 -39198 13587 -38902
rect 12963 -39202 13587 -39198
rect 13623 -38902 13927 -38898
rect 13623 -39198 13627 -38902
rect 13627 -39198 13923 -38902
rect 13923 -39198 13927 -38902
rect 13623 -39202 13927 -39198
rect 13963 -38902 14587 -38898
rect 13963 -39198 13967 -38902
rect 13967 -39198 14583 -38902
rect 14583 -39198 14587 -38902
rect 13963 -39202 14587 -39198
rect 14623 -38902 14927 -38898
rect 14623 -39198 14627 -38902
rect 14627 -39198 14923 -38902
rect 14923 -39198 14927 -38902
rect 14623 -39202 14927 -39198
rect 14963 -38902 15587 -38898
rect 14963 -39198 14967 -38902
rect 14967 -39198 15583 -38902
rect 15583 -39198 15587 -38902
rect 14963 -39202 15587 -39198
rect 15623 -38902 15927 -38898
rect 15623 -39198 15627 -38902
rect 15627 -39198 15923 -38902
rect 15923 -39198 15927 -38902
rect 15623 -39202 15927 -39198
rect 15963 -38902 16587 -38898
rect 15963 -39198 15967 -38902
rect 15967 -39198 16583 -38902
rect 16583 -39198 16587 -38902
rect 15963 -39202 16587 -39198
rect 16623 -38902 16927 -38898
rect 16623 -39198 16627 -38902
rect 16627 -39198 16923 -38902
rect 16923 -39198 16927 -38902
rect 16623 -39202 16927 -39198
rect 16963 -38902 17587 -38898
rect 16963 -39198 16967 -38902
rect 16967 -39198 17583 -38902
rect 17583 -39198 17587 -38902
rect 16963 -39202 17587 -39198
rect 17623 -38902 17927 -38898
rect 17623 -39198 17627 -38902
rect 17627 -39198 17923 -38902
rect 17923 -39198 17927 -38902
rect 17623 -39202 17927 -39198
rect 17963 -38902 18587 -38898
rect 17963 -39198 17967 -38902
rect 17967 -39198 18583 -38902
rect 18583 -39198 18587 -38902
rect 17963 -39202 18587 -39198
rect 18623 -38902 18927 -38898
rect 18623 -39198 18627 -38902
rect 18627 -39198 18923 -38902
rect 18923 -39198 18927 -38902
rect 18623 -39202 18927 -39198
rect 18963 -38902 19587 -38898
rect 18963 -39198 18967 -38902
rect 18967 -39198 19583 -38902
rect 19583 -39198 19587 -38902
rect 18963 -39202 19587 -39198
rect 19623 -38902 19927 -38898
rect 19623 -39198 19627 -38902
rect 19627 -39198 19923 -38902
rect 19923 -39198 19927 -38902
rect 19623 -39202 19927 -39198
rect 19963 -38902 20587 -38898
rect 19963 -39198 19967 -38902
rect 19967 -39198 20583 -38902
rect 20583 -39198 20587 -38902
rect 19963 -39202 20587 -39198
rect 20623 -38902 20927 -38898
rect 20623 -39198 20627 -38902
rect 20627 -39198 20923 -38902
rect 20923 -39198 20927 -38902
rect 20623 -39202 20927 -39198
rect 20963 -38902 21587 -38898
rect 20963 -39198 20967 -38902
rect 20967 -39198 21583 -38902
rect 21583 -39198 21587 -38902
rect 20963 -39202 21587 -39198
rect 21623 -38902 21927 -38898
rect 21623 -39198 21627 -38902
rect 21627 -39198 21923 -38902
rect 21923 -39198 21927 -38902
rect 21623 -39202 21927 -39198
rect 21963 -38902 22587 -38898
rect 21963 -39198 21967 -38902
rect 21967 -39198 22583 -38902
rect 22583 -39198 22587 -38902
rect 21963 -39202 22587 -39198
rect 22623 -38902 22927 -38898
rect 22623 -39198 22627 -38902
rect 22627 -39198 22923 -38902
rect 22923 -39198 22927 -38902
rect 22623 -39202 22927 -39198
rect 22963 -38902 23587 -38898
rect 22963 -39198 22967 -38902
rect 22967 -39198 23583 -38902
rect 23583 -39198 23587 -38902
rect 22963 -39202 23587 -39198
rect 23623 -38902 23927 -38898
rect 23623 -39198 23627 -38902
rect 23627 -39198 23923 -38902
rect 23923 -39198 23927 -38902
rect 23623 -39202 23927 -39198
rect 23963 -38902 24587 -38898
rect 23963 -39198 23967 -38902
rect 23967 -39198 24583 -38902
rect 24583 -39198 24587 -38902
rect 23963 -39202 24587 -39198
rect 24623 -38902 24927 -38898
rect 24623 -39198 24627 -38902
rect 24627 -39198 24923 -38902
rect 24923 -39198 24927 -38902
rect 24623 -39202 24927 -39198
rect 24963 -38902 25587 -38898
rect 24963 -39198 24967 -38902
rect 24967 -39198 25583 -38902
rect 25583 -39198 25587 -38902
rect 24963 -39202 25587 -39198
rect 25623 -38902 25927 -38898
rect 25623 -39198 25627 -38902
rect 25627 -39198 25923 -38902
rect 25923 -39198 25927 -38902
rect 25623 -39202 25927 -39198
rect 25963 -38902 26587 -38898
rect 25963 -39198 25967 -38902
rect 25967 -39198 26583 -38902
rect 26583 -39198 26587 -38902
rect 25963 -39202 26587 -39198
rect 26623 -38902 26927 -38898
rect 26623 -39198 26627 -38902
rect 26627 -39198 26923 -38902
rect 26923 -39198 26927 -38902
rect 26623 -39202 26927 -39198
rect 26963 -38902 27587 -38898
rect 26963 -39198 26967 -38902
rect 26967 -39198 27583 -38902
rect 27583 -39198 27587 -38902
rect 26963 -39202 27587 -39198
rect 27623 -38902 27927 -38898
rect 27623 -39198 27627 -38902
rect 27627 -39198 27923 -38902
rect 27923 -39198 27927 -38902
rect 27623 -39202 27927 -39198
rect 27963 -38902 28587 -38898
rect 27963 -39198 27967 -38902
rect 27967 -39198 28583 -38902
rect 28583 -39198 28587 -38902
rect 27963 -39202 28587 -39198
rect 28623 -38902 28927 -38898
rect 28623 -39198 28627 -38902
rect 28627 -39198 28923 -38902
rect 28923 -39198 28927 -38902
rect 28623 -39202 28927 -39198
rect 28963 -38902 29587 -38898
rect 28963 -39198 28967 -38902
rect 28967 -39198 29583 -38902
rect 29583 -39198 29587 -38902
rect 28963 -39202 29587 -39198
rect 29623 -38902 29927 -38898
rect 29623 -39198 29627 -38902
rect 29627 -39198 29923 -38902
rect 29923 -39198 29927 -38902
rect 29623 -39202 29927 -39198
rect 29963 -38902 30587 -38898
rect 29963 -39198 29967 -38902
rect 29967 -39198 30583 -38902
rect 30583 -39198 30587 -38902
rect 29963 -39202 30587 -39198
rect 30623 -38902 30927 -38898
rect 30623 -39198 30627 -38902
rect 30627 -39198 30923 -38902
rect 30923 -39198 30927 -38902
rect 30623 -39202 30927 -39198
rect 30963 -38902 31587 -38898
rect 30963 -39198 30967 -38902
rect 30967 -39198 31583 -38902
rect 31583 -39198 31587 -38902
rect 30963 -39202 31587 -39198
rect 31623 -38902 31927 -38898
rect 31623 -39198 31627 -38902
rect 31627 -39198 31923 -38902
rect 31923 -39198 31927 -38902
rect 31623 -39202 31927 -39198
rect 31963 -38902 32587 -38898
rect 31963 -39198 31967 -38902
rect 31967 -39198 32583 -38902
rect 32583 -39198 32587 -38902
rect 31963 -39202 32587 -39198
rect 32623 -38902 32927 -38898
rect 32623 -39198 32627 -38902
rect 32627 -39198 32923 -38902
rect 32923 -39198 32927 -38902
rect 32623 -39202 32927 -39198
rect 32963 -38902 33587 -38898
rect 32963 -39198 32967 -38902
rect 32967 -39198 33583 -38902
rect 33583 -39198 33587 -38902
rect 32963 -39202 33587 -39198
rect 33623 -38902 33927 -38898
rect 33623 -39198 33627 -38902
rect 33627 -39198 33923 -38902
rect 33923 -39198 33927 -38902
rect 33623 -39202 33927 -39198
rect 33963 -38902 34267 -38898
rect 33963 -39198 33967 -38902
rect 33967 -39198 34263 -38902
rect 34263 -39198 34267 -38902
rect 33963 -39202 34267 -39198
rect 8623 -39242 8927 -39238
rect 8623 -39858 8627 -39242
rect 8627 -39858 8923 -39242
rect 8923 -39858 8927 -39242
rect 8623 -39862 8927 -39858
rect 9623 -39242 9927 -39238
rect 9623 -39858 9627 -39242
rect 9627 -39858 9923 -39242
rect 9923 -39858 9927 -39242
rect 9623 -39862 9927 -39858
rect 10623 -39242 10927 -39238
rect 10623 -39858 10627 -39242
rect 10627 -39858 10923 -39242
rect 10923 -39858 10927 -39242
rect 10623 -39862 10927 -39858
rect 11623 -39242 11927 -39238
rect 11623 -39858 11627 -39242
rect 11627 -39858 11923 -39242
rect 11923 -39858 11927 -39242
rect 11623 -39862 11927 -39858
rect 12623 -39242 12927 -39238
rect 12623 -39858 12627 -39242
rect 12627 -39858 12923 -39242
rect 12923 -39858 12927 -39242
rect 12623 -39862 12927 -39858
rect 13623 -39242 13927 -39238
rect 13623 -39858 13627 -39242
rect 13627 -39858 13923 -39242
rect 13923 -39858 13927 -39242
rect 13623 -39862 13927 -39858
rect 14623 -39242 14927 -39238
rect 14623 -39858 14627 -39242
rect 14627 -39858 14923 -39242
rect 14923 -39858 14927 -39242
rect 14623 -39862 14927 -39858
rect 15623 -39242 15927 -39238
rect 15623 -39858 15627 -39242
rect 15627 -39858 15923 -39242
rect 15923 -39858 15927 -39242
rect 15623 -39862 15927 -39858
rect 16623 -39242 16927 -39238
rect 16623 -39858 16627 -39242
rect 16627 -39858 16923 -39242
rect 16923 -39858 16927 -39242
rect 16623 -39862 16927 -39858
rect 17623 -39242 17927 -39238
rect 17623 -39858 17627 -39242
rect 17627 -39858 17923 -39242
rect 17923 -39858 17927 -39242
rect 17623 -39862 17927 -39858
rect 18623 -39242 18927 -39238
rect 18623 -39858 18627 -39242
rect 18627 -39858 18923 -39242
rect 18923 -39858 18927 -39242
rect 18623 -39862 18927 -39858
rect 19623 -39242 19927 -39238
rect 19623 -39858 19627 -39242
rect 19627 -39858 19923 -39242
rect 19923 -39858 19927 -39242
rect 19623 -39862 19927 -39858
rect 20623 -39242 20927 -39238
rect 20623 -39858 20627 -39242
rect 20627 -39858 20923 -39242
rect 20923 -39858 20927 -39242
rect 20623 -39862 20927 -39858
rect 21623 -39242 21927 -39238
rect 21623 -39858 21627 -39242
rect 21627 -39858 21923 -39242
rect 21923 -39858 21927 -39242
rect 21623 -39862 21927 -39858
rect 22623 -39242 22927 -39238
rect 22623 -39858 22627 -39242
rect 22627 -39858 22923 -39242
rect 22923 -39858 22927 -39242
rect 22623 -39862 22927 -39858
rect 23623 -39242 23927 -39238
rect 23623 -39858 23627 -39242
rect 23627 -39858 23923 -39242
rect 23923 -39858 23927 -39242
rect 23623 -39862 23927 -39858
rect 24623 -39242 24927 -39238
rect 24623 -39858 24627 -39242
rect 24627 -39858 24923 -39242
rect 24923 -39858 24927 -39242
rect 24623 -39862 24927 -39858
rect 25623 -39242 25927 -39238
rect 25623 -39858 25627 -39242
rect 25627 -39858 25923 -39242
rect 25923 -39858 25927 -39242
rect 25623 -39862 25927 -39858
rect 26623 -39242 26927 -39238
rect 26623 -39858 26627 -39242
rect 26627 -39858 26923 -39242
rect 26923 -39858 26927 -39242
rect 26623 -39862 26927 -39858
rect 27623 -39242 27927 -39238
rect 27623 -39858 27627 -39242
rect 27627 -39858 27923 -39242
rect 27923 -39858 27927 -39242
rect 27623 -39862 27927 -39858
rect 28623 -39242 28927 -39238
rect 28623 -39858 28627 -39242
rect 28627 -39858 28923 -39242
rect 28923 -39858 28927 -39242
rect 28623 -39862 28927 -39858
rect 29623 -39242 29927 -39238
rect 29623 -39858 29627 -39242
rect 29627 -39858 29923 -39242
rect 29923 -39858 29927 -39242
rect 29623 -39862 29927 -39858
rect 30623 -39242 30927 -39238
rect 30623 -39858 30627 -39242
rect 30627 -39858 30923 -39242
rect 30923 -39858 30927 -39242
rect 30623 -39862 30927 -39858
rect 31623 -39242 31927 -39238
rect 31623 -39858 31627 -39242
rect 31627 -39858 31923 -39242
rect 31923 -39858 31927 -39242
rect 31623 -39862 31927 -39858
rect 32623 -39242 32927 -39238
rect 32623 -39858 32627 -39242
rect 32627 -39858 32923 -39242
rect 32923 -39858 32927 -39242
rect 32623 -39862 32927 -39858
rect 33623 -39242 33927 -39238
rect 33623 -39858 33627 -39242
rect 33627 -39858 33923 -39242
rect 33923 -39858 33927 -39242
rect 33623 -39862 33927 -39858
rect 8283 -39902 8587 -39898
rect 8283 -40198 8287 -39902
rect 8287 -40198 8583 -39902
rect 8583 -40198 8587 -39902
rect 8283 -40202 8587 -40198
rect 8623 -39902 8927 -39898
rect 8623 -40198 8627 -39902
rect 8627 -40198 8923 -39902
rect 8923 -40198 8927 -39902
rect 8623 -40202 8927 -40198
rect 8963 -39902 9587 -39898
rect 8963 -40198 8967 -39902
rect 8967 -40198 9583 -39902
rect 9583 -40198 9587 -39902
rect 8963 -40202 9587 -40198
rect 9623 -39902 9927 -39898
rect 9623 -40198 9627 -39902
rect 9627 -40198 9923 -39902
rect 9923 -40198 9927 -39902
rect 9623 -40202 9927 -40198
rect 9963 -39902 10587 -39898
rect 9963 -40198 9967 -39902
rect 9967 -40198 10583 -39902
rect 10583 -40198 10587 -39902
rect 9963 -40202 10587 -40198
rect 10623 -39902 10927 -39898
rect 10623 -40198 10627 -39902
rect 10627 -40198 10923 -39902
rect 10923 -40198 10927 -39902
rect 10623 -40202 10927 -40198
rect 10963 -39902 11587 -39898
rect 10963 -40198 10967 -39902
rect 10967 -40198 11583 -39902
rect 11583 -40198 11587 -39902
rect 10963 -40202 11587 -40198
rect 11623 -39902 11927 -39898
rect 11623 -40198 11627 -39902
rect 11627 -40198 11923 -39902
rect 11923 -40198 11927 -39902
rect 11623 -40202 11927 -40198
rect 11963 -39902 12587 -39898
rect 11963 -40198 11967 -39902
rect 11967 -40198 12583 -39902
rect 12583 -40198 12587 -39902
rect 11963 -40202 12587 -40198
rect 12623 -39902 12927 -39898
rect 12623 -40198 12627 -39902
rect 12627 -40198 12923 -39902
rect 12923 -40198 12927 -39902
rect 12623 -40202 12927 -40198
rect 12963 -39902 13587 -39898
rect 12963 -40198 12967 -39902
rect 12967 -40198 13583 -39902
rect 13583 -40198 13587 -39902
rect 12963 -40202 13587 -40198
rect 13623 -39902 13927 -39898
rect 13623 -40198 13627 -39902
rect 13627 -40198 13923 -39902
rect 13923 -40198 13927 -39902
rect 13623 -40202 13927 -40198
rect 13963 -39902 14587 -39898
rect 13963 -40198 13967 -39902
rect 13967 -40198 14583 -39902
rect 14583 -40198 14587 -39902
rect 13963 -40202 14587 -40198
rect 14623 -39902 14927 -39898
rect 14623 -40198 14627 -39902
rect 14627 -40198 14923 -39902
rect 14923 -40198 14927 -39902
rect 14623 -40202 14927 -40198
rect 14963 -39902 15587 -39898
rect 14963 -40198 14967 -39902
rect 14967 -40198 15583 -39902
rect 15583 -40198 15587 -39902
rect 14963 -40202 15587 -40198
rect 15623 -39902 15927 -39898
rect 15623 -40198 15627 -39902
rect 15627 -40198 15923 -39902
rect 15923 -40198 15927 -39902
rect 15623 -40202 15927 -40198
rect 15963 -39902 16587 -39898
rect 15963 -40198 15967 -39902
rect 15967 -40198 16583 -39902
rect 16583 -40198 16587 -39902
rect 15963 -40202 16587 -40198
rect 16623 -39902 16927 -39898
rect 16623 -40198 16627 -39902
rect 16627 -40198 16923 -39902
rect 16923 -40198 16927 -39902
rect 16623 -40202 16927 -40198
rect 16963 -39902 17587 -39898
rect 16963 -40198 16967 -39902
rect 16967 -40198 17583 -39902
rect 17583 -40198 17587 -39902
rect 16963 -40202 17587 -40198
rect 17623 -39902 17927 -39898
rect 17623 -40198 17627 -39902
rect 17627 -40198 17923 -39902
rect 17923 -40198 17927 -39902
rect 17623 -40202 17927 -40198
rect 17963 -39902 18587 -39898
rect 17963 -40198 17967 -39902
rect 17967 -40198 18583 -39902
rect 18583 -40198 18587 -39902
rect 17963 -40202 18587 -40198
rect 18623 -39902 18927 -39898
rect 18623 -40198 18627 -39902
rect 18627 -40198 18923 -39902
rect 18923 -40198 18927 -39902
rect 18623 -40202 18927 -40198
rect 18963 -39902 19587 -39898
rect 18963 -40198 18967 -39902
rect 18967 -40198 19583 -39902
rect 19583 -40198 19587 -39902
rect 18963 -40202 19587 -40198
rect 19623 -39902 19927 -39898
rect 19623 -40198 19627 -39902
rect 19627 -40198 19923 -39902
rect 19923 -40198 19927 -39902
rect 19623 -40202 19927 -40198
rect 19963 -39902 20587 -39898
rect 19963 -40198 19967 -39902
rect 19967 -40198 20583 -39902
rect 20583 -40198 20587 -39902
rect 19963 -40202 20587 -40198
rect 20623 -39902 20927 -39898
rect 20623 -40198 20627 -39902
rect 20627 -40198 20923 -39902
rect 20923 -40198 20927 -39902
rect 20623 -40202 20927 -40198
rect 20963 -39902 21587 -39898
rect 20963 -40198 20967 -39902
rect 20967 -40198 21583 -39902
rect 21583 -40198 21587 -39902
rect 20963 -40202 21587 -40198
rect 21623 -39902 21927 -39898
rect 21623 -40198 21627 -39902
rect 21627 -40198 21923 -39902
rect 21923 -40198 21927 -39902
rect 21623 -40202 21927 -40198
rect 21963 -39902 22587 -39898
rect 21963 -40198 21967 -39902
rect 21967 -40198 22583 -39902
rect 22583 -40198 22587 -39902
rect 21963 -40202 22587 -40198
rect 22623 -39902 22927 -39898
rect 22623 -40198 22627 -39902
rect 22627 -40198 22923 -39902
rect 22923 -40198 22927 -39902
rect 22623 -40202 22927 -40198
rect 22963 -39902 23587 -39898
rect 22963 -40198 22967 -39902
rect 22967 -40198 23583 -39902
rect 23583 -40198 23587 -39902
rect 22963 -40202 23587 -40198
rect 23623 -39902 23927 -39898
rect 23623 -40198 23627 -39902
rect 23627 -40198 23923 -39902
rect 23923 -40198 23927 -39902
rect 23623 -40202 23927 -40198
rect 23963 -39902 24587 -39898
rect 23963 -40198 23967 -39902
rect 23967 -40198 24583 -39902
rect 24583 -40198 24587 -39902
rect 23963 -40202 24587 -40198
rect 24623 -39902 24927 -39898
rect 24623 -40198 24627 -39902
rect 24627 -40198 24923 -39902
rect 24923 -40198 24927 -39902
rect 24623 -40202 24927 -40198
rect 24963 -39902 25587 -39898
rect 24963 -40198 24967 -39902
rect 24967 -40198 25583 -39902
rect 25583 -40198 25587 -39902
rect 24963 -40202 25587 -40198
rect 25623 -39902 25927 -39898
rect 25623 -40198 25627 -39902
rect 25627 -40198 25923 -39902
rect 25923 -40198 25927 -39902
rect 25623 -40202 25927 -40198
rect 25963 -39902 26587 -39898
rect 25963 -40198 25967 -39902
rect 25967 -40198 26583 -39902
rect 26583 -40198 26587 -39902
rect 25963 -40202 26587 -40198
rect 26623 -39902 26927 -39898
rect 26623 -40198 26627 -39902
rect 26627 -40198 26923 -39902
rect 26923 -40198 26927 -39902
rect 26623 -40202 26927 -40198
rect 26963 -39902 27587 -39898
rect 26963 -40198 26967 -39902
rect 26967 -40198 27583 -39902
rect 27583 -40198 27587 -39902
rect 26963 -40202 27587 -40198
rect 27623 -39902 27927 -39898
rect 27623 -40198 27627 -39902
rect 27627 -40198 27923 -39902
rect 27923 -40198 27927 -39902
rect 27623 -40202 27927 -40198
rect 27963 -39902 28587 -39898
rect 27963 -40198 27967 -39902
rect 27967 -40198 28583 -39902
rect 28583 -40198 28587 -39902
rect 27963 -40202 28587 -40198
rect 28623 -39902 28927 -39898
rect 28623 -40198 28627 -39902
rect 28627 -40198 28923 -39902
rect 28923 -40198 28927 -39902
rect 28623 -40202 28927 -40198
rect 28963 -39902 29587 -39898
rect 28963 -40198 28967 -39902
rect 28967 -40198 29583 -39902
rect 29583 -40198 29587 -39902
rect 28963 -40202 29587 -40198
rect 29623 -39902 29927 -39898
rect 29623 -40198 29627 -39902
rect 29627 -40198 29923 -39902
rect 29923 -40198 29927 -39902
rect 29623 -40202 29927 -40198
rect 29963 -39902 30587 -39898
rect 29963 -40198 29967 -39902
rect 29967 -40198 30583 -39902
rect 30583 -40198 30587 -39902
rect 29963 -40202 30587 -40198
rect 30623 -39902 30927 -39898
rect 30623 -40198 30627 -39902
rect 30627 -40198 30923 -39902
rect 30923 -40198 30927 -39902
rect 30623 -40202 30927 -40198
rect 30963 -39902 31587 -39898
rect 30963 -40198 30967 -39902
rect 30967 -40198 31583 -39902
rect 31583 -40198 31587 -39902
rect 30963 -40202 31587 -40198
rect 31623 -39902 31927 -39898
rect 31623 -40198 31627 -39902
rect 31627 -40198 31923 -39902
rect 31923 -40198 31927 -39902
rect 31623 -40202 31927 -40198
rect 31963 -39902 32587 -39898
rect 31963 -40198 31967 -39902
rect 31967 -40198 32583 -39902
rect 32583 -40198 32587 -39902
rect 31963 -40202 32587 -40198
rect 32623 -39902 32927 -39898
rect 32623 -40198 32627 -39902
rect 32627 -40198 32923 -39902
rect 32923 -40198 32927 -39902
rect 32623 -40202 32927 -40198
rect 32963 -39902 33587 -39898
rect 32963 -40198 32967 -39902
rect 32967 -40198 33583 -39902
rect 33583 -40198 33587 -39902
rect 32963 -40202 33587 -40198
rect 33623 -39902 33927 -39898
rect 33623 -40198 33627 -39902
rect 33627 -40198 33923 -39902
rect 33923 -40198 33927 -39902
rect 33623 -40202 33927 -40198
rect 33963 -39902 34267 -39898
rect 33963 -40198 33967 -39902
rect 33967 -40198 34263 -39902
rect 34263 -40198 34267 -39902
rect 33963 -40202 34267 -40198
rect 8623 -40242 8927 -40238
rect 8623 -40858 8627 -40242
rect 8627 -40858 8923 -40242
rect 8923 -40858 8927 -40242
rect 8623 -40862 8927 -40858
rect 9623 -40242 9927 -40238
rect 9623 -40858 9627 -40242
rect 9627 -40858 9923 -40242
rect 9923 -40858 9927 -40242
rect 9623 -40862 9927 -40858
rect 10623 -40242 10927 -40238
rect 10623 -40858 10627 -40242
rect 10627 -40858 10923 -40242
rect 10923 -40858 10927 -40242
rect 10623 -40862 10927 -40858
rect 11623 -40242 11927 -40238
rect 11623 -40858 11627 -40242
rect 11627 -40858 11923 -40242
rect 11923 -40858 11927 -40242
rect 11623 -40862 11927 -40858
rect 12623 -40242 12927 -40238
rect 12623 -40858 12627 -40242
rect 12627 -40858 12923 -40242
rect 12923 -40858 12927 -40242
rect 12623 -40862 12927 -40858
rect 13623 -40242 13927 -40238
rect 13623 -40858 13627 -40242
rect 13627 -40858 13923 -40242
rect 13923 -40858 13927 -40242
rect 13623 -40862 13927 -40858
rect 14623 -40242 14927 -40238
rect 14623 -40858 14627 -40242
rect 14627 -40858 14923 -40242
rect 14923 -40858 14927 -40242
rect 14623 -40862 14927 -40858
rect 15623 -40242 15927 -40238
rect 15623 -40858 15627 -40242
rect 15627 -40858 15923 -40242
rect 15923 -40858 15927 -40242
rect 15623 -40862 15927 -40858
rect 16623 -40242 16927 -40238
rect 16623 -40858 16627 -40242
rect 16627 -40858 16923 -40242
rect 16923 -40858 16927 -40242
rect 16623 -40862 16927 -40858
rect 17623 -40242 17927 -40238
rect 17623 -40858 17627 -40242
rect 17627 -40858 17923 -40242
rect 17923 -40858 17927 -40242
rect 17623 -40862 17927 -40858
rect 18623 -40242 18927 -40238
rect 18623 -40858 18627 -40242
rect 18627 -40858 18923 -40242
rect 18923 -40858 18927 -40242
rect 18623 -40862 18927 -40858
rect 19623 -40242 19927 -40238
rect 19623 -40858 19627 -40242
rect 19627 -40858 19923 -40242
rect 19923 -40858 19927 -40242
rect 19623 -40862 19927 -40858
rect 20623 -40242 20927 -40238
rect 20623 -40858 20627 -40242
rect 20627 -40858 20923 -40242
rect 20923 -40858 20927 -40242
rect 20623 -40862 20927 -40858
rect 21623 -40242 21927 -40238
rect 21623 -40858 21627 -40242
rect 21627 -40858 21923 -40242
rect 21923 -40858 21927 -40242
rect 21623 -40862 21927 -40858
rect 22623 -40242 22927 -40238
rect 22623 -40858 22627 -40242
rect 22627 -40858 22923 -40242
rect 22923 -40858 22927 -40242
rect 22623 -40862 22927 -40858
rect 23623 -40242 23927 -40238
rect 23623 -40858 23627 -40242
rect 23627 -40858 23923 -40242
rect 23923 -40858 23927 -40242
rect 23623 -40862 23927 -40858
rect 24623 -40242 24927 -40238
rect 24623 -40858 24627 -40242
rect 24627 -40858 24923 -40242
rect 24923 -40858 24927 -40242
rect 24623 -40862 24927 -40858
rect 25623 -40242 25927 -40238
rect 25623 -40858 25627 -40242
rect 25627 -40858 25923 -40242
rect 25923 -40858 25927 -40242
rect 25623 -40862 25927 -40858
rect 26623 -40242 26927 -40238
rect 26623 -40858 26627 -40242
rect 26627 -40858 26923 -40242
rect 26923 -40858 26927 -40242
rect 26623 -40862 26927 -40858
rect 27623 -40242 27927 -40238
rect 27623 -40858 27627 -40242
rect 27627 -40858 27923 -40242
rect 27923 -40858 27927 -40242
rect 27623 -40862 27927 -40858
rect 28623 -40242 28927 -40238
rect 28623 -40858 28627 -40242
rect 28627 -40858 28923 -40242
rect 28923 -40858 28927 -40242
rect 28623 -40862 28927 -40858
rect 29623 -40242 29927 -40238
rect 29623 -40858 29627 -40242
rect 29627 -40858 29923 -40242
rect 29923 -40858 29927 -40242
rect 29623 -40862 29927 -40858
rect 30623 -40242 30927 -40238
rect 30623 -40858 30627 -40242
rect 30627 -40858 30923 -40242
rect 30923 -40858 30927 -40242
rect 30623 -40862 30927 -40858
rect 31623 -40242 31927 -40238
rect 31623 -40858 31627 -40242
rect 31627 -40858 31923 -40242
rect 31923 -40858 31927 -40242
rect 31623 -40862 31927 -40858
rect 32623 -40242 32927 -40238
rect 32623 -40858 32627 -40242
rect 32627 -40858 32923 -40242
rect 32923 -40858 32927 -40242
rect 32623 -40862 32927 -40858
rect 33623 -40242 33927 -40238
rect 33623 -40858 33627 -40242
rect 33627 -40858 33923 -40242
rect 33923 -40858 33927 -40242
rect 33623 -40862 33927 -40858
rect 8283 -40902 8587 -40898
rect 8283 -41198 8287 -40902
rect 8287 -41198 8583 -40902
rect 8583 -41198 8587 -40902
rect 8283 -41202 8587 -41198
rect 8623 -40902 8927 -40898
rect 8623 -41198 8627 -40902
rect 8627 -41198 8923 -40902
rect 8923 -41198 8927 -40902
rect 8623 -41202 8927 -41198
rect 8963 -40902 9587 -40898
rect 8963 -41198 8967 -40902
rect 8967 -41198 9583 -40902
rect 9583 -41198 9587 -40902
rect 8963 -41202 9587 -41198
rect 9623 -40902 9927 -40898
rect 9623 -41198 9627 -40902
rect 9627 -41198 9923 -40902
rect 9923 -41198 9927 -40902
rect 9623 -41202 9927 -41198
rect 9963 -40902 10587 -40898
rect 9963 -41198 9967 -40902
rect 9967 -41198 10583 -40902
rect 10583 -41198 10587 -40902
rect 9963 -41202 10587 -41198
rect 10623 -40902 10927 -40898
rect 10623 -41198 10627 -40902
rect 10627 -41198 10923 -40902
rect 10923 -41198 10927 -40902
rect 10623 -41202 10927 -41198
rect 10963 -40902 11587 -40898
rect 10963 -41198 10967 -40902
rect 10967 -41198 11583 -40902
rect 11583 -41198 11587 -40902
rect 10963 -41202 11587 -41198
rect 11623 -40902 11927 -40898
rect 11623 -41198 11627 -40902
rect 11627 -41198 11923 -40902
rect 11923 -41198 11927 -40902
rect 11623 -41202 11927 -41198
rect 11963 -40902 12587 -40898
rect 11963 -41198 11967 -40902
rect 11967 -41198 12583 -40902
rect 12583 -41198 12587 -40902
rect 11963 -41202 12587 -41198
rect 12623 -40902 12927 -40898
rect 12623 -41198 12627 -40902
rect 12627 -41198 12923 -40902
rect 12923 -41198 12927 -40902
rect 12623 -41202 12927 -41198
rect 12963 -40902 13587 -40898
rect 12963 -41198 12967 -40902
rect 12967 -41198 13583 -40902
rect 13583 -41198 13587 -40902
rect 12963 -41202 13587 -41198
rect 13623 -40902 13927 -40898
rect 13623 -41198 13627 -40902
rect 13627 -41198 13923 -40902
rect 13923 -41198 13927 -40902
rect 13623 -41202 13927 -41198
rect 13963 -40902 14587 -40898
rect 13963 -41198 13967 -40902
rect 13967 -41198 14583 -40902
rect 14583 -41198 14587 -40902
rect 13963 -41202 14587 -41198
rect 14623 -40902 14927 -40898
rect 14623 -41198 14627 -40902
rect 14627 -41198 14923 -40902
rect 14923 -41198 14927 -40902
rect 14623 -41202 14927 -41198
rect 14963 -40902 15587 -40898
rect 14963 -41198 14967 -40902
rect 14967 -41198 15583 -40902
rect 15583 -41198 15587 -40902
rect 14963 -41202 15587 -41198
rect 15623 -40902 15927 -40898
rect 15623 -41198 15627 -40902
rect 15627 -41198 15923 -40902
rect 15923 -41198 15927 -40902
rect 15623 -41202 15927 -41198
rect 15963 -40902 16587 -40898
rect 15963 -41198 15967 -40902
rect 15967 -41198 16583 -40902
rect 16583 -41198 16587 -40902
rect 15963 -41202 16587 -41198
rect 16623 -40902 16927 -40898
rect 16623 -41198 16627 -40902
rect 16627 -41198 16923 -40902
rect 16923 -41198 16927 -40902
rect 16623 -41202 16927 -41198
rect 16963 -40902 17587 -40898
rect 16963 -41198 16967 -40902
rect 16967 -41198 17583 -40902
rect 17583 -41198 17587 -40902
rect 16963 -41202 17587 -41198
rect 17623 -40902 17927 -40898
rect 17623 -41198 17627 -40902
rect 17627 -41198 17923 -40902
rect 17923 -41198 17927 -40902
rect 17623 -41202 17927 -41198
rect 17963 -40902 18587 -40898
rect 17963 -41198 17967 -40902
rect 17967 -41198 18583 -40902
rect 18583 -41198 18587 -40902
rect 17963 -41202 18587 -41198
rect 18623 -40902 18927 -40898
rect 18623 -41198 18627 -40902
rect 18627 -41198 18923 -40902
rect 18923 -41198 18927 -40902
rect 18623 -41202 18927 -41198
rect 18963 -40902 19587 -40898
rect 18963 -41198 18967 -40902
rect 18967 -41198 19583 -40902
rect 19583 -41198 19587 -40902
rect 18963 -41202 19587 -41198
rect 19623 -40902 19927 -40898
rect 19623 -41198 19627 -40902
rect 19627 -41198 19923 -40902
rect 19923 -41198 19927 -40902
rect 19623 -41202 19927 -41198
rect 19963 -40902 20587 -40898
rect 19963 -41198 19967 -40902
rect 19967 -41198 20583 -40902
rect 20583 -41198 20587 -40902
rect 19963 -41202 20587 -41198
rect 20623 -40902 20927 -40898
rect 20623 -41198 20627 -40902
rect 20627 -41198 20923 -40902
rect 20923 -41198 20927 -40902
rect 20623 -41202 20927 -41198
rect 20963 -40902 21587 -40898
rect 20963 -41198 20967 -40902
rect 20967 -41198 21583 -40902
rect 21583 -41198 21587 -40902
rect 20963 -41202 21587 -41198
rect 21623 -40902 21927 -40898
rect 21623 -41198 21627 -40902
rect 21627 -41198 21923 -40902
rect 21923 -41198 21927 -40902
rect 21623 -41202 21927 -41198
rect 21963 -40902 22587 -40898
rect 21963 -41198 21967 -40902
rect 21967 -41198 22583 -40902
rect 22583 -41198 22587 -40902
rect 21963 -41202 22587 -41198
rect 22623 -40902 22927 -40898
rect 22623 -41198 22627 -40902
rect 22627 -41198 22923 -40902
rect 22923 -41198 22927 -40902
rect 22623 -41202 22927 -41198
rect 22963 -40902 23587 -40898
rect 22963 -41198 22967 -40902
rect 22967 -41198 23583 -40902
rect 23583 -41198 23587 -40902
rect 22963 -41202 23587 -41198
rect 23623 -40902 23927 -40898
rect 23623 -41198 23627 -40902
rect 23627 -41198 23923 -40902
rect 23923 -41198 23927 -40902
rect 23623 -41202 23927 -41198
rect 23963 -40902 24587 -40898
rect 23963 -41198 23967 -40902
rect 23967 -41198 24583 -40902
rect 24583 -41198 24587 -40902
rect 23963 -41202 24587 -41198
rect 24623 -40902 24927 -40898
rect 24623 -41198 24627 -40902
rect 24627 -41198 24923 -40902
rect 24923 -41198 24927 -40902
rect 24623 -41202 24927 -41198
rect 24963 -40902 25587 -40898
rect 24963 -41198 24967 -40902
rect 24967 -41198 25583 -40902
rect 25583 -41198 25587 -40902
rect 24963 -41202 25587 -41198
rect 25623 -40902 25927 -40898
rect 25623 -41198 25627 -40902
rect 25627 -41198 25923 -40902
rect 25923 -41198 25927 -40902
rect 25623 -41202 25927 -41198
rect 25963 -40902 26587 -40898
rect 25963 -41198 25967 -40902
rect 25967 -41198 26583 -40902
rect 26583 -41198 26587 -40902
rect 25963 -41202 26587 -41198
rect 26623 -40902 26927 -40898
rect 26623 -41198 26627 -40902
rect 26627 -41198 26923 -40902
rect 26923 -41198 26927 -40902
rect 26623 -41202 26927 -41198
rect 26963 -40902 27587 -40898
rect 26963 -41198 26967 -40902
rect 26967 -41198 27583 -40902
rect 27583 -41198 27587 -40902
rect 26963 -41202 27587 -41198
rect 27623 -40902 27927 -40898
rect 27623 -41198 27627 -40902
rect 27627 -41198 27923 -40902
rect 27923 -41198 27927 -40902
rect 27623 -41202 27927 -41198
rect 27963 -40902 28587 -40898
rect 27963 -41198 27967 -40902
rect 27967 -41198 28583 -40902
rect 28583 -41198 28587 -40902
rect 27963 -41202 28587 -41198
rect 28623 -40902 28927 -40898
rect 28623 -41198 28627 -40902
rect 28627 -41198 28923 -40902
rect 28923 -41198 28927 -40902
rect 28623 -41202 28927 -41198
rect 28963 -40902 29587 -40898
rect 28963 -41198 28967 -40902
rect 28967 -41198 29583 -40902
rect 29583 -41198 29587 -40902
rect 28963 -41202 29587 -41198
rect 29623 -40902 29927 -40898
rect 29623 -41198 29627 -40902
rect 29627 -41198 29923 -40902
rect 29923 -41198 29927 -40902
rect 29623 -41202 29927 -41198
rect 29963 -40902 30587 -40898
rect 29963 -41198 29967 -40902
rect 29967 -41198 30583 -40902
rect 30583 -41198 30587 -40902
rect 29963 -41202 30587 -41198
rect 30623 -40902 30927 -40898
rect 30623 -41198 30627 -40902
rect 30627 -41198 30923 -40902
rect 30923 -41198 30927 -40902
rect 30623 -41202 30927 -41198
rect 30963 -40902 31587 -40898
rect 30963 -41198 30967 -40902
rect 30967 -41198 31583 -40902
rect 31583 -41198 31587 -40902
rect 30963 -41202 31587 -41198
rect 31623 -40902 31927 -40898
rect 31623 -41198 31627 -40902
rect 31627 -41198 31923 -40902
rect 31923 -41198 31927 -40902
rect 31623 -41202 31927 -41198
rect 31963 -40902 32587 -40898
rect 31963 -41198 31967 -40902
rect 31967 -41198 32583 -40902
rect 32583 -41198 32587 -40902
rect 31963 -41202 32587 -41198
rect 32623 -40902 32927 -40898
rect 32623 -41198 32627 -40902
rect 32627 -41198 32923 -40902
rect 32923 -41198 32927 -40902
rect 32623 -41202 32927 -41198
rect 32963 -40902 33587 -40898
rect 32963 -41198 32967 -40902
rect 32967 -41198 33583 -40902
rect 33583 -41198 33587 -40902
rect 32963 -41202 33587 -41198
rect 33623 -40902 33927 -40898
rect 33623 -41198 33627 -40902
rect 33627 -41198 33923 -40902
rect 33923 -41198 33927 -40902
rect 33623 -41202 33927 -41198
rect 33963 -40902 34267 -40898
rect 33963 -41198 33967 -40902
rect 33967 -41198 34263 -40902
rect 34263 -41198 34267 -40902
rect 33963 -41202 34267 -41198
rect 8623 -41242 8927 -41238
rect 8623 -41858 8627 -41242
rect 8627 -41858 8923 -41242
rect 8923 -41858 8927 -41242
rect 8623 -41862 8927 -41858
rect 9623 -41242 9927 -41238
rect 9623 -41858 9627 -41242
rect 9627 -41858 9923 -41242
rect 9923 -41858 9927 -41242
rect 9623 -41862 9927 -41858
rect 10623 -41242 10927 -41238
rect 10623 -41858 10627 -41242
rect 10627 -41858 10923 -41242
rect 10923 -41858 10927 -41242
rect 10623 -41862 10927 -41858
rect 11623 -41242 11927 -41238
rect 11623 -41858 11627 -41242
rect 11627 -41858 11923 -41242
rect 11923 -41858 11927 -41242
rect 11623 -41862 11927 -41858
rect 12623 -41242 12927 -41238
rect 12623 -41858 12627 -41242
rect 12627 -41858 12923 -41242
rect 12923 -41858 12927 -41242
rect 12623 -41862 12927 -41858
rect 13623 -41242 13927 -41238
rect 13623 -41858 13627 -41242
rect 13627 -41858 13923 -41242
rect 13923 -41858 13927 -41242
rect 13623 -41862 13927 -41858
rect 14623 -41242 14927 -41238
rect 14623 -41858 14627 -41242
rect 14627 -41858 14923 -41242
rect 14923 -41858 14927 -41242
rect 14623 -41862 14927 -41858
rect 15623 -41242 15927 -41238
rect 15623 -41858 15627 -41242
rect 15627 -41858 15923 -41242
rect 15923 -41858 15927 -41242
rect 15623 -41862 15927 -41858
rect 16623 -41242 16927 -41238
rect 16623 -41858 16627 -41242
rect 16627 -41858 16923 -41242
rect 16923 -41858 16927 -41242
rect 16623 -41862 16927 -41858
rect 17623 -41242 17927 -41238
rect 17623 -41858 17627 -41242
rect 17627 -41858 17923 -41242
rect 17923 -41858 17927 -41242
rect 17623 -41862 17927 -41858
rect 18623 -41242 18927 -41238
rect 18623 -41858 18627 -41242
rect 18627 -41858 18923 -41242
rect 18923 -41858 18927 -41242
rect 18623 -41862 18927 -41858
rect 19623 -41242 19927 -41238
rect 19623 -41858 19627 -41242
rect 19627 -41858 19923 -41242
rect 19923 -41858 19927 -41242
rect 19623 -41862 19927 -41858
rect 20623 -41242 20927 -41238
rect 20623 -41858 20627 -41242
rect 20627 -41858 20923 -41242
rect 20923 -41858 20927 -41242
rect 20623 -41862 20927 -41858
rect 21623 -41242 21927 -41238
rect 21623 -41858 21627 -41242
rect 21627 -41858 21923 -41242
rect 21923 -41858 21927 -41242
rect 21623 -41862 21927 -41858
rect 22623 -41242 22927 -41238
rect 22623 -41858 22627 -41242
rect 22627 -41858 22923 -41242
rect 22923 -41858 22927 -41242
rect 22623 -41862 22927 -41858
rect 23623 -41242 23927 -41238
rect 23623 -41858 23627 -41242
rect 23627 -41858 23923 -41242
rect 23923 -41858 23927 -41242
rect 23623 -41862 23927 -41858
rect 24623 -41242 24927 -41238
rect 24623 -41858 24627 -41242
rect 24627 -41858 24923 -41242
rect 24923 -41858 24927 -41242
rect 24623 -41862 24927 -41858
rect 25623 -41242 25927 -41238
rect 25623 -41858 25627 -41242
rect 25627 -41858 25923 -41242
rect 25923 -41858 25927 -41242
rect 25623 -41862 25927 -41858
rect 26623 -41242 26927 -41238
rect 26623 -41858 26627 -41242
rect 26627 -41858 26923 -41242
rect 26923 -41858 26927 -41242
rect 26623 -41862 26927 -41858
rect 27623 -41242 27927 -41238
rect 27623 -41858 27627 -41242
rect 27627 -41858 27923 -41242
rect 27923 -41858 27927 -41242
rect 27623 -41862 27927 -41858
rect 28623 -41242 28927 -41238
rect 28623 -41858 28627 -41242
rect 28627 -41858 28923 -41242
rect 28923 -41858 28927 -41242
rect 28623 -41862 28927 -41858
rect 29623 -41242 29927 -41238
rect 29623 -41858 29627 -41242
rect 29627 -41858 29923 -41242
rect 29923 -41858 29927 -41242
rect 29623 -41862 29927 -41858
rect 30623 -41242 30927 -41238
rect 30623 -41858 30627 -41242
rect 30627 -41858 30923 -41242
rect 30923 -41858 30927 -41242
rect 30623 -41862 30927 -41858
rect 31623 -41242 31927 -41238
rect 31623 -41858 31627 -41242
rect 31627 -41858 31923 -41242
rect 31923 -41858 31927 -41242
rect 31623 -41862 31927 -41858
rect 32623 -41242 32927 -41238
rect 32623 -41858 32627 -41242
rect 32627 -41858 32923 -41242
rect 32923 -41858 32927 -41242
rect 32623 -41862 32927 -41858
rect 33623 -41242 33927 -41238
rect 33623 -41858 33627 -41242
rect 33627 -41858 33923 -41242
rect 33923 -41858 33927 -41242
rect 33623 -41862 33927 -41858
rect 8283 -41902 8587 -41898
rect 8283 -42198 8287 -41902
rect 8287 -42198 8583 -41902
rect 8583 -42198 8587 -41902
rect 8283 -42202 8587 -42198
rect 8623 -41902 8927 -41898
rect 8623 -42198 8627 -41902
rect 8627 -42198 8923 -41902
rect 8923 -42198 8927 -41902
rect 8623 -42202 8927 -42198
rect 8963 -41902 9587 -41898
rect 8963 -42198 8967 -41902
rect 8967 -42198 9583 -41902
rect 9583 -42198 9587 -41902
rect 8963 -42202 9587 -42198
rect 9623 -41902 9927 -41898
rect 9623 -42198 9627 -41902
rect 9627 -42198 9923 -41902
rect 9923 -42198 9927 -41902
rect 9623 -42202 9927 -42198
rect 9963 -41902 10587 -41898
rect 9963 -42198 9967 -41902
rect 9967 -42198 10583 -41902
rect 10583 -42198 10587 -41902
rect 9963 -42202 10587 -42198
rect 10623 -41902 10927 -41898
rect 10623 -42198 10627 -41902
rect 10627 -42198 10923 -41902
rect 10923 -42198 10927 -41902
rect 10623 -42202 10927 -42198
rect 10963 -41902 11587 -41898
rect 10963 -42198 10967 -41902
rect 10967 -42198 11583 -41902
rect 11583 -42198 11587 -41902
rect 10963 -42202 11587 -42198
rect 11623 -41902 11927 -41898
rect 11623 -42198 11627 -41902
rect 11627 -42198 11923 -41902
rect 11923 -42198 11927 -41902
rect 11623 -42202 11927 -42198
rect 11963 -41902 12587 -41898
rect 11963 -42198 11967 -41902
rect 11967 -42198 12583 -41902
rect 12583 -42198 12587 -41902
rect 11963 -42202 12587 -42198
rect 12623 -41902 12927 -41898
rect 12623 -42198 12627 -41902
rect 12627 -42198 12923 -41902
rect 12923 -42198 12927 -41902
rect 12623 -42202 12927 -42198
rect 12963 -41902 13587 -41898
rect 12963 -42198 12967 -41902
rect 12967 -42198 13583 -41902
rect 13583 -42198 13587 -41902
rect 12963 -42202 13587 -42198
rect 13623 -41902 13927 -41898
rect 13623 -42198 13627 -41902
rect 13627 -42198 13923 -41902
rect 13923 -42198 13927 -41902
rect 13623 -42202 13927 -42198
rect 13963 -41902 14587 -41898
rect 13963 -42198 13967 -41902
rect 13967 -42198 14583 -41902
rect 14583 -42198 14587 -41902
rect 13963 -42202 14587 -42198
rect 14623 -41902 14927 -41898
rect 14623 -42198 14627 -41902
rect 14627 -42198 14923 -41902
rect 14923 -42198 14927 -41902
rect 14623 -42202 14927 -42198
rect 14963 -41902 15587 -41898
rect 14963 -42198 14967 -41902
rect 14967 -42198 15583 -41902
rect 15583 -42198 15587 -41902
rect 14963 -42202 15587 -42198
rect 15623 -41902 15927 -41898
rect 15623 -42198 15627 -41902
rect 15627 -42198 15923 -41902
rect 15923 -42198 15927 -41902
rect 15623 -42202 15927 -42198
rect 15963 -41902 16587 -41898
rect 15963 -42198 15967 -41902
rect 15967 -42198 16583 -41902
rect 16583 -42198 16587 -41902
rect 15963 -42202 16587 -42198
rect 16623 -41902 16927 -41898
rect 16623 -42198 16627 -41902
rect 16627 -42198 16923 -41902
rect 16923 -42198 16927 -41902
rect 16623 -42202 16927 -42198
rect 16963 -41902 17587 -41898
rect 16963 -42198 16967 -41902
rect 16967 -42198 17583 -41902
rect 17583 -42198 17587 -41902
rect 16963 -42202 17587 -42198
rect 17623 -41902 17927 -41898
rect 17623 -42198 17627 -41902
rect 17627 -42198 17923 -41902
rect 17923 -42198 17927 -41902
rect 17623 -42202 17927 -42198
rect 17963 -41902 18587 -41898
rect 17963 -42198 17967 -41902
rect 17967 -42198 18583 -41902
rect 18583 -42198 18587 -41902
rect 17963 -42202 18587 -42198
rect 18623 -41902 18927 -41898
rect 18623 -42198 18627 -41902
rect 18627 -42198 18923 -41902
rect 18923 -42198 18927 -41902
rect 18623 -42202 18927 -42198
rect 18963 -41902 19587 -41898
rect 18963 -42198 18967 -41902
rect 18967 -42198 19583 -41902
rect 19583 -42198 19587 -41902
rect 18963 -42202 19587 -42198
rect 19623 -41902 19927 -41898
rect 19623 -42198 19627 -41902
rect 19627 -42198 19923 -41902
rect 19923 -42198 19927 -41902
rect 19623 -42202 19927 -42198
rect 19963 -41902 20587 -41898
rect 19963 -42198 19967 -41902
rect 19967 -42198 20583 -41902
rect 20583 -42198 20587 -41902
rect 19963 -42202 20587 -42198
rect 20623 -41902 20927 -41898
rect 20623 -42198 20627 -41902
rect 20627 -42198 20923 -41902
rect 20923 -42198 20927 -41902
rect 20623 -42202 20927 -42198
rect 20963 -41902 21587 -41898
rect 20963 -42198 20967 -41902
rect 20967 -42198 21583 -41902
rect 21583 -42198 21587 -41902
rect 20963 -42202 21587 -42198
rect 21623 -41902 21927 -41898
rect 21623 -42198 21627 -41902
rect 21627 -42198 21923 -41902
rect 21923 -42198 21927 -41902
rect 21623 -42202 21927 -42198
rect 21963 -41902 22587 -41898
rect 21963 -42198 21967 -41902
rect 21967 -42198 22583 -41902
rect 22583 -42198 22587 -41902
rect 21963 -42202 22587 -42198
rect 22623 -41902 22927 -41898
rect 22623 -42198 22627 -41902
rect 22627 -42198 22923 -41902
rect 22923 -42198 22927 -41902
rect 22623 -42202 22927 -42198
rect 22963 -41902 23587 -41898
rect 22963 -42198 22967 -41902
rect 22967 -42198 23583 -41902
rect 23583 -42198 23587 -41902
rect 22963 -42202 23587 -42198
rect 23623 -41902 23927 -41898
rect 23623 -42198 23627 -41902
rect 23627 -42198 23923 -41902
rect 23923 -42198 23927 -41902
rect 23623 -42202 23927 -42198
rect 23963 -41902 24587 -41898
rect 23963 -42198 23967 -41902
rect 23967 -42198 24583 -41902
rect 24583 -42198 24587 -41902
rect 23963 -42202 24587 -42198
rect 24623 -41902 24927 -41898
rect 24623 -42198 24627 -41902
rect 24627 -42198 24923 -41902
rect 24923 -42198 24927 -41902
rect 24623 -42202 24927 -42198
rect 24963 -41902 25587 -41898
rect 24963 -42198 24967 -41902
rect 24967 -42198 25583 -41902
rect 25583 -42198 25587 -41902
rect 24963 -42202 25587 -42198
rect 25623 -41902 25927 -41898
rect 25623 -42198 25627 -41902
rect 25627 -42198 25923 -41902
rect 25923 -42198 25927 -41902
rect 25623 -42202 25927 -42198
rect 25963 -41902 26587 -41898
rect 25963 -42198 25967 -41902
rect 25967 -42198 26583 -41902
rect 26583 -42198 26587 -41902
rect 25963 -42202 26587 -42198
rect 26623 -41902 26927 -41898
rect 26623 -42198 26627 -41902
rect 26627 -42198 26923 -41902
rect 26923 -42198 26927 -41902
rect 26623 -42202 26927 -42198
rect 26963 -41902 27587 -41898
rect 26963 -42198 26967 -41902
rect 26967 -42198 27583 -41902
rect 27583 -42198 27587 -41902
rect 26963 -42202 27587 -42198
rect 27623 -41902 27927 -41898
rect 27623 -42198 27627 -41902
rect 27627 -42198 27923 -41902
rect 27923 -42198 27927 -41902
rect 27623 -42202 27927 -42198
rect 27963 -41902 28587 -41898
rect 27963 -42198 27967 -41902
rect 27967 -42198 28583 -41902
rect 28583 -42198 28587 -41902
rect 27963 -42202 28587 -42198
rect 28623 -41902 28927 -41898
rect 28623 -42198 28627 -41902
rect 28627 -42198 28923 -41902
rect 28923 -42198 28927 -41902
rect 28623 -42202 28927 -42198
rect 28963 -41902 29587 -41898
rect 28963 -42198 28967 -41902
rect 28967 -42198 29583 -41902
rect 29583 -42198 29587 -41902
rect 28963 -42202 29587 -42198
rect 29623 -41902 29927 -41898
rect 29623 -42198 29627 -41902
rect 29627 -42198 29923 -41902
rect 29923 -42198 29927 -41902
rect 29623 -42202 29927 -42198
rect 29963 -41902 30587 -41898
rect 29963 -42198 29967 -41902
rect 29967 -42198 30583 -41902
rect 30583 -42198 30587 -41902
rect 29963 -42202 30587 -42198
rect 30623 -41902 30927 -41898
rect 30623 -42198 30627 -41902
rect 30627 -42198 30923 -41902
rect 30923 -42198 30927 -41902
rect 30623 -42202 30927 -42198
rect 30963 -41902 31587 -41898
rect 30963 -42198 30967 -41902
rect 30967 -42198 31583 -41902
rect 31583 -42198 31587 -41902
rect 30963 -42202 31587 -42198
rect 31623 -41902 31927 -41898
rect 31623 -42198 31627 -41902
rect 31627 -42198 31923 -41902
rect 31923 -42198 31927 -41902
rect 31623 -42202 31927 -42198
rect 31963 -41902 32587 -41898
rect 31963 -42198 31967 -41902
rect 31967 -42198 32583 -41902
rect 32583 -42198 32587 -41902
rect 31963 -42202 32587 -42198
rect 32623 -41902 32927 -41898
rect 32623 -42198 32627 -41902
rect 32627 -42198 32923 -41902
rect 32923 -42198 32927 -41902
rect 32623 -42202 32927 -42198
rect 32963 -41902 33587 -41898
rect 32963 -42198 32967 -41902
rect 32967 -42198 33583 -41902
rect 33583 -42198 33587 -41902
rect 32963 -42202 33587 -42198
rect 33623 -41902 33927 -41898
rect 33623 -42198 33627 -41902
rect 33627 -42198 33923 -41902
rect 33923 -42198 33927 -41902
rect 33623 -42202 33927 -42198
rect 33963 -41902 34267 -41898
rect 33963 -42198 33967 -41902
rect 33967 -42198 34263 -41902
rect 34263 -42198 34267 -41902
rect 33963 -42202 34267 -42198
rect 8623 -42242 8927 -42238
rect 8623 -42858 8627 -42242
rect 8627 -42858 8923 -42242
rect 8923 -42858 8927 -42242
rect 8623 -42862 8927 -42858
rect 9623 -42242 9927 -42238
rect 9623 -42858 9627 -42242
rect 9627 -42858 9923 -42242
rect 9923 -42858 9927 -42242
rect 9623 -42862 9927 -42858
rect 10623 -42242 10927 -42238
rect 10623 -42858 10627 -42242
rect 10627 -42858 10923 -42242
rect 10923 -42858 10927 -42242
rect 10623 -42862 10927 -42858
rect 11623 -42242 11927 -42238
rect 11623 -42858 11627 -42242
rect 11627 -42858 11923 -42242
rect 11923 -42858 11927 -42242
rect 11623 -42862 11927 -42858
rect 12623 -42242 12927 -42238
rect 12623 -42858 12627 -42242
rect 12627 -42858 12923 -42242
rect 12923 -42858 12927 -42242
rect 12623 -42862 12927 -42858
rect 13623 -42242 13927 -42238
rect 13623 -42858 13627 -42242
rect 13627 -42858 13923 -42242
rect 13923 -42858 13927 -42242
rect 13623 -42862 13927 -42858
rect 14623 -42242 14927 -42238
rect 14623 -42858 14627 -42242
rect 14627 -42858 14923 -42242
rect 14923 -42858 14927 -42242
rect 14623 -42862 14927 -42858
rect 15623 -42242 15927 -42238
rect 15623 -42858 15627 -42242
rect 15627 -42858 15923 -42242
rect 15923 -42858 15927 -42242
rect 15623 -42862 15927 -42858
rect 16623 -42242 16927 -42238
rect 16623 -42858 16627 -42242
rect 16627 -42858 16923 -42242
rect 16923 -42858 16927 -42242
rect 16623 -42862 16927 -42858
rect 17623 -42242 17927 -42238
rect 17623 -42858 17627 -42242
rect 17627 -42858 17923 -42242
rect 17923 -42858 17927 -42242
rect 17623 -42862 17927 -42858
rect 18623 -42242 18927 -42238
rect 18623 -42858 18627 -42242
rect 18627 -42858 18923 -42242
rect 18923 -42858 18927 -42242
rect 18623 -42862 18927 -42858
rect 19623 -42242 19927 -42238
rect 19623 -42858 19627 -42242
rect 19627 -42858 19923 -42242
rect 19923 -42858 19927 -42242
rect 19623 -42862 19927 -42858
rect 20623 -42242 20927 -42238
rect 20623 -42858 20627 -42242
rect 20627 -42858 20923 -42242
rect 20923 -42858 20927 -42242
rect 20623 -42862 20927 -42858
rect 21623 -42242 21927 -42238
rect 21623 -42858 21627 -42242
rect 21627 -42858 21923 -42242
rect 21923 -42858 21927 -42242
rect 21623 -42862 21927 -42858
rect 22623 -42242 22927 -42238
rect 22623 -42858 22627 -42242
rect 22627 -42858 22923 -42242
rect 22923 -42858 22927 -42242
rect 22623 -42862 22927 -42858
rect 23623 -42242 23927 -42238
rect 23623 -42858 23627 -42242
rect 23627 -42858 23923 -42242
rect 23923 -42858 23927 -42242
rect 23623 -42862 23927 -42858
rect 24623 -42242 24927 -42238
rect 24623 -42858 24627 -42242
rect 24627 -42858 24923 -42242
rect 24923 -42858 24927 -42242
rect 24623 -42862 24927 -42858
rect 25623 -42242 25927 -42238
rect 25623 -42858 25627 -42242
rect 25627 -42858 25923 -42242
rect 25923 -42858 25927 -42242
rect 25623 -42862 25927 -42858
rect 26623 -42242 26927 -42238
rect 26623 -42858 26627 -42242
rect 26627 -42858 26923 -42242
rect 26923 -42858 26927 -42242
rect 26623 -42862 26927 -42858
rect 27623 -42242 27927 -42238
rect 27623 -42858 27627 -42242
rect 27627 -42858 27923 -42242
rect 27923 -42858 27927 -42242
rect 27623 -42862 27927 -42858
rect 28623 -42242 28927 -42238
rect 28623 -42858 28627 -42242
rect 28627 -42858 28923 -42242
rect 28923 -42858 28927 -42242
rect 28623 -42862 28927 -42858
rect 29623 -42242 29927 -42238
rect 29623 -42858 29627 -42242
rect 29627 -42858 29923 -42242
rect 29923 -42858 29927 -42242
rect 29623 -42862 29927 -42858
rect 30623 -42242 30927 -42238
rect 30623 -42858 30627 -42242
rect 30627 -42858 30923 -42242
rect 30923 -42858 30927 -42242
rect 30623 -42862 30927 -42858
rect 31623 -42242 31927 -42238
rect 31623 -42858 31627 -42242
rect 31627 -42858 31923 -42242
rect 31923 -42858 31927 -42242
rect 31623 -42862 31927 -42858
rect 32623 -42242 32927 -42238
rect 32623 -42858 32627 -42242
rect 32627 -42858 32923 -42242
rect 32923 -42858 32927 -42242
rect 32623 -42862 32927 -42858
rect 33623 -42242 33927 -42238
rect 33623 -42858 33627 -42242
rect 33627 -42858 33923 -42242
rect 33923 -42858 33927 -42242
rect 33623 -42862 33927 -42858
rect 8283 -42902 8587 -42898
rect 8283 -43198 8287 -42902
rect 8287 -43198 8583 -42902
rect 8583 -43198 8587 -42902
rect 8283 -43202 8587 -43198
rect 8623 -42902 8927 -42898
rect 8623 -43198 8627 -42902
rect 8627 -43198 8923 -42902
rect 8923 -43198 8927 -42902
rect 8623 -43202 8927 -43198
rect 8963 -42902 9587 -42898
rect 8963 -43198 8967 -42902
rect 8967 -43198 9583 -42902
rect 9583 -43198 9587 -42902
rect 8963 -43202 9587 -43198
rect 9623 -42902 9927 -42898
rect 9623 -43198 9627 -42902
rect 9627 -43198 9923 -42902
rect 9923 -43198 9927 -42902
rect 9623 -43202 9927 -43198
rect 9963 -42902 10587 -42898
rect 9963 -43198 9967 -42902
rect 9967 -43198 10583 -42902
rect 10583 -43198 10587 -42902
rect 9963 -43202 10587 -43198
rect 10623 -42902 10927 -42898
rect 10623 -43198 10627 -42902
rect 10627 -43198 10923 -42902
rect 10923 -43198 10927 -42902
rect 10623 -43202 10927 -43198
rect 10963 -42902 11587 -42898
rect 10963 -43198 10967 -42902
rect 10967 -43198 11583 -42902
rect 11583 -43198 11587 -42902
rect 10963 -43202 11587 -43198
rect 11623 -42902 11927 -42898
rect 11623 -43198 11627 -42902
rect 11627 -43198 11923 -42902
rect 11923 -43198 11927 -42902
rect 11623 -43202 11927 -43198
rect 11963 -42902 12587 -42898
rect 11963 -43198 11967 -42902
rect 11967 -43198 12583 -42902
rect 12583 -43198 12587 -42902
rect 11963 -43202 12587 -43198
rect 12623 -42902 12927 -42898
rect 12623 -43198 12627 -42902
rect 12627 -43198 12923 -42902
rect 12923 -43198 12927 -42902
rect 12623 -43202 12927 -43198
rect 12963 -42902 13587 -42898
rect 12963 -43198 12967 -42902
rect 12967 -43198 13583 -42902
rect 13583 -43198 13587 -42902
rect 12963 -43202 13587 -43198
rect 13623 -42902 13927 -42898
rect 13623 -43198 13627 -42902
rect 13627 -43198 13923 -42902
rect 13923 -43198 13927 -42902
rect 13623 -43202 13927 -43198
rect 13963 -42902 14587 -42898
rect 13963 -43198 13967 -42902
rect 13967 -43198 14583 -42902
rect 14583 -43198 14587 -42902
rect 13963 -43202 14587 -43198
rect 14623 -42902 14927 -42898
rect 14623 -43198 14627 -42902
rect 14627 -43198 14923 -42902
rect 14923 -43198 14927 -42902
rect 14623 -43202 14927 -43198
rect 14963 -42902 15587 -42898
rect 14963 -43198 14967 -42902
rect 14967 -43198 15583 -42902
rect 15583 -43198 15587 -42902
rect 14963 -43202 15587 -43198
rect 15623 -42902 15927 -42898
rect 15623 -43198 15627 -42902
rect 15627 -43198 15923 -42902
rect 15923 -43198 15927 -42902
rect 15623 -43202 15927 -43198
rect 15963 -42902 16587 -42898
rect 15963 -43198 15967 -42902
rect 15967 -43198 16583 -42902
rect 16583 -43198 16587 -42902
rect 15963 -43202 16587 -43198
rect 16623 -42902 16927 -42898
rect 16623 -43198 16627 -42902
rect 16627 -43198 16923 -42902
rect 16923 -43198 16927 -42902
rect 16623 -43202 16927 -43198
rect 16963 -42902 17587 -42898
rect 16963 -43198 16967 -42902
rect 16967 -43198 17583 -42902
rect 17583 -43198 17587 -42902
rect 16963 -43202 17587 -43198
rect 17623 -42902 17927 -42898
rect 17623 -43198 17627 -42902
rect 17627 -43198 17923 -42902
rect 17923 -43198 17927 -42902
rect 17623 -43202 17927 -43198
rect 17963 -42902 18587 -42898
rect 17963 -43198 17967 -42902
rect 17967 -43198 18583 -42902
rect 18583 -43198 18587 -42902
rect 17963 -43202 18587 -43198
rect 18623 -42902 18927 -42898
rect 18623 -43198 18627 -42902
rect 18627 -43198 18923 -42902
rect 18923 -43198 18927 -42902
rect 18623 -43202 18927 -43198
rect 18963 -42902 19587 -42898
rect 18963 -43198 18967 -42902
rect 18967 -43198 19583 -42902
rect 19583 -43198 19587 -42902
rect 18963 -43202 19587 -43198
rect 19623 -42902 19927 -42898
rect 19623 -43198 19627 -42902
rect 19627 -43198 19923 -42902
rect 19923 -43198 19927 -42902
rect 19623 -43202 19927 -43198
rect 19963 -42902 20587 -42898
rect 19963 -43198 19967 -42902
rect 19967 -43198 20583 -42902
rect 20583 -43198 20587 -42902
rect 19963 -43202 20587 -43198
rect 20623 -42902 20927 -42898
rect 20623 -43198 20627 -42902
rect 20627 -43198 20923 -42902
rect 20923 -43198 20927 -42902
rect 20623 -43202 20927 -43198
rect 20963 -42902 21587 -42898
rect 20963 -43198 20967 -42902
rect 20967 -43198 21583 -42902
rect 21583 -43198 21587 -42902
rect 20963 -43202 21587 -43198
rect 21623 -42902 21927 -42898
rect 21623 -43198 21627 -42902
rect 21627 -43198 21923 -42902
rect 21923 -43198 21927 -42902
rect 21623 -43202 21927 -43198
rect 21963 -42902 22587 -42898
rect 21963 -43198 21967 -42902
rect 21967 -43198 22583 -42902
rect 22583 -43198 22587 -42902
rect 21963 -43202 22587 -43198
rect 22623 -42902 22927 -42898
rect 22623 -43198 22627 -42902
rect 22627 -43198 22923 -42902
rect 22923 -43198 22927 -42902
rect 22623 -43202 22927 -43198
rect 22963 -42902 23587 -42898
rect 22963 -43198 22967 -42902
rect 22967 -43198 23583 -42902
rect 23583 -43198 23587 -42902
rect 22963 -43202 23587 -43198
rect 23623 -42902 23927 -42898
rect 23623 -43198 23627 -42902
rect 23627 -43198 23923 -42902
rect 23923 -43198 23927 -42902
rect 23623 -43202 23927 -43198
rect 23963 -42902 24587 -42898
rect 23963 -43198 23967 -42902
rect 23967 -43198 24583 -42902
rect 24583 -43198 24587 -42902
rect 23963 -43202 24587 -43198
rect 24623 -42902 24927 -42898
rect 24623 -43198 24627 -42902
rect 24627 -43198 24923 -42902
rect 24923 -43198 24927 -42902
rect 24623 -43202 24927 -43198
rect 24963 -42902 25587 -42898
rect 24963 -43198 24967 -42902
rect 24967 -43198 25583 -42902
rect 25583 -43198 25587 -42902
rect 24963 -43202 25587 -43198
rect 25623 -42902 25927 -42898
rect 25623 -43198 25627 -42902
rect 25627 -43198 25923 -42902
rect 25923 -43198 25927 -42902
rect 25623 -43202 25927 -43198
rect 25963 -42902 26587 -42898
rect 25963 -43198 25967 -42902
rect 25967 -43198 26583 -42902
rect 26583 -43198 26587 -42902
rect 25963 -43202 26587 -43198
rect 26623 -42902 26927 -42898
rect 26623 -43198 26627 -42902
rect 26627 -43198 26923 -42902
rect 26923 -43198 26927 -42902
rect 26623 -43202 26927 -43198
rect 26963 -42902 27587 -42898
rect 26963 -43198 26967 -42902
rect 26967 -43198 27583 -42902
rect 27583 -43198 27587 -42902
rect 26963 -43202 27587 -43198
rect 27623 -42902 27927 -42898
rect 27623 -43198 27627 -42902
rect 27627 -43198 27923 -42902
rect 27923 -43198 27927 -42902
rect 27623 -43202 27927 -43198
rect 27963 -42902 28587 -42898
rect 27963 -43198 27967 -42902
rect 27967 -43198 28583 -42902
rect 28583 -43198 28587 -42902
rect 27963 -43202 28587 -43198
rect 28623 -42902 28927 -42898
rect 28623 -43198 28627 -42902
rect 28627 -43198 28923 -42902
rect 28923 -43198 28927 -42902
rect 28623 -43202 28927 -43198
rect 28963 -42902 29587 -42898
rect 28963 -43198 28967 -42902
rect 28967 -43198 29583 -42902
rect 29583 -43198 29587 -42902
rect 28963 -43202 29587 -43198
rect 29623 -42902 29927 -42898
rect 29623 -43198 29627 -42902
rect 29627 -43198 29923 -42902
rect 29923 -43198 29927 -42902
rect 29623 -43202 29927 -43198
rect 29963 -42902 30587 -42898
rect 29963 -43198 29967 -42902
rect 29967 -43198 30583 -42902
rect 30583 -43198 30587 -42902
rect 29963 -43202 30587 -43198
rect 30623 -42902 30927 -42898
rect 30623 -43198 30627 -42902
rect 30627 -43198 30923 -42902
rect 30923 -43198 30927 -42902
rect 30623 -43202 30927 -43198
rect 30963 -42902 31587 -42898
rect 30963 -43198 30967 -42902
rect 30967 -43198 31583 -42902
rect 31583 -43198 31587 -42902
rect 30963 -43202 31587 -43198
rect 31623 -42902 31927 -42898
rect 31623 -43198 31627 -42902
rect 31627 -43198 31923 -42902
rect 31923 -43198 31927 -42902
rect 31623 -43202 31927 -43198
rect 31963 -42902 32587 -42898
rect 31963 -43198 31967 -42902
rect 31967 -43198 32583 -42902
rect 32583 -43198 32587 -42902
rect 31963 -43202 32587 -43198
rect 32623 -42902 32927 -42898
rect 32623 -43198 32627 -42902
rect 32627 -43198 32923 -42902
rect 32923 -43198 32927 -42902
rect 32623 -43202 32927 -43198
rect 32963 -42902 33587 -42898
rect 32963 -43198 32967 -42902
rect 32967 -43198 33583 -42902
rect 33583 -43198 33587 -42902
rect 32963 -43202 33587 -43198
rect 33623 -42902 33927 -42898
rect 33623 -43198 33627 -42902
rect 33627 -43198 33923 -42902
rect 33923 -43198 33927 -42902
rect 33623 -43202 33927 -43198
rect 33963 -42902 34267 -42898
rect 33963 -43198 33967 -42902
rect 33967 -43198 34263 -42902
rect 34263 -43198 34267 -42902
rect 33963 -43202 34267 -43198
rect 8623 -43242 8927 -43238
rect 8623 -43858 8627 -43242
rect 8627 -43858 8923 -43242
rect 8923 -43858 8927 -43242
rect 8623 -43862 8927 -43858
rect 9623 -43242 9927 -43238
rect 9623 -43858 9627 -43242
rect 9627 -43858 9923 -43242
rect 9923 -43858 9927 -43242
rect 9623 -43862 9927 -43858
rect 10623 -43242 10927 -43238
rect 10623 -43858 10627 -43242
rect 10627 -43858 10923 -43242
rect 10923 -43858 10927 -43242
rect 10623 -43862 10927 -43858
rect 11623 -43242 11927 -43238
rect 11623 -43858 11627 -43242
rect 11627 -43858 11923 -43242
rect 11923 -43858 11927 -43242
rect 11623 -43862 11927 -43858
rect 12623 -43242 12927 -43238
rect 12623 -43858 12627 -43242
rect 12627 -43858 12923 -43242
rect 12923 -43858 12927 -43242
rect 12623 -43862 12927 -43858
rect 13623 -43242 13927 -43238
rect 13623 -43858 13627 -43242
rect 13627 -43858 13923 -43242
rect 13923 -43858 13927 -43242
rect 13623 -43862 13927 -43858
rect 14623 -43242 14927 -43238
rect 14623 -43858 14627 -43242
rect 14627 -43858 14923 -43242
rect 14923 -43858 14927 -43242
rect 14623 -43862 14927 -43858
rect 15623 -43242 15927 -43238
rect 15623 -43858 15627 -43242
rect 15627 -43858 15923 -43242
rect 15923 -43858 15927 -43242
rect 15623 -43862 15927 -43858
rect 16623 -43242 16927 -43238
rect 16623 -43858 16627 -43242
rect 16627 -43858 16923 -43242
rect 16923 -43858 16927 -43242
rect 16623 -43862 16927 -43858
rect 17623 -43242 17927 -43238
rect 17623 -43858 17627 -43242
rect 17627 -43858 17923 -43242
rect 17923 -43858 17927 -43242
rect 17623 -43862 17927 -43858
rect 18623 -43242 18927 -43238
rect 18623 -43858 18627 -43242
rect 18627 -43858 18923 -43242
rect 18923 -43858 18927 -43242
rect 18623 -43862 18927 -43858
rect 19623 -43242 19927 -43238
rect 19623 -43858 19627 -43242
rect 19627 -43858 19923 -43242
rect 19923 -43858 19927 -43242
rect 19623 -43862 19927 -43858
rect 20623 -43242 20927 -43238
rect 20623 -43858 20627 -43242
rect 20627 -43858 20923 -43242
rect 20923 -43858 20927 -43242
rect 20623 -43862 20927 -43858
rect 21623 -43242 21927 -43238
rect 21623 -43858 21627 -43242
rect 21627 -43858 21923 -43242
rect 21923 -43858 21927 -43242
rect 21623 -43862 21927 -43858
rect 22623 -43242 22927 -43238
rect 22623 -43858 22627 -43242
rect 22627 -43858 22923 -43242
rect 22923 -43858 22927 -43242
rect 22623 -43862 22927 -43858
rect 23623 -43242 23927 -43238
rect 23623 -43858 23627 -43242
rect 23627 -43858 23923 -43242
rect 23923 -43858 23927 -43242
rect 23623 -43862 23927 -43858
rect 24623 -43242 24927 -43238
rect 24623 -43858 24627 -43242
rect 24627 -43858 24923 -43242
rect 24923 -43858 24927 -43242
rect 24623 -43862 24927 -43858
rect 25623 -43242 25927 -43238
rect 25623 -43858 25627 -43242
rect 25627 -43858 25923 -43242
rect 25923 -43858 25927 -43242
rect 25623 -43862 25927 -43858
rect 26623 -43242 26927 -43238
rect 26623 -43858 26627 -43242
rect 26627 -43858 26923 -43242
rect 26923 -43858 26927 -43242
rect 26623 -43862 26927 -43858
rect 27623 -43242 27927 -43238
rect 27623 -43858 27627 -43242
rect 27627 -43858 27923 -43242
rect 27923 -43858 27927 -43242
rect 27623 -43862 27927 -43858
rect 28623 -43242 28927 -43238
rect 28623 -43858 28627 -43242
rect 28627 -43858 28923 -43242
rect 28923 -43858 28927 -43242
rect 28623 -43862 28927 -43858
rect 29623 -43242 29927 -43238
rect 29623 -43858 29627 -43242
rect 29627 -43858 29923 -43242
rect 29923 -43858 29927 -43242
rect 29623 -43862 29927 -43858
rect 30623 -43242 30927 -43238
rect 30623 -43858 30627 -43242
rect 30627 -43858 30923 -43242
rect 30923 -43858 30927 -43242
rect 30623 -43862 30927 -43858
rect 31623 -43242 31927 -43238
rect 31623 -43858 31627 -43242
rect 31627 -43858 31923 -43242
rect 31923 -43858 31927 -43242
rect 31623 -43862 31927 -43858
rect 32623 -43242 32927 -43238
rect 32623 -43858 32627 -43242
rect 32627 -43858 32923 -43242
rect 32923 -43858 32927 -43242
rect 32623 -43862 32927 -43858
rect 33623 -43242 33927 -43238
rect 33623 -43858 33627 -43242
rect 33627 -43858 33923 -43242
rect 33923 -43858 33927 -43242
rect 33623 -43862 33927 -43858
rect 8283 -43902 8587 -43898
rect 8283 -44198 8287 -43902
rect 8287 -44198 8583 -43902
rect 8583 -44198 8587 -43902
rect 8283 -44202 8587 -44198
rect 8623 -43902 8927 -43898
rect 8623 -44198 8627 -43902
rect 8627 -44198 8923 -43902
rect 8923 -44198 8927 -43902
rect 8623 -44202 8927 -44198
rect 8963 -43902 9587 -43898
rect 8963 -44198 8967 -43902
rect 8967 -44198 9583 -43902
rect 9583 -44198 9587 -43902
rect 8963 -44202 9587 -44198
rect 9623 -43902 9927 -43898
rect 9623 -44198 9627 -43902
rect 9627 -44198 9923 -43902
rect 9923 -44198 9927 -43902
rect 9623 -44202 9927 -44198
rect 9963 -43902 10587 -43898
rect 9963 -44198 9967 -43902
rect 9967 -44198 10583 -43902
rect 10583 -44198 10587 -43902
rect 9963 -44202 10587 -44198
rect 10623 -43902 10927 -43898
rect 10623 -44198 10627 -43902
rect 10627 -44198 10923 -43902
rect 10923 -44198 10927 -43902
rect 10623 -44202 10927 -44198
rect 10963 -43902 11587 -43898
rect 10963 -44198 10967 -43902
rect 10967 -44198 11583 -43902
rect 11583 -44198 11587 -43902
rect 10963 -44202 11587 -44198
rect 11623 -43902 11927 -43898
rect 11623 -44198 11627 -43902
rect 11627 -44198 11923 -43902
rect 11923 -44198 11927 -43902
rect 11623 -44202 11927 -44198
rect 11963 -43902 12587 -43898
rect 11963 -44198 11967 -43902
rect 11967 -44198 12583 -43902
rect 12583 -44198 12587 -43902
rect 11963 -44202 12587 -44198
rect 12623 -43902 12927 -43898
rect 12623 -44198 12627 -43902
rect 12627 -44198 12923 -43902
rect 12923 -44198 12927 -43902
rect 12623 -44202 12927 -44198
rect 12963 -43902 13587 -43898
rect 12963 -44198 12967 -43902
rect 12967 -44198 13583 -43902
rect 13583 -44198 13587 -43902
rect 12963 -44202 13587 -44198
rect 13623 -43902 13927 -43898
rect 13623 -44198 13627 -43902
rect 13627 -44198 13923 -43902
rect 13923 -44198 13927 -43902
rect 13623 -44202 13927 -44198
rect 13963 -43902 14587 -43898
rect 13963 -44198 13967 -43902
rect 13967 -44198 14583 -43902
rect 14583 -44198 14587 -43902
rect 13963 -44202 14587 -44198
rect 14623 -43902 14927 -43898
rect 14623 -44198 14627 -43902
rect 14627 -44198 14923 -43902
rect 14923 -44198 14927 -43902
rect 14623 -44202 14927 -44198
rect 14963 -43902 15587 -43898
rect 14963 -44198 14967 -43902
rect 14967 -44198 15583 -43902
rect 15583 -44198 15587 -43902
rect 14963 -44202 15587 -44198
rect 15623 -43902 15927 -43898
rect 15623 -44198 15627 -43902
rect 15627 -44198 15923 -43902
rect 15923 -44198 15927 -43902
rect 15623 -44202 15927 -44198
rect 15963 -43902 16587 -43898
rect 15963 -44198 15967 -43902
rect 15967 -44198 16583 -43902
rect 16583 -44198 16587 -43902
rect 15963 -44202 16587 -44198
rect 16623 -43902 16927 -43898
rect 16623 -44198 16627 -43902
rect 16627 -44198 16923 -43902
rect 16923 -44198 16927 -43902
rect 16623 -44202 16927 -44198
rect 16963 -43902 17587 -43898
rect 16963 -44198 16967 -43902
rect 16967 -44198 17583 -43902
rect 17583 -44198 17587 -43902
rect 16963 -44202 17587 -44198
rect 17623 -43902 17927 -43898
rect 17623 -44198 17627 -43902
rect 17627 -44198 17923 -43902
rect 17923 -44198 17927 -43902
rect 17623 -44202 17927 -44198
rect 17963 -43902 18587 -43898
rect 17963 -44198 17967 -43902
rect 17967 -44198 18583 -43902
rect 18583 -44198 18587 -43902
rect 17963 -44202 18587 -44198
rect 18623 -43902 18927 -43898
rect 18623 -44198 18627 -43902
rect 18627 -44198 18923 -43902
rect 18923 -44198 18927 -43902
rect 18623 -44202 18927 -44198
rect 18963 -43902 19587 -43898
rect 18963 -44198 18967 -43902
rect 18967 -44198 19583 -43902
rect 19583 -44198 19587 -43902
rect 18963 -44202 19587 -44198
rect 19623 -43902 19927 -43898
rect 19623 -44198 19627 -43902
rect 19627 -44198 19923 -43902
rect 19923 -44198 19927 -43902
rect 19623 -44202 19927 -44198
rect 19963 -43902 20587 -43898
rect 19963 -44198 19967 -43902
rect 19967 -44198 20583 -43902
rect 20583 -44198 20587 -43902
rect 19963 -44202 20587 -44198
rect 20623 -43902 20927 -43898
rect 20623 -44198 20627 -43902
rect 20627 -44198 20923 -43902
rect 20923 -44198 20927 -43902
rect 20623 -44202 20927 -44198
rect 20963 -43902 21587 -43898
rect 20963 -44198 20967 -43902
rect 20967 -44198 21583 -43902
rect 21583 -44198 21587 -43902
rect 20963 -44202 21587 -44198
rect 21623 -43902 21927 -43898
rect 21623 -44198 21627 -43902
rect 21627 -44198 21923 -43902
rect 21923 -44198 21927 -43902
rect 21623 -44202 21927 -44198
rect 21963 -43902 22587 -43898
rect 21963 -44198 21967 -43902
rect 21967 -44198 22583 -43902
rect 22583 -44198 22587 -43902
rect 21963 -44202 22587 -44198
rect 22623 -43902 22927 -43898
rect 22623 -44198 22627 -43902
rect 22627 -44198 22923 -43902
rect 22923 -44198 22927 -43902
rect 22623 -44202 22927 -44198
rect 22963 -43902 23587 -43898
rect 22963 -44198 22967 -43902
rect 22967 -44198 23583 -43902
rect 23583 -44198 23587 -43902
rect 22963 -44202 23587 -44198
rect 23623 -43902 23927 -43898
rect 23623 -44198 23627 -43902
rect 23627 -44198 23923 -43902
rect 23923 -44198 23927 -43902
rect 23623 -44202 23927 -44198
rect 23963 -43902 24587 -43898
rect 23963 -44198 23967 -43902
rect 23967 -44198 24583 -43902
rect 24583 -44198 24587 -43902
rect 23963 -44202 24587 -44198
rect 24623 -43902 24927 -43898
rect 24623 -44198 24627 -43902
rect 24627 -44198 24923 -43902
rect 24923 -44198 24927 -43902
rect 24623 -44202 24927 -44198
rect 24963 -43902 25587 -43898
rect 24963 -44198 24967 -43902
rect 24967 -44198 25583 -43902
rect 25583 -44198 25587 -43902
rect 24963 -44202 25587 -44198
rect 25623 -43902 25927 -43898
rect 25623 -44198 25627 -43902
rect 25627 -44198 25923 -43902
rect 25923 -44198 25927 -43902
rect 25623 -44202 25927 -44198
rect 25963 -43902 26587 -43898
rect 25963 -44198 25967 -43902
rect 25967 -44198 26583 -43902
rect 26583 -44198 26587 -43902
rect 25963 -44202 26587 -44198
rect 26623 -43902 26927 -43898
rect 26623 -44198 26627 -43902
rect 26627 -44198 26923 -43902
rect 26923 -44198 26927 -43902
rect 26623 -44202 26927 -44198
rect 26963 -43902 27587 -43898
rect 26963 -44198 26967 -43902
rect 26967 -44198 27583 -43902
rect 27583 -44198 27587 -43902
rect 26963 -44202 27587 -44198
rect 27623 -43902 27927 -43898
rect 27623 -44198 27627 -43902
rect 27627 -44198 27923 -43902
rect 27923 -44198 27927 -43902
rect 27623 -44202 27927 -44198
rect 27963 -43902 28587 -43898
rect 27963 -44198 27967 -43902
rect 27967 -44198 28583 -43902
rect 28583 -44198 28587 -43902
rect 27963 -44202 28587 -44198
rect 28623 -43902 28927 -43898
rect 28623 -44198 28627 -43902
rect 28627 -44198 28923 -43902
rect 28923 -44198 28927 -43902
rect 28623 -44202 28927 -44198
rect 28963 -43902 29587 -43898
rect 28963 -44198 28967 -43902
rect 28967 -44198 29583 -43902
rect 29583 -44198 29587 -43902
rect 28963 -44202 29587 -44198
rect 29623 -43902 29927 -43898
rect 29623 -44198 29627 -43902
rect 29627 -44198 29923 -43902
rect 29923 -44198 29927 -43902
rect 29623 -44202 29927 -44198
rect 29963 -43902 30587 -43898
rect 29963 -44198 29967 -43902
rect 29967 -44198 30583 -43902
rect 30583 -44198 30587 -43902
rect 29963 -44202 30587 -44198
rect 30623 -43902 30927 -43898
rect 30623 -44198 30627 -43902
rect 30627 -44198 30923 -43902
rect 30923 -44198 30927 -43902
rect 30623 -44202 30927 -44198
rect 30963 -43902 31587 -43898
rect 30963 -44198 30967 -43902
rect 30967 -44198 31583 -43902
rect 31583 -44198 31587 -43902
rect 30963 -44202 31587 -44198
rect 31623 -43902 31927 -43898
rect 31623 -44198 31627 -43902
rect 31627 -44198 31923 -43902
rect 31923 -44198 31927 -43902
rect 31623 -44202 31927 -44198
rect 31963 -43902 32587 -43898
rect 31963 -44198 31967 -43902
rect 31967 -44198 32583 -43902
rect 32583 -44198 32587 -43902
rect 31963 -44202 32587 -44198
rect 32623 -43902 32927 -43898
rect 32623 -44198 32627 -43902
rect 32627 -44198 32923 -43902
rect 32923 -44198 32927 -43902
rect 32623 -44202 32927 -44198
rect 32963 -43902 33587 -43898
rect 32963 -44198 32967 -43902
rect 32967 -44198 33583 -43902
rect 33583 -44198 33587 -43902
rect 32963 -44202 33587 -44198
rect 33623 -43902 33927 -43898
rect 33623 -44198 33627 -43902
rect 33627 -44198 33923 -43902
rect 33923 -44198 33927 -43902
rect 33623 -44202 33927 -44198
rect 33963 -43902 34267 -43898
rect 33963 -44198 33967 -43902
rect 33967 -44198 34263 -43902
rect 34263 -44198 34267 -43902
rect 33963 -44202 34267 -44198
rect 8623 -44242 8927 -44238
rect 8623 -44858 8627 -44242
rect 8627 -44858 8923 -44242
rect 8923 -44858 8927 -44242
rect 8623 -44862 8927 -44858
rect 9623 -44242 9927 -44238
rect 9623 -44858 9627 -44242
rect 9627 -44858 9923 -44242
rect 9923 -44858 9927 -44242
rect 9623 -44862 9927 -44858
rect 10623 -44242 10927 -44238
rect 10623 -44858 10627 -44242
rect 10627 -44858 10923 -44242
rect 10923 -44858 10927 -44242
rect 10623 -44862 10927 -44858
rect 11623 -44242 11927 -44238
rect 11623 -44858 11627 -44242
rect 11627 -44858 11923 -44242
rect 11923 -44858 11927 -44242
rect 11623 -44862 11927 -44858
rect 12623 -44242 12927 -44238
rect 12623 -44858 12627 -44242
rect 12627 -44858 12923 -44242
rect 12923 -44858 12927 -44242
rect 12623 -44862 12927 -44858
rect 13623 -44242 13927 -44238
rect 13623 -44858 13627 -44242
rect 13627 -44858 13923 -44242
rect 13923 -44858 13927 -44242
rect 13623 -44862 13927 -44858
rect 14623 -44242 14927 -44238
rect 14623 -44858 14627 -44242
rect 14627 -44858 14923 -44242
rect 14923 -44858 14927 -44242
rect 14623 -44862 14927 -44858
rect 15623 -44242 15927 -44238
rect 15623 -44858 15627 -44242
rect 15627 -44858 15923 -44242
rect 15923 -44858 15927 -44242
rect 15623 -44862 15927 -44858
rect 16623 -44242 16927 -44238
rect 16623 -44858 16627 -44242
rect 16627 -44858 16923 -44242
rect 16923 -44858 16927 -44242
rect 16623 -44862 16927 -44858
rect 17623 -44242 17927 -44238
rect 17623 -44858 17627 -44242
rect 17627 -44858 17923 -44242
rect 17923 -44858 17927 -44242
rect 17623 -44862 17927 -44858
rect 18623 -44242 18927 -44238
rect 18623 -44858 18627 -44242
rect 18627 -44858 18923 -44242
rect 18923 -44858 18927 -44242
rect 18623 -44862 18927 -44858
rect 19623 -44242 19927 -44238
rect 19623 -44858 19627 -44242
rect 19627 -44858 19923 -44242
rect 19923 -44858 19927 -44242
rect 19623 -44862 19927 -44858
rect 20623 -44242 20927 -44238
rect 20623 -44858 20627 -44242
rect 20627 -44858 20923 -44242
rect 20923 -44858 20927 -44242
rect 20623 -44862 20927 -44858
rect 21623 -44242 21927 -44238
rect 21623 -44858 21627 -44242
rect 21627 -44858 21923 -44242
rect 21923 -44858 21927 -44242
rect 21623 -44862 21927 -44858
rect 22623 -44242 22927 -44238
rect 22623 -44858 22627 -44242
rect 22627 -44858 22923 -44242
rect 22923 -44858 22927 -44242
rect 22623 -44862 22927 -44858
rect 23623 -44242 23927 -44238
rect 23623 -44858 23627 -44242
rect 23627 -44858 23923 -44242
rect 23923 -44858 23927 -44242
rect 23623 -44862 23927 -44858
rect 24623 -44242 24927 -44238
rect 24623 -44858 24627 -44242
rect 24627 -44858 24923 -44242
rect 24923 -44858 24927 -44242
rect 24623 -44862 24927 -44858
rect 25623 -44242 25927 -44238
rect 25623 -44858 25627 -44242
rect 25627 -44858 25923 -44242
rect 25923 -44858 25927 -44242
rect 25623 -44862 25927 -44858
rect 26623 -44242 26927 -44238
rect 26623 -44858 26627 -44242
rect 26627 -44858 26923 -44242
rect 26923 -44858 26927 -44242
rect 26623 -44862 26927 -44858
rect 27623 -44242 27927 -44238
rect 27623 -44858 27627 -44242
rect 27627 -44858 27923 -44242
rect 27923 -44858 27927 -44242
rect 27623 -44862 27927 -44858
rect 28623 -44242 28927 -44238
rect 28623 -44858 28627 -44242
rect 28627 -44858 28923 -44242
rect 28923 -44858 28927 -44242
rect 28623 -44862 28927 -44858
rect 29623 -44242 29927 -44238
rect 29623 -44858 29627 -44242
rect 29627 -44858 29923 -44242
rect 29923 -44858 29927 -44242
rect 29623 -44862 29927 -44858
rect 30623 -44242 30927 -44238
rect 30623 -44858 30627 -44242
rect 30627 -44858 30923 -44242
rect 30923 -44858 30927 -44242
rect 30623 -44862 30927 -44858
rect 31623 -44242 31927 -44238
rect 31623 -44858 31627 -44242
rect 31627 -44858 31923 -44242
rect 31923 -44858 31927 -44242
rect 31623 -44862 31927 -44858
rect 32623 -44242 32927 -44238
rect 32623 -44858 32627 -44242
rect 32627 -44858 32923 -44242
rect 32923 -44858 32927 -44242
rect 32623 -44862 32927 -44858
rect 33623 -44242 33927 -44238
rect 33623 -44858 33627 -44242
rect 33627 -44858 33923 -44242
rect 33923 -44858 33927 -44242
rect 33623 -44862 33927 -44858
rect -74817 -44902 -74513 -44898
rect -74817 -45198 -74813 -44902
rect -74813 -45198 -74517 -44902
rect -74517 -45198 -74513 -44902
rect -74817 -45202 -74513 -45198
rect -74477 -44902 -74173 -44898
rect -74477 -45198 -74473 -44902
rect -74473 -45198 -74177 -44902
rect -74177 -45198 -74173 -44902
rect -74477 -45202 -74173 -45198
rect -74137 -44902 -73513 -44898
rect -74137 -45198 -74133 -44902
rect -74133 -45198 -73517 -44902
rect -73517 -45198 -73513 -44902
rect -74137 -45202 -73513 -45198
rect -73477 -44902 -73173 -44898
rect -73477 -45198 -73473 -44902
rect -73473 -45198 -73177 -44902
rect -73177 -45198 -73173 -44902
rect -73477 -45202 -73173 -45198
rect -73137 -44902 -72513 -44898
rect -73137 -45198 -73133 -44902
rect -73133 -45198 -72517 -44902
rect -72517 -45198 -72513 -44902
rect -73137 -45202 -72513 -45198
rect -72477 -44902 -72173 -44898
rect -72477 -45198 -72473 -44902
rect -72473 -45198 -72177 -44902
rect -72177 -45198 -72173 -44902
rect -72477 -45202 -72173 -45198
rect -72137 -44902 -71513 -44898
rect -72137 -45198 -72133 -44902
rect -72133 -45198 -71517 -44902
rect -71517 -45198 -71513 -44902
rect -72137 -45202 -71513 -45198
rect -71477 -44902 -71173 -44898
rect -71477 -45198 -71473 -44902
rect -71473 -45198 -71177 -44902
rect -71177 -45198 -71173 -44902
rect -71477 -45202 -71173 -45198
rect -71137 -44902 -70513 -44898
rect -71137 -45198 -71133 -44902
rect -71133 -45198 -70517 -44902
rect -70517 -45198 -70513 -44902
rect -71137 -45202 -70513 -45198
rect -70477 -44902 -70173 -44898
rect -70477 -45198 -70473 -44902
rect -70473 -45198 -70177 -44902
rect -70177 -45198 -70173 -44902
rect -70477 -45202 -70173 -45198
rect -70137 -44902 -69513 -44898
rect -70137 -45198 -70133 -44902
rect -70133 -45198 -69517 -44902
rect -69517 -45198 -69513 -44902
rect -70137 -45202 -69513 -45198
rect -69477 -44902 -69173 -44898
rect -69477 -45198 -69473 -44902
rect -69473 -45198 -69177 -44902
rect -69177 -45198 -69173 -44902
rect -69477 -45202 -69173 -45198
rect -69137 -44902 -68513 -44898
rect -69137 -45198 -69133 -44902
rect -69133 -45198 -68517 -44902
rect -68517 -45198 -68513 -44902
rect -69137 -45202 -68513 -45198
rect -68477 -44902 -68173 -44898
rect -68477 -45198 -68473 -44902
rect -68473 -45198 -68177 -44902
rect -68177 -45198 -68173 -44902
rect -68477 -45202 -68173 -45198
rect -68137 -44902 -67513 -44898
rect -68137 -45198 -68133 -44902
rect -68133 -45198 -67517 -44902
rect -67517 -45198 -67513 -44902
rect -68137 -45202 -67513 -45198
rect -67477 -44902 -67173 -44898
rect -67477 -45198 -67473 -44902
rect -67473 -45198 -67177 -44902
rect -67177 -45198 -67173 -44902
rect -67477 -45202 -67173 -45198
rect -67137 -44902 -66513 -44898
rect -67137 -45198 -67133 -44902
rect -67133 -45198 -66517 -44902
rect -66517 -45198 -66513 -44902
rect -67137 -45202 -66513 -45198
rect -66477 -44902 -66173 -44898
rect -66477 -45198 -66473 -44902
rect -66473 -45198 -66177 -44902
rect -66177 -45198 -66173 -44902
rect -66477 -45202 -66173 -45198
rect -66137 -44902 -65513 -44898
rect -66137 -45198 -66133 -44902
rect -66133 -45198 -65517 -44902
rect -65517 -45198 -65513 -44902
rect -66137 -45202 -65513 -45198
rect -65477 -44902 -65173 -44898
rect -65477 -45198 -65473 -44902
rect -65473 -45198 -65177 -44902
rect -65177 -45198 -65173 -44902
rect -65477 -45202 -65173 -45198
rect -65137 -44902 -64513 -44898
rect -65137 -45198 -65133 -44902
rect -65133 -45198 -64517 -44902
rect -64517 -45198 -64513 -44902
rect -65137 -45202 -64513 -45198
rect -64477 -44902 -64173 -44898
rect -64477 -45198 -64473 -44902
rect -64473 -45198 -64177 -44902
rect -64177 -45198 -64173 -44902
rect -64477 -45202 -64173 -45198
rect -64137 -44902 -63513 -44898
rect -64137 -45198 -64133 -44902
rect -64133 -45198 -63517 -44902
rect -63517 -45198 -63513 -44902
rect -64137 -45202 -63513 -45198
rect -63477 -44902 -63173 -44898
rect -63477 -45198 -63473 -44902
rect -63473 -45198 -63177 -44902
rect -63177 -45198 -63173 -44902
rect -63477 -45202 -63173 -45198
rect -63137 -44902 -62513 -44898
rect -63137 -45198 -63133 -44902
rect -63133 -45198 -62517 -44902
rect -62517 -45198 -62513 -44902
rect -63137 -45202 -62513 -45198
rect -62477 -44902 -62173 -44898
rect -62477 -45198 -62473 -44902
rect -62473 -45198 -62177 -44902
rect -62177 -45198 -62173 -44902
rect -62477 -45202 -62173 -45198
rect -62137 -44902 -61513 -44898
rect -62137 -45198 -62133 -44902
rect -62133 -45198 -61517 -44902
rect -61517 -45198 -61513 -44902
rect -62137 -45202 -61513 -45198
rect -61477 -44902 -61173 -44898
rect -61477 -45198 -61473 -44902
rect -61473 -45198 -61177 -44902
rect -61177 -45198 -61173 -44902
rect -61477 -45202 -61173 -45198
rect -61137 -44902 -60513 -44898
rect -61137 -45198 -61133 -44902
rect -61133 -45198 -60517 -44902
rect -60517 -45198 -60513 -44902
rect -61137 -45202 -60513 -45198
rect -60477 -44902 -60173 -44898
rect -60477 -45198 -60473 -44902
rect -60473 -45198 -60177 -44902
rect -60177 -45198 -60173 -44902
rect -60477 -45202 -60173 -45198
rect -60137 -44902 -59513 -44898
rect -60137 -45198 -60133 -44902
rect -60133 -45198 -59517 -44902
rect -59517 -45198 -59513 -44902
rect -60137 -45202 -59513 -45198
rect -59477 -44902 -59173 -44898
rect -59477 -45198 -59473 -44902
rect -59473 -45198 -59177 -44902
rect -59177 -45198 -59173 -44902
rect -59477 -45202 -59173 -45198
rect -59137 -44902 -58513 -44898
rect -59137 -45198 -59133 -44902
rect -59133 -45198 -58517 -44902
rect -58517 -45198 -58513 -44902
rect -59137 -45202 -58513 -45198
rect -58477 -44902 -58173 -44898
rect -58477 -45198 -58473 -44902
rect -58473 -45198 -58177 -44902
rect -58177 -45198 -58173 -44902
rect -58477 -45202 -58173 -45198
rect -58137 -44902 -57513 -44898
rect -58137 -45198 -58133 -44902
rect -58133 -45198 -57517 -44902
rect -57517 -45198 -57513 -44902
rect -58137 -45202 -57513 -45198
rect -57477 -44902 -57173 -44898
rect -57477 -45198 -57473 -44902
rect -57473 -45198 -57177 -44902
rect -57177 -45198 -57173 -44902
rect -57477 -45202 -57173 -45198
rect -57137 -44902 -56513 -44898
rect -57137 -45198 -57133 -44902
rect -57133 -45198 -56517 -44902
rect -56517 -45198 -56513 -44902
rect -57137 -45202 -56513 -45198
rect -56477 -44902 -56173 -44898
rect -56477 -45198 -56473 -44902
rect -56473 -45198 -56177 -44902
rect -56177 -45198 -56173 -44902
rect -56477 -45202 -56173 -45198
rect -56137 -44902 -55513 -44898
rect -56137 -45198 -56133 -44902
rect -56133 -45198 -55517 -44902
rect -55517 -45198 -55513 -44902
rect -56137 -45202 -55513 -45198
rect -55477 -44902 -55173 -44898
rect -55477 -45198 -55473 -44902
rect -55473 -45198 -55177 -44902
rect -55177 -45198 -55173 -44902
rect -55477 -45202 -55173 -45198
rect -55137 -44902 -54513 -44898
rect -55137 -45198 -55133 -44902
rect -55133 -45198 -54517 -44902
rect -54517 -45198 -54513 -44902
rect -55137 -45202 -54513 -45198
rect -54477 -44902 -54173 -44898
rect -54477 -45198 -54473 -44902
rect -54473 -45198 -54177 -44902
rect -54177 -45198 -54173 -44902
rect -54477 -45202 -54173 -45198
rect -54137 -44902 -53513 -44898
rect -54137 -45198 -54133 -44902
rect -54133 -45198 -53517 -44902
rect -53517 -45198 -53513 -44902
rect -54137 -45202 -53513 -45198
rect -53477 -44902 -53173 -44898
rect -53477 -45198 -53473 -44902
rect -53473 -45198 -53177 -44902
rect -53177 -45198 -53173 -44902
rect -53477 -45202 -53173 -45198
rect -53137 -44902 -52513 -44898
rect -53137 -45198 -53133 -44902
rect -53133 -45198 -52517 -44902
rect -52517 -45198 -52513 -44902
rect -53137 -45202 -52513 -45198
rect -52477 -44902 -52173 -44898
rect -52477 -45198 -52473 -44902
rect -52473 -45198 -52177 -44902
rect -52177 -45198 -52173 -44902
rect -52477 -45202 -52173 -45198
rect -52137 -44902 -51513 -44898
rect -52137 -45198 -52133 -44902
rect -52133 -45198 -51517 -44902
rect -51517 -45198 -51513 -44902
rect -52137 -45202 -51513 -45198
rect -51477 -44902 -51173 -44898
rect -51477 -45198 -51473 -44902
rect -51473 -45198 -51177 -44902
rect -51177 -45198 -51173 -44902
rect -51477 -45202 -51173 -45198
rect -51137 -44902 -50513 -44898
rect -51137 -45198 -51133 -44902
rect -51133 -45198 -50517 -44902
rect -50517 -45198 -50513 -44902
rect -51137 -45202 -50513 -45198
rect -50477 -44902 -50173 -44898
rect -50477 -45198 -50473 -44902
rect -50473 -45198 -50177 -44902
rect -50177 -45198 -50173 -44902
rect -50477 -45202 -50173 -45198
rect -50137 -44902 -49513 -44898
rect -50137 -45198 -50133 -44902
rect -50133 -45198 -49517 -44902
rect -49517 -45198 -49513 -44902
rect -50137 -45202 -49513 -45198
rect -49477 -44902 -49173 -44898
rect -49477 -45198 -49473 -44902
rect -49473 -45198 -49177 -44902
rect -49177 -45198 -49173 -44902
rect -49477 -45202 -49173 -45198
rect -49137 -44902 -48833 -44898
rect -49137 -45198 -49133 -44902
rect -49133 -45198 -48837 -44902
rect -48837 -45198 -48833 -44902
rect -49137 -45202 -48833 -45198
rect 8283 -44902 8587 -44898
rect 8283 -45198 8287 -44902
rect 8287 -45198 8583 -44902
rect 8583 -45198 8587 -44902
rect 8283 -45202 8587 -45198
rect 8623 -44902 8927 -44898
rect 8623 -45198 8627 -44902
rect 8627 -45198 8923 -44902
rect 8923 -45198 8927 -44902
rect 8623 -45202 8927 -45198
rect 8963 -44902 9587 -44898
rect 8963 -45198 8967 -44902
rect 8967 -45198 9583 -44902
rect 9583 -45198 9587 -44902
rect 8963 -45202 9587 -45198
rect 9623 -44902 9927 -44898
rect 9623 -45198 9627 -44902
rect 9627 -45198 9923 -44902
rect 9923 -45198 9927 -44902
rect 9623 -45202 9927 -45198
rect 9963 -44902 10587 -44898
rect 9963 -45198 9967 -44902
rect 9967 -45198 10583 -44902
rect 10583 -45198 10587 -44902
rect 9963 -45202 10587 -45198
rect 10623 -44902 10927 -44898
rect 10623 -45198 10627 -44902
rect 10627 -45198 10923 -44902
rect 10923 -45198 10927 -44902
rect 10623 -45202 10927 -45198
rect 10963 -44902 11587 -44898
rect 10963 -45198 10967 -44902
rect 10967 -45198 11583 -44902
rect 11583 -45198 11587 -44902
rect 10963 -45202 11587 -45198
rect 11623 -44902 11927 -44898
rect 11623 -45198 11627 -44902
rect 11627 -45198 11923 -44902
rect 11923 -45198 11927 -44902
rect 11623 -45202 11927 -45198
rect 11963 -44902 12587 -44898
rect 11963 -45198 11967 -44902
rect 11967 -45198 12583 -44902
rect 12583 -45198 12587 -44902
rect 11963 -45202 12587 -45198
rect 12623 -44902 12927 -44898
rect 12623 -45198 12627 -44902
rect 12627 -45198 12923 -44902
rect 12923 -45198 12927 -44902
rect 12623 -45202 12927 -45198
rect 12963 -44902 13587 -44898
rect 12963 -45198 12967 -44902
rect 12967 -45198 13583 -44902
rect 13583 -45198 13587 -44902
rect 12963 -45202 13587 -45198
rect 13623 -44902 13927 -44898
rect 13623 -45198 13627 -44902
rect 13627 -45198 13923 -44902
rect 13923 -45198 13927 -44902
rect 13623 -45202 13927 -45198
rect 13963 -44902 14587 -44898
rect 13963 -45198 13967 -44902
rect 13967 -45198 14583 -44902
rect 14583 -45198 14587 -44902
rect 13963 -45202 14587 -45198
rect 14623 -44902 14927 -44898
rect 14623 -45198 14627 -44902
rect 14627 -45198 14923 -44902
rect 14923 -45198 14927 -44902
rect 14623 -45202 14927 -45198
rect 14963 -44902 15587 -44898
rect 14963 -45198 14967 -44902
rect 14967 -45198 15583 -44902
rect 15583 -45198 15587 -44902
rect 14963 -45202 15587 -45198
rect 15623 -44902 15927 -44898
rect 15623 -45198 15627 -44902
rect 15627 -45198 15923 -44902
rect 15923 -45198 15927 -44902
rect 15623 -45202 15927 -45198
rect 15963 -44902 16587 -44898
rect 15963 -45198 15967 -44902
rect 15967 -45198 16583 -44902
rect 16583 -45198 16587 -44902
rect 15963 -45202 16587 -45198
rect 16623 -44902 16927 -44898
rect 16623 -45198 16627 -44902
rect 16627 -45198 16923 -44902
rect 16923 -45198 16927 -44902
rect 16623 -45202 16927 -45198
rect 16963 -44902 17587 -44898
rect 16963 -45198 16967 -44902
rect 16967 -45198 17583 -44902
rect 17583 -45198 17587 -44902
rect 16963 -45202 17587 -45198
rect 17623 -44902 17927 -44898
rect 17623 -45198 17627 -44902
rect 17627 -45198 17923 -44902
rect 17923 -45198 17927 -44902
rect 17623 -45202 17927 -45198
rect 17963 -44902 18587 -44898
rect 17963 -45198 17967 -44902
rect 17967 -45198 18583 -44902
rect 18583 -45198 18587 -44902
rect 17963 -45202 18587 -45198
rect 18623 -44902 18927 -44898
rect 18623 -45198 18627 -44902
rect 18627 -45198 18923 -44902
rect 18923 -45198 18927 -44902
rect 18623 -45202 18927 -45198
rect 18963 -44902 19587 -44898
rect 18963 -45198 18967 -44902
rect 18967 -45198 19583 -44902
rect 19583 -45198 19587 -44902
rect 18963 -45202 19587 -45198
rect 19623 -44902 19927 -44898
rect 19623 -45198 19627 -44902
rect 19627 -45198 19923 -44902
rect 19923 -45198 19927 -44902
rect 19623 -45202 19927 -45198
rect 19963 -44902 20587 -44898
rect 19963 -45198 19967 -44902
rect 19967 -45198 20583 -44902
rect 20583 -45198 20587 -44902
rect 19963 -45202 20587 -45198
rect 20623 -44902 20927 -44898
rect 20623 -45198 20627 -44902
rect 20627 -45198 20923 -44902
rect 20923 -45198 20927 -44902
rect 20623 -45202 20927 -45198
rect 20963 -44902 21587 -44898
rect 20963 -45198 20967 -44902
rect 20967 -45198 21583 -44902
rect 21583 -45198 21587 -44902
rect 20963 -45202 21587 -45198
rect 21623 -44902 21927 -44898
rect 21623 -45198 21627 -44902
rect 21627 -45198 21923 -44902
rect 21923 -45198 21927 -44902
rect 21623 -45202 21927 -45198
rect 21963 -44902 22587 -44898
rect 21963 -45198 21967 -44902
rect 21967 -45198 22583 -44902
rect 22583 -45198 22587 -44902
rect 21963 -45202 22587 -45198
rect 22623 -44902 22927 -44898
rect 22623 -45198 22627 -44902
rect 22627 -45198 22923 -44902
rect 22923 -45198 22927 -44902
rect 22623 -45202 22927 -45198
rect 22963 -44902 23587 -44898
rect 22963 -45198 22967 -44902
rect 22967 -45198 23583 -44902
rect 23583 -45198 23587 -44902
rect 22963 -45202 23587 -45198
rect 23623 -44902 23927 -44898
rect 23623 -45198 23627 -44902
rect 23627 -45198 23923 -44902
rect 23923 -45198 23927 -44902
rect 23623 -45202 23927 -45198
rect 23963 -44902 24587 -44898
rect 23963 -45198 23967 -44902
rect 23967 -45198 24583 -44902
rect 24583 -45198 24587 -44902
rect 23963 -45202 24587 -45198
rect 24623 -44902 24927 -44898
rect 24623 -45198 24627 -44902
rect 24627 -45198 24923 -44902
rect 24923 -45198 24927 -44902
rect 24623 -45202 24927 -45198
rect 24963 -44902 25587 -44898
rect 24963 -45198 24967 -44902
rect 24967 -45198 25583 -44902
rect 25583 -45198 25587 -44902
rect 24963 -45202 25587 -45198
rect 25623 -44902 25927 -44898
rect 25623 -45198 25627 -44902
rect 25627 -45198 25923 -44902
rect 25923 -45198 25927 -44902
rect 25623 -45202 25927 -45198
rect 25963 -44902 26587 -44898
rect 25963 -45198 25967 -44902
rect 25967 -45198 26583 -44902
rect 26583 -45198 26587 -44902
rect 25963 -45202 26587 -45198
rect 26623 -44902 26927 -44898
rect 26623 -45198 26627 -44902
rect 26627 -45198 26923 -44902
rect 26923 -45198 26927 -44902
rect 26623 -45202 26927 -45198
rect 26963 -44902 27587 -44898
rect 26963 -45198 26967 -44902
rect 26967 -45198 27583 -44902
rect 27583 -45198 27587 -44902
rect 26963 -45202 27587 -45198
rect 27623 -44902 27927 -44898
rect 27623 -45198 27627 -44902
rect 27627 -45198 27923 -44902
rect 27923 -45198 27927 -44902
rect 27623 -45202 27927 -45198
rect 27963 -44902 28587 -44898
rect 27963 -45198 27967 -44902
rect 27967 -45198 28583 -44902
rect 28583 -45198 28587 -44902
rect 27963 -45202 28587 -45198
rect 28623 -44902 28927 -44898
rect 28623 -45198 28627 -44902
rect 28627 -45198 28923 -44902
rect 28923 -45198 28927 -44902
rect 28623 -45202 28927 -45198
rect 28963 -44902 29587 -44898
rect 28963 -45198 28967 -44902
rect 28967 -45198 29583 -44902
rect 29583 -45198 29587 -44902
rect 28963 -45202 29587 -45198
rect 29623 -44902 29927 -44898
rect 29623 -45198 29627 -44902
rect 29627 -45198 29923 -44902
rect 29923 -45198 29927 -44902
rect 29623 -45202 29927 -45198
rect 29963 -44902 30587 -44898
rect 29963 -45198 29967 -44902
rect 29967 -45198 30583 -44902
rect 30583 -45198 30587 -44902
rect 29963 -45202 30587 -45198
rect 30623 -44902 30927 -44898
rect 30623 -45198 30627 -44902
rect 30627 -45198 30923 -44902
rect 30923 -45198 30927 -44902
rect 30623 -45202 30927 -45198
rect 30963 -44902 31587 -44898
rect 30963 -45198 30967 -44902
rect 30967 -45198 31583 -44902
rect 31583 -45198 31587 -44902
rect 30963 -45202 31587 -45198
rect 31623 -44902 31927 -44898
rect 31623 -45198 31627 -44902
rect 31627 -45198 31923 -44902
rect 31923 -45198 31927 -44902
rect 31623 -45202 31927 -45198
rect 31963 -44902 32587 -44898
rect 31963 -45198 31967 -44902
rect 31967 -45198 32583 -44902
rect 32583 -45198 32587 -44902
rect 31963 -45202 32587 -45198
rect 32623 -44902 32927 -44898
rect 32623 -45198 32627 -44902
rect 32627 -45198 32923 -44902
rect 32923 -45198 32927 -44902
rect 32623 -45202 32927 -45198
rect 32963 -44902 33587 -44898
rect 32963 -45198 32967 -44902
rect 32967 -45198 33583 -44902
rect 33583 -45198 33587 -44902
rect 32963 -45202 33587 -45198
rect 33623 -44902 33927 -44898
rect 33623 -45198 33627 -44902
rect 33627 -45198 33923 -44902
rect 33923 -45198 33927 -44902
rect 33623 -45202 33927 -45198
rect 33963 -44902 34267 -44898
rect 33963 -45198 33967 -44902
rect 33967 -45198 34263 -44902
rect 34263 -45198 34267 -44902
rect 33963 -45202 34267 -45198
rect -74477 -45242 -74173 -45238
rect -74477 -45858 -74473 -45242
rect -74473 -45858 -74177 -45242
rect -74177 -45858 -74173 -45242
rect -74477 -45862 -74173 -45858
rect -73477 -45242 -73173 -45238
rect -73477 -45858 -73473 -45242
rect -73473 -45858 -73177 -45242
rect -73177 -45858 -73173 -45242
rect -73477 -45862 -73173 -45858
rect -72477 -45242 -72173 -45238
rect -72477 -45858 -72473 -45242
rect -72473 -45858 -72177 -45242
rect -72177 -45858 -72173 -45242
rect -72477 -45862 -72173 -45858
rect -71477 -45242 -71173 -45238
rect -71477 -45858 -71473 -45242
rect -71473 -45858 -71177 -45242
rect -71177 -45858 -71173 -45242
rect -71477 -45862 -71173 -45858
rect -70477 -45242 -70173 -45238
rect -70477 -45858 -70473 -45242
rect -70473 -45858 -70177 -45242
rect -70177 -45858 -70173 -45242
rect -70477 -45862 -70173 -45858
rect -69477 -45242 -69173 -45238
rect -69477 -45858 -69473 -45242
rect -69473 -45858 -69177 -45242
rect -69177 -45858 -69173 -45242
rect -69477 -45862 -69173 -45858
rect -68477 -45242 -68173 -45238
rect -68477 -45858 -68473 -45242
rect -68473 -45858 -68177 -45242
rect -68177 -45858 -68173 -45242
rect -68477 -45862 -68173 -45858
rect -67477 -45242 -67173 -45238
rect -67477 -45858 -67473 -45242
rect -67473 -45858 -67177 -45242
rect -67177 -45858 -67173 -45242
rect -67477 -45862 -67173 -45858
rect -66477 -45242 -66173 -45238
rect -66477 -45858 -66473 -45242
rect -66473 -45858 -66177 -45242
rect -66177 -45858 -66173 -45242
rect -66477 -45862 -66173 -45858
rect -65477 -45242 -65173 -45238
rect -65477 -45858 -65473 -45242
rect -65473 -45858 -65177 -45242
rect -65177 -45858 -65173 -45242
rect -65477 -45862 -65173 -45858
rect -64477 -45242 -64173 -45238
rect -64477 -45858 -64473 -45242
rect -64473 -45858 -64177 -45242
rect -64177 -45858 -64173 -45242
rect -64477 -45862 -64173 -45858
rect -63477 -45242 -63173 -45238
rect -63477 -45858 -63473 -45242
rect -63473 -45858 -63177 -45242
rect -63177 -45858 -63173 -45242
rect -63477 -45862 -63173 -45858
rect -62477 -45242 -62173 -45238
rect -62477 -45858 -62473 -45242
rect -62473 -45858 -62177 -45242
rect -62177 -45858 -62173 -45242
rect -62477 -45862 -62173 -45858
rect -61477 -45242 -61173 -45238
rect -61477 -45858 -61473 -45242
rect -61473 -45858 -61177 -45242
rect -61177 -45858 -61173 -45242
rect -61477 -45862 -61173 -45858
rect -60477 -45242 -60173 -45238
rect -60477 -45858 -60473 -45242
rect -60473 -45858 -60177 -45242
rect -60177 -45858 -60173 -45242
rect -60477 -45862 -60173 -45858
rect -59477 -45242 -59173 -45238
rect -59477 -45858 -59473 -45242
rect -59473 -45858 -59177 -45242
rect -59177 -45858 -59173 -45242
rect -59477 -45862 -59173 -45858
rect -58477 -45242 -58173 -45238
rect -58477 -45858 -58473 -45242
rect -58473 -45858 -58177 -45242
rect -58177 -45858 -58173 -45242
rect -58477 -45862 -58173 -45858
rect -57477 -45242 -57173 -45238
rect -57477 -45858 -57473 -45242
rect -57473 -45858 -57177 -45242
rect -57177 -45858 -57173 -45242
rect -57477 -45862 -57173 -45858
rect -56477 -45242 -56173 -45238
rect -56477 -45858 -56473 -45242
rect -56473 -45858 -56177 -45242
rect -56177 -45858 -56173 -45242
rect -56477 -45862 -56173 -45858
rect -55477 -45242 -55173 -45238
rect -55477 -45858 -55473 -45242
rect -55473 -45858 -55177 -45242
rect -55177 -45858 -55173 -45242
rect -55477 -45862 -55173 -45858
rect -54477 -45242 -54173 -45238
rect -54477 -45858 -54473 -45242
rect -54473 -45858 -54177 -45242
rect -54177 -45858 -54173 -45242
rect -54477 -45862 -54173 -45858
rect -53477 -45242 -53173 -45238
rect -53477 -45858 -53473 -45242
rect -53473 -45858 -53177 -45242
rect -53177 -45858 -53173 -45242
rect -53477 -45862 -53173 -45858
rect -52477 -45242 -52173 -45238
rect -52477 -45858 -52473 -45242
rect -52473 -45858 -52177 -45242
rect -52177 -45858 -52173 -45242
rect -52477 -45862 -52173 -45858
rect -51477 -45242 -51173 -45238
rect -51477 -45858 -51473 -45242
rect -51473 -45858 -51177 -45242
rect -51177 -45858 -51173 -45242
rect -51477 -45862 -51173 -45858
rect -50477 -45242 -50173 -45238
rect -50477 -45858 -50473 -45242
rect -50473 -45858 -50177 -45242
rect -50177 -45858 -50173 -45242
rect -50477 -45862 -50173 -45858
rect -49477 -45242 -49173 -45238
rect -49477 -45858 -49473 -45242
rect -49473 -45858 -49177 -45242
rect -49177 -45858 -49173 -45242
rect -49477 -45862 -49173 -45858
rect 8623 -45242 8927 -45238
rect 8623 -45858 8627 -45242
rect 8627 -45858 8923 -45242
rect 8923 -45858 8927 -45242
rect 8623 -45862 8927 -45858
rect 9623 -45242 9927 -45238
rect 9623 -45858 9627 -45242
rect 9627 -45858 9923 -45242
rect 9923 -45858 9927 -45242
rect 9623 -45862 9927 -45858
rect 10623 -45242 10927 -45238
rect 10623 -45858 10627 -45242
rect 10627 -45858 10923 -45242
rect 10923 -45858 10927 -45242
rect 10623 -45862 10927 -45858
rect 11623 -45242 11927 -45238
rect 11623 -45858 11627 -45242
rect 11627 -45858 11923 -45242
rect 11923 -45858 11927 -45242
rect 11623 -45862 11927 -45858
rect 12623 -45242 12927 -45238
rect 12623 -45858 12627 -45242
rect 12627 -45858 12923 -45242
rect 12923 -45858 12927 -45242
rect 12623 -45862 12927 -45858
rect 13623 -45242 13927 -45238
rect 13623 -45858 13627 -45242
rect 13627 -45858 13923 -45242
rect 13923 -45858 13927 -45242
rect 13623 -45862 13927 -45858
rect 14623 -45242 14927 -45238
rect 14623 -45858 14627 -45242
rect 14627 -45858 14923 -45242
rect 14923 -45858 14927 -45242
rect 14623 -45862 14927 -45858
rect 15623 -45242 15927 -45238
rect 15623 -45858 15627 -45242
rect 15627 -45858 15923 -45242
rect 15923 -45858 15927 -45242
rect 15623 -45862 15927 -45858
rect 16623 -45242 16927 -45238
rect 16623 -45858 16627 -45242
rect 16627 -45858 16923 -45242
rect 16923 -45858 16927 -45242
rect 16623 -45862 16927 -45858
rect 17623 -45242 17927 -45238
rect 17623 -45858 17627 -45242
rect 17627 -45858 17923 -45242
rect 17923 -45858 17927 -45242
rect 17623 -45862 17927 -45858
rect 18623 -45242 18927 -45238
rect 18623 -45858 18627 -45242
rect 18627 -45858 18923 -45242
rect 18923 -45858 18927 -45242
rect 18623 -45862 18927 -45858
rect 19623 -45242 19927 -45238
rect 19623 -45858 19627 -45242
rect 19627 -45858 19923 -45242
rect 19923 -45858 19927 -45242
rect 19623 -45862 19927 -45858
rect 20623 -45242 20927 -45238
rect 20623 -45858 20627 -45242
rect 20627 -45858 20923 -45242
rect 20923 -45858 20927 -45242
rect 20623 -45862 20927 -45858
rect 21623 -45242 21927 -45238
rect 21623 -45858 21627 -45242
rect 21627 -45858 21923 -45242
rect 21923 -45858 21927 -45242
rect 21623 -45862 21927 -45858
rect 22623 -45242 22927 -45238
rect 22623 -45858 22627 -45242
rect 22627 -45858 22923 -45242
rect 22923 -45858 22927 -45242
rect 22623 -45862 22927 -45858
rect 23623 -45242 23927 -45238
rect 23623 -45858 23627 -45242
rect 23627 -45858 23923 -45242
rect 23923 -45858 23927 -45242
rect 23623 -45862 23927 -45858
rect 24623 -45242 24927 -45238
rect 24623 -45858 24627 -45242
rect 24627 -45858 24923 -45242
rect 24923 -45858 24927 -45242
rect 24623 -45862 24927 -45858
rect 25623 -45242 25927 -45238
rect 25623 -45858 25627 -45242
rect 25627 -45858 25923 -45242
rect 25923 -45858 25927 -45242
rect 25623 -45862 25927 -45858
rect 26623 -45242 26927 -45238
rect 26623 -45858 26627 -45242
rect 26627 -45858 26923 -45242
rect 26923 -45858 26927 -45242
rect 26623 -45862 26927 -45858
rect 27623 -45242 27927 -45238
rect 27623 -45858 27627 -45242
rect 27627 -45858 27923 -45242
rect 27923 -45858 27927 -45242
rect 27623 -45862 27927 -45858
rect 28623 -45242 28927 -45238
rect 28623 -45858 28627 -45242
rect 28627 -45858 28923 -45242
rect 28923 -45858 28927 -45242
rect 28623 -45862 28927 -45858
rect 29623 -45242 29927 -45238
rect 29623 -45858 29627 -45242
rect 29627 -45858 29923 -45242
rect 29923 -45858 29927 -45242
rect 29623 -45862 29927 -45858
rect 30623 -45242 30927 -45238
rect 30623 -45858 30627 -45242
rect 30627 -45858 30923 -45242
rect 30923 -45858 30927 -45242
rect 30623 -45862 30927 -45858
rect 31623 -45242 31927 -45238
rect 31623 -45858 31627 -45242
rect 31627 -45858 31923 -45242
rect 31923 -45858 31927 -45242
rect 31623 -45862 31927 -45858
rect 32623 -45242 32927 -45238
rect 32623 -45858 32627 -45242
rect 32627 -45858 32923 -45242
rect 32923 -45858 32927 -45242
rect 32623 -45862 32927 -45858
rect 33623 -45242 33927 -45238
rect 33623 -45858 33627 -45242
rect 33627 -45858 33923 -45242
rect 33923 -45858 33927 -45242
rect 33623 -45862 33927 -45858
rect -74817 -45902 -74513 -45898
rect -74817 -46198 -74813 -45902
rect -74813 -46198 -74517 -45902
rect -74517 -46198 -74513 -45902
rect -74817 -46202 -74513 -46198
rect -74477 -45902 -74173 -45898
rect -74477 -46198 -74473 -45902
rect -74473 -46198 -74177 -45902
rect -74177 -46198 -74173 -45902
rect -74477 -46202 -74173 -46198
rect -74137 -45902 -73513 -45898
rect -74137 -46198 -74133 -45902
rect -74133 -46198 -73517 -45902
rect -73517 -46198 -73513 -45902
rect -74137 -46202 -73513 -46198
rect -73477 -45902 -73173 -45898
rect -73477 -46198 -73473 -45902
rect -73473 -46198 -73177 -45902
rect -73177 -46198 -73173 -45902
rect -73477 -46202 -73173 -46198
rect -73137 -45902 -72513 -45898
rect -73137 -46198 -73133 -45902
rect -73133 -46198 -72517 -45902
rect -72517 -46198 -72513 -45902
rect -73137 -46202 -72513 -46198
rect -72477 -45902 -72173 -45898
rect -72477 -46198 -72473 -45902
rect -72473 -46198 -72177 -45902
rect -72177 -46198 -72173 -45902
rect -72477 -46202 -72173 -46198
rect -72137 -45902 -71513 -45898
rect -72137 -46198 -72133 -45902
rect -72133 -46198 -71517 -45902
rect -71517 -46198 -71513 -45902
rect -72137 -46202 -71513 -46198
rect -71477 -45902 -71173 -45898
rect -71477 -46198 -71473 -45902
rect -71473 -46198 -71177 -45902
rect -71177 -46198 -71173 -45902
rect -71477 -46202 -71173 -46198
rect -71137 -45902 -70513 -45898
rect -71137 -46198 -71133 -45902
rect -71133 -46198 -70517 -45902
rect -70517 -46198 -70513 -45902
rect -71137 -46202 -70513 -46198
rect -70477 -45902 -70173 -45898
rect -70477 -46198 -70473 -45902
rect -70473 -46198 -70177 -45902
rect -70177 -46198 -70173 -45902
rect -70477 -46202 -70173 -46198
rect -70137 -45902 -69513 -45898
rect -70137 -46198 -70133 -45902
rect -70133 -46198 -69517 -45902
rect -69517 -46198 -69513 -45902
rect -70137 -46202 -69513 -46198
rect -69477 -45902 -69173 -45898
rect -69477 -46198 -69473 -45902
rect -69473 -46198 -69177 -45902
rect -69177 -46198 -69173 -45902
rect -69477 -46202 -69173 -46198
rect -69137 -45902 -68513 -45898
rect -69137 -46198 -69133 -45902
rect -69133 -46198 -68517 -45902
rect -68517 -46198 -68513 -45902
rect -69137 -46202 -68513 -46198
rect -68477 -45902 -68173 -45898
rect -68477 -46198 -68473 -45902
rect -68473 -46198 -68177 -45902
rect -68177 -46198 -68173 -45902
rect -68477 -46202 -68173 -46198
rect -68137 -45902 -67513 -45898
rect -68137 -46198 -68133 -45902
rect -68133 -46198 -67517 -45902
rect -67517 -46198 -67513 -45902
rect -68137 -46202 -67513 -46198
rect -67477 -45902 -67173 -45898
rect -67477 -46198 -67473 -45902
rect -67473 -46198 -67177 -45902
rect -67177 -46198 -67173 -45902
rect -67477 -46202 -67173 -46198
rect -67137 -45902 -66513 -45898
rect -67137 -46198 -67133 -45902
rect -67133 -46198 -66517 -45902
rect -66517 -46198 -66513 -45902
rect -67137 -46202 -66513 -46198
rect -66477 -45902 -66173 -45898
rect -66477 -46198 -66473 -45902
rect -66473 -46198 -66177 -45902
rect -66177 -46198 -66173 -45902
rect -66477 -46202 -66173 -46198
rect -66137 -45902 -65513 -45898
rect -66137 -46198 -66133 -45902
rect -66133 -46198 -65517 -45902
rect -65517 -46198 -65513 -45902
rect -66137 -46202 -65513 -46198
rect -65477 -45902 -65173 -45898
rect -65477 -46198 -65473 -45902
rect -65473 -46198 -65177 -45902
rect -65177 -46198 -65173 -45902
rect -65477 -46202 -65173 -46198
rect -65137 -45902 -64513 -45898
rect -65137 -46198 -65133 -45902
rect -65133 -46198 -64517 -45902
rect -64517 -46198 -64513 -45902
rect -65137 -46202 -64513 -46198
rect -64477 -45902 -64173 -45898
rect -64477 -46198 -64473 -45902
rect -64473 -46198 -64177 -45902
rect -64177 -46198 -64173 -45902
rect -64477 -46202 -64173 -46198
rect -64137 -45902 -63513 -45898
rect -64137 -46198 -64133 -45902
rect -64133 -46198 -63517 -45902
rect -63517 -46198 -63513 -45902
rect -64137 -46202 -63513 -46198
rect -63477 -45902 -63173 -45898
rect -63477 -46198 -63473 -45902
rect -63473 -46198 -63177 -45902
rect -63177 -46198 -63173 -45902
rect -63477 -46202 -63173 -46198
rect -63137 -45902 -62513 -45898
rect -63137 -46198 -63133 -45902
rect -63133 -46198 -62517 -45902
rect -62517 -46198 -62513 -45902
rect -63137 -46202 -62513 -46198
rect -62477 -45902 -62173 -45898
rect -62477 -46198 -62473 -45902
rect -62473 -46198 -62177 -45902
rect -62177 -46198 -62173 -45902
rect -62477 -46202 -62173 -46198
rect -62137 -45902 -61513 -45898
rect -62137 -46198 -62133 -45902
rect -62133 -46198 -61517 -45902
rect -61517 -46198 -61513 -45902
rect -62137 -46202 -61513 -46198
rect -61477 -45902 -61173 -45898
rect -61477 -46198 -61473 -45902
rect -61473 -46198 -61177 -45902
rect -61177 -46198 -61173 -45902
rect -61477 -46202 -61173 -46198
rect -61137 -45902 -60513 -45898
rect -61137 -46198 -61133 -45902
rect -61133 -46198 -60517 -45902
rect -60517 -46198 -60513 -45902
rect -61137 -46202 -60513 -46198
rect -60477 -45902 -60173 -45898
rect -60477 -46198 -60473 -45902
rect -60473 -46198 -60177 -45902
rect -60177 -46198 -60173 -45902
rect -60477 -46202 -60173 -46198
rect -60137 -45902 -59513 -45898
rect -60137 -46198 -60133 -45902
rect -60133 -46198 -59517 -45902
rect -59517 -46198 -59513 -45902
rect -60137 -46202 -59513 -46198
rect -59477 -45902 -59173 -45898
rect -59477 -46198 -59473 -45902
rect -59473 -46198 -59177 -45902
rect -59177 -46198 -59173 -45902
rect -59477 -46202 -59173 -46198
rect -59137 -45902 -58513 -45898
rect -59137 -46198 -59133 -45902
rect -59133 -46198 -58517 -45902
rect -58517 -46198 -58513 -45902
rect -59137 -46202 -58513 -46198
rect -58477 -45902 -58173 -45898
rect -58477 -46198 -58473 -45902
rect -58473 -46198 -58177 -45902
rect -58177 -46198 -58173 -45902
rect -58477 -46202 -58173 -46198
rect -58137 -45902 -57513 -45898
rect -58137 -46198 -58133 -45902
rect -58133 -46198 -57517 -45902
rect -57517 -46198 -57513 -45902
rect -58137 -46202 -57513 -46198
rect -57477 -45902 -57173 -45898
rect -57477 -46198 -57473 -45902
rect -57473 -46198 -57177 -45902
rect -57177 -46198 -57173 -45902
rect -57477 -46202 -57173 -46198
rect -57137 -45902 -56513 -45898
rect -57137 -46198 -57133 -45902
rect -57133 -46198 -56517 -45902
rect -56517 -46198 -56513 -45902
rect -57137 -46202 -56513 -46198
rect -56477 -45902 -56173 -45898
rect -56477 -46198 -56473 -45902
rect -56473 -46198 -56177 -45902
rect -56177 -46198 -56173 -45902
rect -56477 -46202 -56173 -46198
rect -56137 -45902 -55513 -45898
rect -56137 -46198 -56133 -45902
rect -56133 -46198 -55517 -45902
rect -55517 -46198 -55513 -45902
rect -56137 -46202 -55513 -46198
rect -55477 -45902 -55173 -45898
rect -55477 -46198 -55473 -45902
rect -55473 -46198 -55177 -45902
rect -55177 -46198 -55173 -45902
rect -55477 -46202 -55173 -46198
rect -55137 -45902 -54513 -45898
rect -55137 -46198 -55133 -45902
rect -55133 -46198 -54517 -45902
rect -54517 -46198 -54513 -45902
rect -55137 -46202 -54513 -46198
rect -54477 -45902 -54173 -45898
rect -54477 -46198 -54473 -45902
rect -54473 -46198 -54177 -45902
rect -54177 -46198 -54173 -45902
rect -54477 -46202 -54173 -46198
rect -54137 -45902 -53513 -45898
rect -54137 -46198 -54133 -45902
rect -54133 -46198 -53517 -45902
rect -53517 -46198 -53513 -45902
rect -54137 -46202 -53513 -46198
rect -53477 -45902 -53173 -45898
rect -53477 -46198 -53473 -45902
rect -53473 -46198 -53177 -45902
rect -53177 -46198 -53173 -45902
rect -53477 -46202 -53173 -46198
rect -53137 -45902 -52513 -45898
rect -53137 -46198 -53133 -45902
rect -53133 -46198 -52517 -45902
rect -52517 -46198 -52513 -45902
rect -53137 -46202 -52513 -46198
rect -52477 -45902 -52173 -45898
rect -52477 -46198 -52473 -45902
rect -52473 -46198 -52177 -45902
rect -52177 -46198 -52173 -45902
rect -52477 -46202 -52173 -46198
rect -52137 -45902 -51513 -45898
rect -52137 -46198 -52133 -45902
rect -52133 -46198 -51517 -45902
rect -51517 -46198 -51513 -45902
rect -52137 -46202 -51513 -46198
rect -51477 -45902 -51173 -45898
rect -51477 -46198 -51473 -45902
rect -51473 -46198 -51177 -45902
rect -51177 -46198 -51173 -45902
rect -51477 -46202 -51173 -46198
rect -51137 -45902 -50513 -45898
rect -51137 -46198 -51133 -45902
rect -51133 -46198 -50517 -45902
rect -50517 -46198 -50513 -45902
rect -51137 -46202 -50513 -46198
rect -50477 -45902 -50173 -45898
rect -50477 -46198 -50473 -45902
rect -50473 -46198 -50177 -45902
rect -50177 -46198 -50173 -45902
rect -50477 -46202 -50173 -46198
rect -50137 -45902 -49513 -45898
rect -50137 -46198 -50133 -45902
rect -50133 -46198 -49517 -45902
rect -49517 -46198 -49513 -45902
rect -50137 -46202 -49513 -46198
rect -49477 -45902 -49173 -45898
rect -49477 -46198 -49473 -45902
rect -49473 -46198 -49177 -45902
rect -49177 -46198 -49173 -45902
rect -49477 -46202 -49173 -46198
rect -49137 -45902 -48833 -45898
rect -49137 -46198 -49133 -45902
rect -49133 -46198 -48837 -45902
rect -48837 -46198 -48833 -45902
rect -49137 -46202 -48833 -46198
rect 8283 -45902 8587 -45898
rect 8283 -46198 8287 -45902
rect 8287 -46198 8583 -45902
rect 8583 -46198 8587 -45902
rect 8283 -46202 8587 -46198
rect 8623 -45902 8927 -45898
rect 8623 -46198 8627 -45902
rect 8627 -46198 8923 -45902
rect 8923 -46198 8927 -45902
rect 8623 -46202 8927 -46198
rect 8963 -45902 9587 -45898
rect 8963 -46198 8967 -45902
rect 8967 -46198 9583 -45902
rect 9583 -46198 9587 -45902
rect 8963 -46202 9587 -46198
rect 9623 -45902 9927 -45898
rect 9623 -46198 9627 -45902
rect 9627 -46198 9923 -45902
rect 9923 -46198 9927 -45902
rect 9623 -46202 9927 -46198
rect 9963 -45902 10587 -45898
rect 9963 -46198 9967 -45902
rect 9967 -46198 10583 -45902
rect 10583 -46198 10587 -45902
rect 9963 -46202 10587 -46198
rect 10623 -45902 10927 -45898
rect 10623 -46198 10627 -45902
rect 10627 -46198 10923 -45902
rect 10923 -46198 10927 -45902
rect 10623 -46202 10927 -46198
rect 10963 -45902 11587 -45898
rect 10963 -46198 10967 -45902
rect 10967 -46198 11583 -45902
rect 11583 -46198 11587 -45902
rect 10963 -46202 11587 -46198
rect 11623 -45902 11927 -45898
rect 11623 -46198 11627 -45902
rect 11627 -46198 11923 -45902
rect 11923 -46198 11927 -45902
rect 11623 -46202 11927 -46198
rect 11963 -45902 12587 -45898
rect 11963 -46198 11967 -45902
rect 11967 -46198 12583 -45902
rect 12583 -46198 12587 -45902
rect 11963 -46202 12587 -46198
rect 12623 -45902 12927 -45898
rect 12623 -46198 12627 -45902
rect 12627 -46198 12923 -45902
rect 12923 -46198 12927 -45902
rect 12623 -46202 12927 -46198
rect 12963 -45902 13587 -45898
rect 12963 -46198 12967 -45902
rect 12967 -46198 13583 -45902
rect 13583 -46198 13587 -45902
rect 12963 -46202 13587 -46198
rect 13623 -45902 13927 -45898
rect 13623 -46198 13627 -45902
rect 13627 -46198 13923 -45902
rect 13923 -46198 13927 -45902
rect 13623 -46202 13927 -46198
rect 13963 -45902 14587 -45898
rect 13963 -46198 13967 -45902
rect 13967 -46198 14583 -45902
rect 14583 -46198 14587 -45902
rect 13963 -46202 14587 -46198
rect 14623 -45902 14927 -45898
rect 14623 -46198 14627 -45902
rect 14627 -46198 14923 -45902
rect 14923 -46198 14927 -45902
rect 14623 -46202 14927 -46198
rect 14963 -45902 15587 -45898
rect 14963 -46198 14967 -45902
rect 14967 -46198 15583 -45902
rect 15583 -46198 15587 -45902
rect 14963 -46202 15587 -46198
rect 15623 -45902 15927 -45898
rect 15623 -46198 15627 -45902
rect 15627 -46198 15923 -45902
rect 15923 -46198 15927 -45902
rect 15623 -46202 15927 -46198
rect 15963 -45902 16587 -45898
rect 15963 -46198 15967 -45902
rect 15967 -46198 16583 -45902
rect 16583 -46198 16587 -45902
rect 15963 -46202 16587 -46198
rect 16623 -45902 16927 -45898
rect 16623 -46198 16627 -45902
rect 16627 -46198 16923 -45902
rect 16923 -46198 16927 -45902
rect 16623 -46202 16927 -46198
rect 16963 -45902 17587 -45898
rect 16963 -46198 16967 -45902
rect 16967 -46198 17583 -45902
rect 17583 -46198 17587 -45902
rect 16963 -46202 17587 -46198
rect 17623 -45902 17927 -45898
rect 17623 -46198 17627 -45902
rect 17627 -46198 17923 -45902
rect 17923 -46198 17927 -45902
rect 17623 -46202 17927 -46198
rect 17963 -45902 18587 -45898
rect 17963 -46198 17967 -45902
rect 17967 -46198 18583 -45902
rect 18583 -46198 18587 -45902
rect 17963 -46202 18587 -46198
rect 18623 -45902 18927 -45898
rect 18623 -46198 18627 -45902
rect 18627 -46198 18923 -45902
rect 18923 -46198 18927 -45902
rect 18623 -46202 18927 -46198
rect 18963 -45902 19587 -45898
rect 18963 -46198 18967 -45902
rect 18967 -46198 19583 -45902
rect 19583 -46198 19587 -45902
rect 18963 -46202 19587 -46198
rect 19623 -45902 19927 -45898
rect 19623 -46198 19627 -45902
rect 19627 -46198 19923 -45902
rect 19923 -46198 19927 -45902
rect 19623 -46202 19927 -46198
rect 19963 -45902 20587 -45898
rect 19963 -46198 19967 -45902
rect 19967 -46198 20583 -45902
rect 20583 -46198 20587 -45902
rect 19963 -46202 20587 -46198
rect 20623 -45902 20927 -45898
rect 20623 -46198 20627 -45902
rect 20627 -46198 20923 -45902
rect 20923 -46198 20927 -45902
rect 20623 -46202 20927 -46198
rect 20963 -45902 21587 -45898
rect 20963 -46198 20967 -45902
rect 20967 -46198 21583 -45902
rect 21583 -46198 21587 -45902
rect 20963 -46202 21587 -46198
rect 21623 -45902 21927 -45898
rect 21623 -46198 21627 -45902
rect 21627 -46198 21923 -45902
rect 21923 -46198 21927 -45902
rect 21623 -46202 21927 -46198
rect 21963 -45902 22587 -45898
rect 21963 -46198 21967 -45902
rect 21967 -46198 22583 -45902
rect 22583 -46198 22587 -45902
rect 21963 -46202 22587 -46198
rect 22623 -45902 22927 -45898
rect 22623 -46198 22627 -45902
rect 22627 -46198 22923 -45902
rect 22923 -46198 22927 -45902
rect 22623 -46202 22927 -46198
rect 22963 -45902 23587 -45898
rect 22963 -46198 22967 -45902
rect 22967 -46198 23583 -45902
rect 23583 -46198 23587 -45902
rect 22963 -46202 23587 -46198
rect 23623 -45902 23927 -45898
rect 23623 -46198 23627 -45902
rect 23627 -46198 23923 -45902
rect 23923 -46198 23927 -45902
rect 23623 -46202 23927 -46198
rect 23963 -45902 24587 -45898
rect 23963 -46198 23967 -45902
rect 23967 -46198 24583 -45902
rect 24583 -46198 24587 -45902
rect 23963 -46202 24587 -46198
rect 24623 -45902 24927 -45898
rect 24623 -46198 24627 -45902
rect 24627 -46198 24923 -45902
rect 24923 -46198 24927 -45902
rect 24623 -46202 24927 -46198
rect 24963 -45902 25587 -45898
rect 24963 -46198 24967 -45902
rect 24967 -46198 25583 -45902
rect 25583 -46198 25587 -45902
rect 24963 -46202 25587 -46198
rect 25623 -45902 25927 -45898
rect 25623 -46198 25627 -45902
rect 25627 -46198 25923 -45902
rect 25923 -46198 25927 -45902
rect 25623 -46202 25927 -46198
rect 25963 -45902 26587 -45898
rect 25963 -46198 25967 -45902
rect 25967 -46198 26583 -45902
rect 26583 -46198 26587 -45902
rect 25963 -46202 26587 -46198
rect 26623 -45902 26927 -45898
rect 26623 -46198 26627 -45902
rect 26627 -46198 26923 -45902
rect 26923 -46198 26927 -45902
rect 26623 -46202 26927 -46198
rect 26963 -45902 27587 -45898
rect 26963 -46198 26967 -45902
rect 26967 -46198 27583 -45902
rect 27583 -46198 27587 -45902
rect 26963 -46202 27587 -46198
rect 27623 -45902 27927 -45898
rect 27623 -46198 27627 -45902
rect 27627 -46198 27923 -45902
rect 27923 -46198 27927 -45902
rect 27623 -46202 27927 -46198
rect 27963 -45902 28587 -45898
rect 27963 -46198 27967 -45902
rect 27967 -46198 28583 -45902
rect 28583 -46198 28587 -45902
rect 27963 -46202 28587 -46198
rect 28623 -45902 28927 -45898
rect 28623 -46198 28627 -45902
rect 28627 -46198 28923 -45902
rect 28923 -46198 28927 -45902
rect 28623 -46202 28927 -46198
rect 28963 -45902 29587 -45898
rect 28963 -46198 28967 -45902
rect 28967 -46198 29583 -45902
rect 29583 -46198 29587 -45902
rect 28963 -46202 29587 -46198
rect 29623 -45902 29927 -45898
rect 29623 -46198 29627 -45902
rect 29627 -46198 29923 -45902
rect 29923 -46198 29927 -45902
rect 29623 -46202 29927 -46198
rect 29963 -45902 30587 -45898
rect 29963 -46198 29967 -45902
rect 29967 -46198 30583 -45902
rect 30583 -46198 30587 -45902
rect 29963 -46202 30587 -46198
rect 30623 -45902 30927 -45898
rect 30623 -46198 30627 -45902
rect 30627 -46198 30923 -45902
rect 30923 -46198 30927 -45902
rect 30623 -46202 30927 -46198
rect 30963 -45902 31587 -45898
rect 30963 -46198 30967 -45902
rect 30967 -46198 31583 -45902
rect 31583 -46198 31587 -45902
rect 30963 -46202 31587 -46198
rect 31623 -45902 31927 -45898
rect 31623 -46198 31627 -45902
rect 31627 -46198 31923 -45902
rect 31923 -46198 31927 -45902
rect 31623 -46202 31927 -46198
rect 31963 -45902 32587 -45898
rect 31963 -46198 31967 -45902
rect 31967 -46198 32583 -45902
rect 32583 -46198 32587 -45902
rect 31963 -46202 32587 -46198
rect 32623 -45902 32927 -45898
rect 32623 -46198 32627 -45902
rect 32627 -46198 32923 -45902
rect 32923 -46198 32927 -45902
rect 32623 -46202 32927 -46198
rect 32963 -45902 33587 -45898
rect 32963 -46198 32967 -45902
rect 32967 -46198 33583 -45902
rect 33583 -46198 33587 -45902
rect 32963 -46202 33587 -46198
rect 33623 -45902 33927 -45898
rect 33623 -46198 33627 -45902
rect 33627 -46198 33923 -45902
rect 33923 -46198 33927 -45902
rect 33623 -46202 33927 -46198
rect 33963 -45902 34267 -45898
rect 33963 -46198 33967 -45902
rect 33967 -46198 34263 -45902
rect 34263 -46198 34267 -45902
rect 33963 -46202 34267 -46198
rect -74477 -46242 -74173 -46238
rect -74477 -46538 -74473 -46242
rect -74473 -46538 -74177 -46242
rect -74177 -46538 -74173 -46242
rect -74477 -46542 -74173 -46538
rect -73477 -46242 -73173 -46238
rect -73477 -46538 -73473 -46242
rect -73473 -46538 -73177 -46242
rect -73177 -46538 -73173 -46242
rect -73477 -46542 -73173 -46538
rect -72477 -46242 -72173 -46238
rect -72477 -46538 -72473 -46242
rect -72473 -46538 -72177 -46242
rect -72177 -46538 -72173 -46242
rect -72477 -46542 -72173 -46538
rect -71477 -46242 -71173 -46238
rect -71477 -46538 -71473 -46242
rect -71473 -46538 -71177 -46242
rect -71177 -46538 -71173 -46242
rect -71477 -46542 -71173 -46538
rect -70477 -46242 -70173 -46238
rect -70477 -46538 -70473 -46242
rect -70473 -46538 -70177 -46242
rect -70177 -46538 -70173 -46242
rect -70477 -46542 -70173 -46538
rect -69477 -46242 -69173 -46238
rect -69477 -46538 -69473 -46242
rect -69473 -46538 -69177 -46242
rect -69177 -46538 -69173 -46242
rect -69477 -46542 -69173 -46538
rect -68477 -46242 -68173 -46238
rect -68477 -46538 -68473 -46242
rect -68473 -46538 -68177 -46242
rect -68177 -46538 -68173 -46242
rect -68477 -46542 -68173 -46538
rect -67477 -46242 -67173 -46238
rect -67477 -46538 -67473 -46242
rect -67473 -46538 -67177 -46242
rect -67177 -46538 -67173 -46242
rect -67477 -46542 -67173 -46538
rect -66477 -46242 -66173 -46238
rect -66477 -46538 -66473 -46242
rect -66473 -46538 -66177 -46242
rect -66177 -46538 -66173 -46242
rect -66477 -46542 -66173 -46538
rect -65477 -46242 -65173 -46238
rect -65477 -46538 -65473 -46242
rect -65473 -46538 -65177 -46242
rect -65177 -46538 -65173 -46242
rect -65477 -46542 -65173 -46538
rect -64477 -46242 -64173 -46238
rect -64477 -46538 -64473 -46242
rect -64473 -46538 -64177 -46242
rect -64177 -46538 -64173 -46242
rect -64477 -46542 -64173 -46538
rect -63477 -46242 -63173 -46238
rect -63477 -46538 -63473 -46242
rect -63473 -46538 -63177 -46242
rect -63177 -46538 -63173 -46242
rect -63477 -46542 -63173 -46538
rect -62477 -46242 -62173 -46238
rect -62477 -46538 -62473 -46242
rect -62473 -46538 -62177 -46242
rect -62177 -46538 -62173 -46242
rect -62477 -46542 -62173 -46538
rect -61477 -46242 -61173 -46238
rect -61477 -46538 -61473 -46242
rect -61473 -46538 -61177 -46242
rect -61177 -46538 -61173 -46242
rect -61477 -46542 -61173 -46538
rect -60477 -46242 -60173 -46238
rect -60477 -46538 -60473 -46242
rect -60473 -46538 -60177 -46242
rect -60177 -46538 -60173 -46242
rect -60477 -46542 -60173 -46538
rect -59477 -46242 -59173 -46238
rect -59477 -46538 -59473 -46242
rect -59473 -46538 -59177 -46242
rect -59177 -46538 -59173 -46242
rect -59477 -46542 -59173 -46538
rect -58477 -46242 -58173 -46238
rect -58477 -46538 -58473 -46242
rect -58473 -46538 -58177 -46242
rect -58177 -46538 -58173 -46242
rect -58477 -46542 -58173 -46538
rect -57477 -46242 -57173 -46238
rect -57477 -46538 -57473 -46242
rect -57473 -46538 -57177 -46242
rect -57177 -46538 -57173 -46242
rect -57477 -46542 -57173 -46538
rect -56477 -46242 -56173 -46238
rect -56477 -46538 -56473 -46242
rect -56473 -46538 -56177 -46242
rect -56177 -46538 -56173 -46242
rect -56477 -46542 -56173 -46538
rect -55477 -46242 -55173 -46238
rect -55477 -46538 -55473 -46242
rect -55473 -46538 -55177 -46242
rect -55177 -46538 -55173 -46242
rect -55477 -46542 -55173 -46538
rect -54477 -46242 -54173 -46238
rect -54477 -46538 -54473 -46242
rect -54473 -46538 -54177 -46242
rect -54177 -46538 -54173 -46242
rect -54477 -46542 -54173 -46538
rect -53477 -46242 -53173 -46238
rect -53477 -46538 -53473 -46242
rect -53473 -46538 -53177 -46242
rect -53177 -46538 -53173 -46242
rect -53477 -46542 -53173 -46538
rect -52477 -46242 -52173 -46238
rect -52477 -46538 -52473 -46242
rect -52473 -46538 -52177 -46242
rect -52177 -46538 -52173 -46242
rect -52477 -46542 -52173 -46538
rect -51477 -46242 -51173 -46238
rect -51477 -46538 -51473 -46242
rect -51473 -46538 -51177 -46242
rect -51177 -46538 -51173 -46242
rect -51477 -46542 -51173 -46538
rect -50477 -46242 -50173 -46238
rect -50477 -46538 -50473 -46242
rect -50473 -46538 -50177 -46242
rect -50177 -46538 -50173 -46242
rect -50477 -46542 -50173 -46538
rect -49477 -46242 -49173 -46238
rect -49477 -46538 -49473 -46242
rect -49473 -46538 -49177 -46242
rect -49177 -46538 -49173 -46242
rect -49477 -46542 -49173 -46538
rect 8623 -46242 8927 -46238
rect 8623 -46538 8627 -46242
rect 8627 -46538 8923 -46242
rect 8923 -46538 8927 -46242
rect 8623 -46542 8927 -46538
rect 9623 -46242 9927 -46238
rect 9623 -46538 9627 -46242
rect 9627 -46538 9923 -46242
rect 9923 -46538 9927 -46242
rect 9623 -46542 9927 -46538
rect 10623 -46242 10927 -46238
rect 10623 -46538 10627 -46242
rect 10627 -46538 10923 -46242
rect 10923 -46538 10927 -46242
rect 10623 -46542 10927 -46538
rect 11623 -46242 11927 -46238
rect 11623 -46538 11627 -46242
rect 11627 -46538 11923 -46242
rect 11923 -46538 11927 -46242
rect 11623 -46542 11927 -46538
rect 12623 -46242 12927 -46238
rect 12623 -46538 12627 -46242
rect 12627 -46538 12923 -46242
rect 12923 -46538 12927 -46242
rect 12623 -46542 12927 -46538
rect 13623 -46242 13927 -46238
rect 13623 -46538 13627 -46242
rect 13627 -46538 13923 -46242
rect 13923 -46538 13927 -46242
rect 13623 -46542 13927 -46538
rect 14623 -46242 14927 -46238
rect 14623 -46538 14627 -46242
rect 14627 -46538 14923 -46242
rect 14923 -46538 14927 -46242
rect 14623 -46542 14927 -46538
rect 15623 -46242 15927 -46238
rect 15623 -46538 15627 -46242
rect 15627 -46538 15923 -46242
rect 15923 -46538 15927 -46242
rect 15623 -46542 15927 -46538
rect 16623 -46242 16927 -46238
rect 16623 -46538 16627 -46242
rect 16627 -46538 16923 -46242
rect 16923 -46538 16927 -46242
rect 16623 -46542 16927 -46538
rect 17623 -46242 17927 -46238
rect 17623 -46538 17627 -46242
rect 17627 -46538 17923 -46242
rect 17923 -46538 17927 -46242
rect 17623 -46542 17927 -46538
rect 18623 -46242 18927 -46238
rect 18623 -46538 18627 -46242
rect 18627 -46538 18923 -46242
rect 18923 -46538 18927 -46242
rect 18623 -46542 18927 -46538
rect 19623 -46242 19927 -46238
rect 19623 -46538 19627 -46242
rect 19627 -46538 19923 -46242
rect 19923 -46538 19927 -46242
rect 19623 -46542 19927 -46538
rect 20623 -46242 20927 -46238
rect 20623 -46538 20627 -46242
rect 20627 -46538 20923 -46242
rect 20923 -46538 20927 -46242
rect 20623 -46542 20927 -46538
rect 21623 -46242 21927 -46238
rect 21623 -46538 21627 -46242
rect 21627 -46538 21923 -46242
rect 21923 -46538 21927 -46242
rect 21623 -46542 21927 -46538
rect 22623 -46242 22927 -46238
rect 22623 -46538 22627 -46242
rect 22627 -46538 22923 -46242
rect 22923 -46538 22927 -46242
rect 22623 -46542 22927 -46538
rect 23623 -46242 23927 -46238
rect 23623 -46538 23627 -46242
rect 23627 -46538 23923 -46242
rect 23923 -46538 23927 -46242
rect 23623 -46542 23927 -46538
rect 24623 -46242 24927 -46238
rect 24623 -46538 24627 -46242
rect 24627 -46538 24923 -46242
rect 24923 -46538 24927 -46242
rect 24623 -46542 24927 -46538
rect 25623 -46242 25927 -46238
rect 25623 -46538 25627 -46242
rect 25627 -46538 25923 -46242
rect 25923 -46538 25927 -46242
rect 25623 -46542 25927 -46538
rect 26623 -46242 26927 -46238
rect 26623 -46538 26627 -46242
rect 26627 -46538 26923 -46242
rect 26923 -46538 26927 -46242
rect 26623 -46542 26927 -46538
rect 27623 -46242 27927 -46238
rect 27623 -46538 27627 -46242
rect 27627 -46538 27923 -46242
rect 27923 -46538 27927 -46242
rect 27623 -46542 27927 -46538
rect 28623 -46242 28927 -46238
rect 28623 -46538 28627 -46242
rect 28627 -46538 28923 -46242
rect 28923 -46538 28927 -46242
rect 28623 -46542 28927 -46538
rect 29623 -46242 29927 -46238
rect 29623 -46538 29627 -46242
rect 29627 -46538 29923 -46242
rect 29923 -46538 29927 -46242
rect 29623 -46542 29927 -46538
rect 30623 -46242 30927 -46238
rect 30623 -46538 30627 -46242
rect 30627 -46538 30923 -46242
rect 30923 -46538 30927 -46242
rect 30623 -46542 30927 -46538
rect 31623 -46242 31927 -46238
rect 31623 -46538 31627 -46242
rect 31627 -46538 31923 -46242
rect 31923 -46538 31927 -46242
rect 31623 -46542 31927 -46538
rect 32623 -46242 32927 -46238
rect 32623 -46538 32627 -46242
rect 32627 -46538 32923 -46242
rect 32923 -46538 32927 -46242
rect 32623 -46542 32927 -46538
rect 33623 -46242 33927 -46238
rect 33623 -46538 33627 -46242
rect 33627 -46538 33923 -46242
rect 33923 -46538 33927 -46242
rect 33623 -46542 33927 -46538
<< metal4 >>
rect -74485 38542 -74165 38550
rect -74485 38238 -74477 38542
rect -74173 38238 -74165 38542
rect -74485 38210 -74165 38238
rect -73485 38542 -73165 38550
rect -73485 38238 -73477 38542
rect -73173 38238 -73165 38542
rect -73485 38210 -73165 38238
rect -72485 38542 -72165 38550
rect -72485 38238 -72477 38542
rect -72173 38238 -72165 38542
rect -72485 38210 -72165 38238
rect -71485 38542 -71165 38550
rect -71485 38238 -71477 38542
rect -71173 38238 -71165 38542
rect -71485 38210 -71165 38238
rect -70485 38542 -70165 38550
rect -70485 38238 -70477 38542
rect -70173 38238 -70165 38542
rect -70485 38210 -70165 38238
rect -69485 38542 -69165 38550
rect -69485 38238 -69477 38542
rect -69173 38238 -69165 38542
rect -69485 38210 -69165 38238
rect -68485 38542 -68165 38550
rect -68485 38238 -68477 38542
rect -68173 38238 -68165 38542
rect -68485 38210 -68165 38238
rect -67485 38542 -67165 38550
rect -67485 38238 -67477 38542
rect -67173 38238 -67165 38542
rect -67485 38210 -67165 38238
rect -66485 38542 -66165 38550
rect -66485 38238 -66477 38542
rect -66173 38238 -66165 38542
rect -66485 38210 -66165 38238
rect -65485 38542 -65165 38550
rect -65485 38238 -65477 38542
rect -65173 38238 -65165 38542
rect -65485 38210 -65165 38238
rect -64485 38542 -64165 38550
rect -64485 38238 -64477 38542
rect -64173 38238 -64165 38542
rect -64485 38210 -64165 38238
rect -63485 38542 -63165 38550
rect -63485 38238 -63477 38542
rect -63173 38238 -63165 38542
rect -63485 38210 -63165 38238
rect -62485 38542 -62165 38550
rect -62485 38238 -62477 38542
rect -62173 38238 -62165 38542
rect -62485 38210 -62165 38238
rect -61485 38542 -61165 38550
rect -61485 38238 -61477 38542
rect -61173 38238 -61165 38542
rect -61485 38210 -61165 38238
rect -60485 38542 -60165 38550
rect -60485 38238 -60477 38542
rect -60173 38238 -60165 38542
rect -60485 38210 -60165 38238
rect -59485 38542 -59165 38550
rect -59485 38238 -59477 38542
rect -59173 38238 -59165 38542
rect -59485 38210 -59165 38238
rect 9994 38542 10314 38550
rect 9994 38238 10002 38542
rect 10306 38238 10314 38542
rect 9994 38210 10314 38238
rect 10994 38542 11314 38550
rect 10994 38238 11002 38542
rect 11306 38238 11314 38542
rect 10994 38210 11314 38238
rect 11994 38542 12314 38550
rect 11994 38238 12002 38542
rect 12306 38238 12314 38542
rect 11994 38210 12314 38238
rect 12994 38542 13314 38550
rect 12994 38238 13002 38542
rect 13306 38238 13314 38542
rect 12994 38210 13314 38238
rect 13994 38542 14314 38550
rect 13994 38238 14002 38542
rect 14306 38238 14314 38542
rect 13994 38210 14314 38238
rect 14994 38542 15314 38550
rect 14994 38238 15002 38542
rect 15306 38238 15314 38542
rect 14994 38210 15314 38238
rect 15994 38542 16314 38550
rect 15994 38238 16002 38542
rect 16306 38238 16314 38542
rect 15994 38210 16314 38238
rect 16994 38542 17314 38550
rect 16994 38238 17002 38542
rect 17306 38238 17314 38542
rect 16994 38210 17314 38238
rect 17994 38542 18314 38550
rect 17994 38238 18002 38542
rect 18306 38238 18314 38542
rect 17994 38210 18314 38238
rect 18994 38542 19314 38550
rect 18994 38238 19002 38542
rect 19306 38238 19314 38542
rect 18994 38210 19314 38238
rect 19994 38542 20314 38550
rect 19994 38238 20002 38542
rect 20306 38238 20314 38542
rect 19994 38210 20314 38238
rect 20994 38542 21314 38550
rect 20994 38238 21002 38542
rect 21306 38238 21314 38542
rect 20994 38210 21314 38238
rect 21994 38542 22314 38550
rect 21994 38238 22002 38542
rect 22306 38238 22314 38542
rect 21994 38210 22314 38238
rect 22994 38542 23314 38550
rect 22994 38238 23002 38542
rect 23306 38238 23314 38542
rect 22994 38210 23314 38238
rect 23994 38542 24314 38550
rect 23994 38238 24002 38542
rect 24306 38238 24314 38542
rect 23994 38210 24314 38238
rect 24994 38542 25314 38550
rect 24994 38238 25002 38542
rect 25306 38238 25314 38542
rect 24994 38210 25314 38238
rect 25994 38542 26314 38550
rect 25994 38238 26002 38542
rect 26306 38238 26314 38542
rect 25994 38210 26314 38238
rect 26994 38542 27314 38550
rect 26994 38238 27002 38542
rect 27306 38238 27314 38542
rect 26994 38210 27314 38238
rect 27994 38542 28314 38550
rect 27994 38238 28002 38542
rect 28306 38238 28314 38542
rect 27994 38210 28314 38238
rect 28994 38542 29314 38550
rect 28994 38238 29002 38542
rect 29306 38238 29314 38542
rect 28994 38210 29314 38238
rect 29994 38542 30314 38550
rect 29994 38238 30002 38542
rect 30306 38238 30314 38542
rect 29994 38210 30314 38238
rect 30994 38542 31314 38550
rect 30994 38238 31002 38542
rect 31306 38238 31314 38542
rect 30994 38210 31314 38238
rect 31994 38542 32314 38550
rect 31994 38238 32002 38542
rect 32306 38238 32314 38542
rect 31994 38210 32314 38238
rect 32994 38542 33314 38550
rect 32994 38238 33002 38542
rect 33306 38238 33314 38542
rect 32994 38210 33314 38238
rect 33994 38542 34314 38550
rect 33994 38238 34002 38542
rect 34306 38238 34314 38542
rect 33994 38210 34314 38238
rect -74825 38202 -58825 38210
rect -74825 37898 -74817 38202
rect -74513 37898 -74477 38202
rect -74173 37898 -74137 38202
rect -73513 37898 -73477 38202
rect -73173 37898 -73137 38202
rect -72513 37898 -72477 38202
rect -72173 37898 -72137 38202
rect -71513 37898 -71477 38202
rect -71173 37898 -71137 38202
rect -70513 37898 -70477 38202
rect -70173 37898 -70137 38202
rect -69513 37898 -69477 38202
rect -69173 37898 -69137 38202
rect -68513 37898 -68477 38202
rect -68173 37898 -68137 38202
rect -67513 37898 -67477 38202
rect -67173 37898 -67137 38202
rect -66513 37898 -66477 38202
rect -66173 37898 -66137 38202
rect -65513 37898 -65477 38202
rect -65173 37898 -65137 38202
rect -64513 37898 -64477 38202
rect -64173 37898 -64137 38202
rect -63513 37898 -63477 38202
rect -63173 37898 -63137 38202
rect -62513 37898 -62477 38202
rect -62173 37898 -62137 38202
rect -61513 37898 -61477 38202
rect -61173 37898 -61137 38202
rect -60513 37898 -60477 38202
rect -60173 37898 -60137 38202
rect -59513 37898 -59477 38202
rect -59173 37898 -59137 38202
rect -58833 37898 -58825 38202
rect -74825 37890 -58825 37898
rect 9654 38202 34654 38210
rect 9654 37898 9662 38202
rect 9966 37898 10002 38202
rect 10306 37898 10342 38202
rect 10966 37898 11002 38202
rect 11306 37898 11342 38202
rect 11966 37898 12002 38202
rect 12306 37898 12342 38202
rect 12966 37898 13002 38202
rect 13306 37898 13342 38202
rect 13966 37898 14002 38202
rect 14306 37898 14342 38202
rect 14966 37898 15002 38202
rect 15306 37898 15342 38202
rect 15966 37898 16002 38202
rect 16306 37898 16342 38202
rect 16966 37898 17002 38202
rect 17306 37898 17342 38202
rect 17966 37898 18002 38202
rect 18306 37898 18342 38202
rect 18966 37898 19002 38202
rect 19306 37898 19342 38202
rect 19966 37898 20002 38202
rect 20306 37898 20342 38202
rect 20966 37898 21002 38202
rect 21306 37898 21342 38202
rect 21966 37898 22002 38202
rect 22306 37898 22342 38202
rect 22966 37898 23002 38202
rect 23306 37898 23342 38202
rect 23966 37898 24002 38202
rect 24306 37898 24342 38202
rect 24966 37898 25002 38202
rect 25306 37898 25342 38202
rect 25966 37898 26002 38202
rect 26306 37898 26342 38202
rect 26966 37898 27002 38202
rect 27306 37898 27342 38202
rect 27966 37898 28002 38202
rect 28306 37898 28342 38202
rect 28966 37898 29002 38202
rect 29306 37898 29342 38202
rect 29966 37898 30002 38202
rect 30306 37898 30342 38202
rect 30966 37898 31002 38202
rect 31306 37898 31342 38202
rect 31966 37898 32002 38202
rect 32306 37898 32342 38202
rect 32966 37898 33002 38202
rect 33306 37898 33342 38202
rect 33966 37898 34002 38202
rect 34306 37898 34342 38202
rect 34646 37898 34654 38202
rect 9654 37890 34654 37898
rect -74485 37862 -74165 37890
rect -74485 37238 -74477 37862
rect -74173 37238 -74165 37862
rect -74485 37210 -74165 37238
rect -73485 37862 -73165 37890
rect -73485 37238 -73477 37862
rect -73173 37238 -73165 37862
rect -73485 37210 -73165 37238
rect -72485 37862 -72165 37890
rect -72485 37238 -72477 37862
rect -72173 37238 -72165 37862
rect -72485 37210 -72165 37238
rect -71485 37862 -71165 37890
rect -71485 37238 -71477 37862
rect -71173 37238 -71165 37862
rect -71485 37210 -71165 37238
rect -70485 37862 -70165 37890
rect -70485 37238 -70477 37862
rect -70173 37238 -70165 37862
rect -70485 37210 -70165 37238
rect -69485 37862 -69165 37890
rect -69485 37238 -69477 37862
rect -69173 37238 -69165 37862
rect -69485 37210 -69165 37238
rect -68485 37862 -68165 37890
rect -68485 37238 -68477 37862
rect -68173 37238 -68165 37862
rect -68485 37210 -68165 37238
rect -67485 37862 -67165 37890
rect -67485 37238 -67477 37862
rect -67173 37238 -67165 37862
rect -67485 37210 -67165 37238
rect -66485 37862 -66165 37890
rect -66485 37238 -66477 37862
rect -66173 37238 -66165 37862
rect -66485 37210 -66165 37238
rect -65485 37862 -65165 37890
rect -65485 37238 -65477 37862
rect -65173 37238 -65165 37862
rect -65485 37210 -65165 37238
rect -64485 37862 -64165 37890
rect -64485 37238 -64477 37862
rect -64173 37238 -64165 37862
rect -64485 37210 -64165 37238
rect -63485 37862 -63165 37890
rect -63485 37238 -63477 37862
rect -63173 37238 -63165 37862
rect -63485 37210 -63165 37238
rect -62485 37862 -62165 37890
rect -62485 37238 -62477 37862
rect -62173 37238 -62165 37862
rect -62485 37210 -62165 37238
rect -61485 37862 -61165 37890
rect -61485 37238 -61477 37862
rect -61173 37238 -61165 37862
rect -61485 37210 -61165 37238
rect -60485 37862 -60165 37890
rect -60485 37238 -60477 37862
rect -60173 37238 -60165 37862
rect -60485 37210 -60165 37238
rect -59485 37862 -59165 37890
rect -59485 37238 -59477 37862
rect -59173 37238 -59165 37862
rect -59485 37210 -59165 37238
rect 9994 37862 10314 37890
rect 9994 37238 10002 37862
rect 10306 37238 10314 37862
rect 9994 37210 10314 37238
rect 10994 37862 11314 37890
rect 10994 37238 11002 37862
rect 11306 37238 11314 37862
rect 10994 37210 11314 37238
rect 11994 37862 12314 37890
rect 11994 37238 12002 37862
rect 12306 37238 12314 37862
rect 11994 37210 12314 37238
rect 12994 37862 13314 37890
rect 12994 37238 13002 37862
rect 13306 37238 13314 37862
rect 12994 37210 13314 37238
rect 13994 37862 14314 37890
rect 13994 37238 14002 37862
rect 14306 37238 14314 37862
rect 13994 37210 14314 37238
rect 14994 37862 15314 37890
rect 14994 37238 15002 37862
rect 15306 37238 15314 37862
rect 14994 37210 15314 37238
rect 15994 37862 16314 37890
rect 15994 37238 16002 37862
rect 16306 37238 16314 37862
rect 15994 37210 16314 37238
rect 16994 37862 17314 37890
rect 16994 37238 17002 37862
rect 17306 37238 17314 37862
rect 16994 37210 17314 37238
rect 17994 37862 18314 37890
rect 17994 37238 18002 37862
rect 18306 37238 18314 37862
rect 17994 37210 18314 37238
rect 18994 37862 19314 37890
rect 18994 37238 19002 37862
rect 19306 37238 19314 37862
rect 18994 37210 19314 37238
rect 19994 37862 20314 37890
rect 19994 37238 20002 37862
rect 20306 37238 20314 37862
rect 19994 37210 20314 37238
rect 20994 37862 21314 37890
rect 20994 37238 21002 37862
rect 21306 37238 21314 37862
rect 20994 37210 21314 37238
rect 21994 37862 22314 37890
rect 21994 37238 22002 37862
rect 22306 37238 22314 37862
rect 21994 37210 22314 37238
rect 22994 37862 23314 37890
rect 22994 37238 23002 37862
rect 23306 37238 23314 37862
rect 22994 37210 23314 37238
rect 23994 37862 24314 37890
rect 23994 37238 24002 37862
rect 24306 37238 24314 37862
rect 23994 37210 24314 37238
rect 24994 37862 25314 37890
rect 24994 37238 25002 37862
rect 25306 37238 25314 37862
rect 24994 37210 25314 37238
rect 25994 37862 26314 37890
rect 25994 37238 26002 37862
rect 26306 37238 26314 37862
rect 25994 37210 26314 37238
rect 26994 37862 27314 37890
rect 26994 37238 27002 37862
rect 27306 37238 27314 37862
rect 26994 37210 27314 37238
rect 27994 37862 28314 37890
rect 27994 37238 28002 37862
rect 28306 37238 28314 37862
rect 27994 37210 28314 37238
rect 28994 37862 29314 37890
rect 28994 37238 29002 37862
rect 29306 37238 29314 37862
rect 28994 37210 29314 37238
rect 29994 37862 30314 37890
rect 29994 37238 30002 37862
rect 30306 37238 30314 37862
rect 29994 37210 30314 37238
rect 30994 37862 31314 37890
rect 30994 37238 31002 37862
rect 31306 37238 31314 37862
rect 30994 37210 31314 37238
rect 31994 37862 32314 37890
rect 31994 37238 32002 37862
rect 32306 37238 32314 37862
rect 31994 37210 32314 37238
rect 32994 37862 33314 37890
rect 32994 37238 33002 37862
rect 33306 37238 33314 37862
rect 32994 37210 33314 37238
rect 33994 37862 34314 37890
rect 33994 37238 34002 37862
rect 34306 37238 34314 37862
rect 33994 37210 34314 37238
rect -74825 37202 -58825 37210
rect -74825 36898 -74817 37202
rect -74513 36898 -74477 37202
rect -74173 36898 -74137 37202
rect -73513 36898 -73477 37202
rect -73173 36898 -73137 37202
rect -72513 36898 -72477 37202
rect -72173 36898 -72137 37202
rect -71513 36898 -71477 37202
rect -71173 36898 -71137 37202
rect -70513 36898 -70477 37202
rect -70173 36898 -70137 37202
rect -69513 36898 -69477 37202
rect -69173 36898 -69137 37202
rect -68513 36898 -68477 37202
rect -68173 36898 -68137 37202
rect -67513 36898 -67477 37202
rect -67173 36898 -67137 37202
rect -66513 36898 -66477 37202
rect -66173 36898 -66137 37202
rect -65513 36898 -65477 37202
rect -65173 36898 -65137 37202
rect -64513 36898 -64477 37202
rect -64173 36898 -64137 37202
rect -63513 36898 -63477 37202
rect -63173 36898 -63137 37202
rect -62513 36898 -62477 37202
rect -62173 36898 -62137 37202
rect -61513 36898 -61477 37202
rect -61173 36898 -61137 37202
rect -60513 36898 -60477 37202
rect -60173 36898 -60137 37202
rect -59513 36898 -59477 37202
rect -59173 36898 -59137 37202
rect -58833 36898 -58825 37202
rect -74825 36890 -58825 36898
rect 9654 37202 34654 37210
rect 9654 36898 9662 37202
rect 9966 36898 10002 37202
rect 10306 36898 10342 37202
rect 10966 36898 11002 37202
rect 11306 36898 11342 37202
rect 11966 36898 12002 37202
rect 12306 36898 12342 37202
rect 12966 36898 13002 37202
rect 13306 36898 13342 37202
rect 13966 36898 14002 37202
rect 14306 36898 14342 37202
rect 14966 36898 15002 37202
rect 15306 36898 15342 37202
rect 15966 36898 16002 37202
rect 16306 36898 16342 37202
rect 16966 36898 17002 37202
rect 17306 36898 17342 37202
rect 17966 36898 18002 37202
rect 18306 36898 18342 37202
rect 18966 36898 19002 37202
rect 19306 36898 19342 37202
rect 19966 36898 20002 37202
rect 20306 36898 20342 37202
rect 20966 36898 21002 37202
rect 21306 36898 21342 37202
rect 21966 36898 22002 37202
rect 22306 36898 22342 37202
rect 22966 36898 23002 37202
rect 23306 36898 23342 37202
rect 23966 36898 24002 37202
rect 24306 36898 24342 37202
rect 24966 36898 25002 37202
rect 25306 36898 25342 37202
rect 25966 36898 26002 37202
rect 26306 36898 26342 37202
rect 26966 36898 27002 37202
rect 27306 36898 27342 37202
rect 27966 36898 28002 37202
rect 28306 36898 28342 37202
rect 28966 36898 29002 37202
rect 29306 36898 29342 37202
rect 29966 36898 30002 37202
rect 30306 36898 30342 37202
rect 30966 36898 31002 37202
rect 31306 36898 31342 37202
rect 31966 36898 32002 37202
rect 32306 36898 32342 37202
rect 32966 36898 33002 37202
rect 33306 36898 33342 37202
rect 33966 36898 34002 37202
rect 34306 36898 34342 37202
rect 34646 36898 34654 37202
rect 9654 36890 34654 36898
rect -74485 36862 -74165 36890
rect -74485 36238 -74477 36862
rect -74173 36238 -74165 36862
rect -74485 36210 -74165 36238
rect -73485 36862 -73165 36890
rect -73485 36238 -73477 36862
rect -73173 36238 -73165 36862
rect -73485 36210 -73165 36238
rect -72485 36862 -72165 36890
rect -72485 36238 -72477 36862
rect -72173 36238 -72165 36862
rect -72485 36210 -72165 36238
rect -71485 36862 -71165 36890
rect -71485 36238 -71477 36862
rect -71173 36238 -71165 36862
rect -71485 36210 -71165 36238
rect -70485 36862 -70165 36890
rect -70485 36238 -70477 36862
rect -70173 36238 -70165 36862
rect -70485 36210 -70165 36238
rect -69485 36862 -69165 36890
rect -69485 36238 -69477 36862
rect -69173 36238 -69165 36862
rect -69485 36210 -69165 36238
rect -68485 36862 -68165 36890
rect -68485 36238 -68477 36862
rect -68173 36238 -68165 36862
rect -68485 36210 -68165 36238
rect -67485 36862 -67165 36890
rect -67485 36238 -67477 36862
rect -67173 36238 -67165 36862
rect -67485 36210 -67165 36238
rect -66485 36862 -66165 36890
rect -66485 36238 -66477 36862
rect -66173 36238 -66165 36862
rect -66485 36210 -66165 36238
rect -65485 36862 -65165 36890
rect -65485 36238 -65477 36862
rect -65173 36238 -65165 36862
rect -65485 36210 -65165 36238
rect -64485 36862 -64165 36890
rect -64485 36238 -64477 36862
rect -64173 36238 -64165 36862
rect -64485 36210 -64165 36238
rect -63485 36862 -63165 36890
rect -63485 36238 -63477 36862
rect -63173 36238 -63165 36862
rect -63485 36210 -63165 36238
rect -62485 36862 -62165 36890
rect -62485 36238 -62477 36862
rect -62173 36238 -62165 36862
rect -62485 36210 -62165 36238
rect -61485 36862 -61165 36890
rect -61485 36238 -61477 36862
rect -61173 36238 -61165 36862
rect -61485 36210 -61165 36238
rect -60485 36862 -60165 36890
rect -60485 36238 -60477 36862
rect -60173 36238 -60165 36862
rect -60485 36210 -60165 36238
rect -59485 36862 -59165 36890
rect -59485 36238 -59477 36862
rect -59173 36238 -59165 36862
rect -59485 36210 -59165 36238
rect 9994 36862 10314 36890
rect 9994 36238 10002 36862
rect 10306 36238 10314 36862
rect 9994 36210 10314 36238
rect 10994 36862 11314 36890
rect 10994 36238 11002 36862
rect 11306 36238 11314 36862
rect 10994 36210 11314 36238
rect 11994 36862 12314 36890
rect 11994 36238 12002 36862
rect 12306 36238 12314 36862
rect 11994 36210 12314 36238
rect 12994 36862 13314 36890
rect 12994 36238 13002 36862
rect 13306 36238 13314 36862
rect 12994 36210 13314 36238
rect 13994 36862 14314 36890
rect 13994 36238 14002 36862
rect 14306 36238 14314 36862
rect 13994 36210 14314 36238
rect 14994 36862 15314 36890
rect 14994 36238 15002 36862
rect 15306 36238 15314 36862
rect 14994 36210 15314 36238
rect 15994 36862 16314 36890
rect 15994 36238 16002 36862
rect 16306 36238 16314 36862
rect 15994 36210 16314 36238
rect 16994 36862 17314 36890
rect 16994 36238 17002 36862
rect 17306 36238 17314 36862
rect 16994 36210 17314 36238
rect 17994 36862 18314 36890
rect 17994 36238 18002 36862
rect 18306 36238 18314 36862
rect 17994 36210 18314 36238
rect 18994 36862 19314 36890
rect 18994 36238 19002 36862
rect 19306 36238 19314 36862
rect 18994 36210 19314 36238
rect 19994 36862 20314 36890
rect 19994 36238 20002 36862
rect 20306 36238 20314 36862
rect 19994 36210 20314 36238
rect 20994 36862 21314 36890
rect 20994 36238 21002 36862
rect 21306 36238 21314 36862
rect 20994 36210 21314 36238
rect 21994 36862 22314 36890
rect 21994 36238 22002 36862
rect 22306 36238 22314 36862
rect 21994 36210 22314 36238
rect 22994 36862 23314 36890
rect 22994 36238 23002 36862
rect 23306 36238 23314 36862
rect 22994 36210 23314 36238
rect 23994 36862 24314 36890
rect 23994 36238 24002 36862
rect 24306 36238 24314 36862
rect 23994 36210 24314 36238
rect 24994 36862 25314 36890
rect 24994 36238 25002 36862
rect 25306 36238 25314 36862
rect 24994 36210 25314 36238
rect 25994 36862 26314 36890
rect 25994 36238 26002 36862
rect 26306 36238 26314 36862
rect 25994 36210 26314 36238
rect 26994 36862 27314 36890
rect 26994 36238 27002 36862
rect 27306 36238 27314 36862
rect 26994 36210 27314 36238
rect 27994 36862 28314 36890
rect 27994 36238 28002 36862
rect 28306 36238 28314 36862
rect 27994 36210 28314 36238
rect 28994 36862 29314 36890
rect 28994 36238 29002 36862
rect 29306 36238 29314 36862
rect 28994 36210 29314 36238
rect 29994 36862 30314 36890
rect 29994 36238 30002 36862
rect 30306 36238 30314 36862
rect 29994 36210 30314 36238
rect 30994 36862 31314 36890
rect 30994 36238 31002 36862
rect 31306 36238 31314 36862
rect 30994 36210 31314 36238
rect 31994 36862 32314 36890
rect 31994 36238 32002 36862
rect 32306 36238 32314 36862
rect 31994 36210 32314 36238
rect 32994 36862 33314 36890
rect 32994 36238 33002 36862
rect 33306 36238 33314 36862
rect 32994 36210 33314 36238
rect 33994 36862 34314 36890
rect 33994 36238 34002 36862
rect 34306 36238 34314 36862
rect 33994 36210 34314 36238
rect -74825 36202 -58825 36210
rect -74825 35898 -74817 36202
rect -74513 35898 -74477 36202
rect -74173 35898 -74137 36202
rect -73513 35898 -73477 36202
rect -73173 35898 -73137 36202
rect -72513 35898 -72477 36202
rect -72173 35898 -72137 36202
rect -71513 35898 -71477 36202
rect -71173 35898 -71137 36202
rect -70513 35898 -70477 36202
rect -70173 35898 -70137 36202
rect -69513 35898 -69477 36202
rect -69173 35898 -69137 36202
rect -68513 35898 -68477 36202
rect -68173 35898 -68137 36202
rect -67513 35898 -67477 36202
rect -67173 35898 -67137 36202
rect -66513 35898 -66477 36202
rect -66173 35898 -66137 36202
rect -65513 35898 -65477 36202
rect -65173 35898 -65137 36202
rect -64513 35898 -64477 36202
rect -64173 35898 -64137 36202
rect -63513 35898 -63477 36202
rect -63173 35898 -63137 36202
rect -62513 35898 -62477 36202
rect -62173 35898 -62137 36202
rect -61513 35898 -61477 36202
rect -61173 35898 -61137 36202
rect -60513 35898 -60477 36202
rect -60173 35898 -60137 36202
rect -59513 35898 -59477 36202
rect -59173 35898 -59137 36202
rect -58833 35898 -58825 36202
rect -74825 35890 -58825 35898
rect 9654 36202 34654 36210
rect 9654 35898 9662 36202
rect 9966 35898 10002 36202
rect 10306 35898 10342 36202
rect 10966 35898 11002 36202
rect 11306 35898 11342 36202
rect 11966 35898 12002 36202
rect 12306 35898 12342 36202
rect 12966 35898 13002 36202
rect 13306 35898 13342 36202
rect 13966 35898 14002 36202
rect 14306 35898 14342 36202
rect 14966 35898 15002 36202
rect 15306 35898 15342 36202
rect 15966 35898 16002 36202
rect 16306 35898 16342 36202
rect 16966 35898 17002 36202
rect 17306 35898 17342 36202
rect 17966 35898 18002 36202
rect 18306 35898 18342 36202
rect 18966 35898 19002 36202
rect 19306 35898 19342 36202
rect 19966 35898 20002 36202
rect 20306 35898 20342 36202
rect 20966 35898 21002 36202
rect 21306 35898 21342 36202
rect 21966 35898 22002 36202
rect 22306 35898 22342 36202
rect 22966 35898 23002 36202
rect 23306 35898 23342 36202
rect 23966 35898 24002 36202
rect 24306 35898 24342 36202
rect 24966 35898 25002 36202
rect 25306 35898 25342 36202
rect 25966 35898 26002 36202
rect 26306 35898 26342 36202
rect 26966 35898 27002 36202
rect 27306 35898 27342 36202
rect 27966 35898 28002 36202
rect 28306 35898 28342 36202
rect 28966 35898 29002 36202
rect 29306 35898 29342 36202
rect 29966 35898 30002 36202
rect 30306 35898 30342 36202
rect 30966 35898 31002 36202
rect 31306 35898 31342 36202
rect 31966 35898 32002 36202
rect 32306 35898 32342 36202
rect 32966 35898 33002 36202
rect 33306 35898 33342 36202
rect 33966 35898 34002 36202
rect 34306 35898 34342 36202
rect 34646 35898 34654 36202
rect 9654 35890 34654 35898
rect -74485 35862 -74165 35890
rect -74485 35238 -74477 35862
rect -74173 35238 -74165 35862
rect -74485 35210 -74165 35238
rect -73485 35862 -73165 35890
rect -73485 35238 -73477 35862
rect -73173 35238 -73165 35862
rect -73485 35210 -73165 35238
rect -72485 35862 -72165 35890
rect -72485 35238 -72477 35862
rect -72173 35238 -72165 35862
rect -72485 35210 -72165 35238
rect -71485 35862 -71165 35890
rect -71485 35238 -71477 35862
rect -71173 35238 -71165 35862
rect -71485 35210 -71165 35238
rect -70485 35862 -70165 35890
rect -70485 35238 -70477 35862
rect -70173 35238 -70165 35862
rect -70485 35210 -70165 35238
rect -69485 35862 -69165 35890
rect -69485 35238 -69477 35862
rect -69173 35238 -69165 35862
rect -69485 35210 -69165 35238
rect -68485 35862 -68165 35890
rect -68485 35238 -68477 35862
rect -68173 35238 -68165 35862
rect -68485 35210 -68165 35238
rect -67485 35862 -67165 35890
rect -67485 35238 -67477 35862
rect -67173 35238 -67165 35862
rect -67485 35210 -67165 35238
rect -66485 35862 -66165 35890
rect -66485 35238 -66477 35862
rect -66173 35238 -66165 35862
rect -66485 35210 -66165 35238
rect -65485 35862 -65165 35890
rect -65485 35238 -65477 35862
rect -65173 35238 -65165 35862
rect -65485 35210 -65165 35238
rect -64485 35862 -64165 35890
rect -64485 35238 -64477 35862
rect -64173 35238 -64165 35862
rect -64485 35210 -64165 35238
rect -63485 35862 -63165 35890
rect -63485 35238 -63477 35862
rect -63173 35238 -63165 35862
rect -63485 35210 -63165 35238
rect -62485 35862 -62165 35890
rect -62485 35238 -62477 35862
rect -62173 35238 -62165 35862
rect -62485 35210 -62165 35238
rect -61485 35862 -61165 35890
rect -61485 35238 -61477 35862
rect -61173 35238 -61165 35862
rect -61485 35210 -61165 35238
rect -60485 35862 -60165 35890
rect -60485 35238 -60477 35862
rect -60173 35238 -60165 35862
rect -60485 35210 -60165 35238
rect -59485 35862 -59165 35890
rect -59485 35238 -59477 35862
rect -59173 35238 -59165 35862
rect -59485 35210 -59165 35238
rect 9994 35862 10314 35890
rect 9994 35238 10002 35862
rect 10306 35238 10314 35862
rect 9994 35210 10314 35238
rect 10994 35862 11314 35890
rect 10994 35238 11002 35862
rect 11306 35238 11314 35862
rect 10994 35210 11314 35238
rect 11994 35862 12314 35890
rect 11994 35238 12002 35862
rect 12306 35238 12314 35862
rect 11994 35210 12314 35238
rect 12994 35862 13314 35890
rect 12994 35238 13002 35862
rect 13306 35238 13314 35862
rect 12994 35210 13314 35238
rect 13994 35862 14314 35890
rect 13994 35238 14002 35862
rect 14306 35238 14314 35862
rect 13994 35210 14314 35238
rect 14994 35862 15314 35890
rect 14994 35238 15002 35862
rect 15306 35238 15314 35862
rect 14994 35210 15314 35238
rect 15994 35862 16314 35890
rect 15994 35238 16002 35862
rect 16306 35238 16314 35862
rect 15994 35210 16314 35238
rect 16994 35862 17314 35890
rect 16994 35238 17002 35862
rect 17306 35238 17314 35862
rect 16994 35210 17314 35238
rect 17994 35862 18314 35890
rect 17994 35238 18002 35862
rect 18306 35238 18314 35862
rect 17994 35210 18314 35238
rect 18994 35862 19314 35890
rect 18994 35238 19002 35862
rect 19306 35238 19314 35862
rect 18994 35210 19314 35238
rect 19994 35862 20314 35890
rect 19994 35238 20002 35862
rect 20306 35238 20314 35862
rect 19994 35210 20314 35238
rect 20994 35862 21314 35890
rect 20994 35238 21002 35862
rect 21306 35238 21314 35862
rect 20994 35210 21314 35238
rect 21994 35862 22314 35890
rect 21994 35238 22002 35862
rect 22306 35238 22314 35862
rect 21994 35210 22314 35238
rect 22994 35862 23314 35890
rect 22994 35238 23002 35862
rect 23306 35238 23314 35862
rect 22994 35210 23314 35238
rect 23994 35862 24314 35890
rect 23994 35238 24002 35862
rect 24306 35238 24314 35862
rect 23994 35210 24314 35238
rect 24994 35862 25314 35890
rect 24994 35238 25002 35862
rect 25306 35238 25314 35862
rect 24994 35210 25314 35238
rect 25994 35862 26314 35890
rect 25994 35238 26002 35862
rect 26306 35238 26314 35862
rect 25994 35210 26314 35238
rect 26994 35862 27314 35890
rect 26994 35238 27002 35862
rect 27306 35238 27314 35862
rect 26994 35210 27314 35238
rect 27994 35862 28314 35890
rect 27994 35238 28002 35862
rect 28306 35238 28314 35862
rect 27994 35210 28314 35238
rect 28994 35862 29314 35890
rect 28994 35238 29002 35862
rect 29306 35238 29314 35862
rect 28994 35210 29314 35238
rect 29994 35862 30314 35890
rect 29994 35238 30002 35862
rect 30306 35238 30314 35862
rect 29994 35210 30314 35238
rect 30994 35862 31314 35890
rect 30994 35238 31002 35862
rect 31306 35238 31314 35862
rect 30994 35210 31314 35238
rect 31994 35862 32314 35890
rect 31994 35238 32002 35862
rect 32306 35238 32314 35862
rect 31994 35210 32314 35238
rect 32994 35862 33314 35890
rect 32994 35238 33002 35862
rect 33306 35238 33314 35862
rect 32994 35210 33314 35238
rect 33994 35862 34314 35890
rect 33994 35238 34002 35862
rect 34306 35238 34314 35862
rect 33994 35210 34314 35238
rect -74825 35202 -58825 35210
rect -74825 34898 -74817 35202
rect -74513 34898 -74477 35202
rect -74173 34898 -74137 35202
rect -73513 34898 -73477 35202
rect -73173 34898 -73137 35202
rect -72513 34898 -72477 35202
rect -72173 34898 -72137 35202
rect -71513 34898 -71477 35202
rect -71173 34898 -71137 35202
rect -70513 34898 -70477 35202
rect -70173 34898 -70137 35202
rect -69513 34898 -69477 35202
rect -69173 34898 -69137 35202
rect -68513 34898 -68477 35202
rect -68173 34898 -68137 35202
rect -67513 34898 -67477 35202
rect -67173 34898 -67137 35202
rect -66513 34898 -66477 35202
rect -66173 34898 -66137 35202
rect -65513 34898 -65477 35202
rect -65173 34898 -65137 35202
rect -64513 34898 -64477 35202
rect -64173 34898 -64137 35202
rect -63513 34898 -63477 35202
rect -63173 34898 -63137 35202
rect -62513 34898 -62477 35202
rect -62173 34898 -62137 35202
rect -61513 34898 -61477 35202
rect -61173 34898 -61137 35202
rect -60513 34898 -60477 35202
rect -60173 34898 -60137 35202
rect -59513 34898 -59477 35202
rect -59173 34898 -59137 35202
rect -58833 34898 -58825 35202
rect -74825 34890 -58825 34898
rect 9654 35202 34654 35210
rect 9654 34898 9662 35202
rect 9966 34898 10002 35202
rect 10306 34898 10342 35202
rect 10966 34898 11002 35202
rect 11306 34898 11342 35202
rect 11966 34898 12002 35202
rect 12306 34898 12342 35202
rect 12966 34898 13002 35202
rect 13306 34898 13342 35202
rect 13966 34898 14002 35202
rect 14306 34898 14342 35202
rect 14966 34898 15002 35202
rect 15306 34898 15342 35202
rect 15966 34898 16002 35202
rect 16306 34898 16342 35202
rect 16966 34898 17002 35202
rect 17306 34898 17342 35202
rect 17966 34898 18002 35202
rect 18306 34898 18342 35202
rect 18966 34898 19002 35202
rect 19306 34898 19342 35202
rect 19966 34898 20002 35202
rect 20306 34898 20342 35202
rect 20966 34898 21002 35202
rect 21306 34898 21342 35202
rect 21966 34898 22002 35202
rect 22306 34898 22342 35202
rect 22966 34898 23002 35202
rect 23306 34898 23342 35202
rect 23966 34898 24002 35202
rect 24306 34898 24342 35202
rect 24966 34898 25002 35202
rect 25306 34898 25342 35202
rect 25966 34898 26002 35202
rect 26306 34898 26342 35202
rect 26966 34898 27002 35202
rect 27306 34898 27342 35202
rect 27966 34898 28002 35202
rect 28306 34898 28342 35202
rect 28966 34898 29002 35202
rect 29306 34898 29342 35202
rect 29966 34898 30002 35202
rect 30306 34898 30342 35202
rect 30966 34898 31002 35202
rect 31306 34898 31342 35202
rect 31966 34898 32002 35202
rect 32306 34898 32342 35202
rect 32966 34898 33002 35202
rect 33306 34898 33342 35202
rect 33966 34898 34002 35202
rect 34306 34898 34342 35202
rect 34646 34898 34654 35202
rect 9654 34890 34654 34898
rect -74485 34862 -74165 34890
rect -74485 34238 -74477 34862
rect -74173 34238 -74165 34862
rect -74485 34210 -74165 34238
rect -73485 34862 -73165 34890
rect -73485 34238 -73477 34862
rect -73173 34238 -73165 34862
rect -73485 34210 -73165 34238
rect -72485 34862 -72165 34890
rect -72485 34238 -72477 34862
rect -72173 34238 -72165 34862
rect -72485 34210 -72165 34238
rect -71485 34862 -71165 34890
rect -71485 34238 -71477 34862
rect -71173 34238 -71165 34862
rect -71485 34210 -71165 34238
rect -70485 34862 -70165 34890
rect -70485 34238 -70477 34862
rect -70173 34238 -70165 34862
rect -70485 34210 -70165 34238
rect -69485 34862 -69165 34890
rect -69485 34238 -69477 34862
rect -69173 34238 -69165 34862
rect -69485 34210 -69165 34238
rect -68485 34862 -68165 34890
rect -68485 34238 -68477 34862
rect -68173 34238 -68165 34862
rect -68485 34210 -68165 34238
rect -67485 34862 -67165 34890
rect -67485 34238 -67477 34862
rect -67173 34238 -67165 34862
rect -67485 34210 -67165 34238
rect -66485 34862 -66165 34890
rect -66485 34238 -66477 34862
rect -66173 34238 -66165 34862
rect -66485 34210 -66165 34238
rect -65485 34862 -65165 34890
rect -65485 34238 -65477 34862
rect -65173 34238 -65165 34862
rect -65485 34210 -65165 34238
rect -64485 34862 -64165 34890
rect -64485 34238 -64477 34862
rect -64173 34238 -64165 34862
rect -64485 34210 -64165 34238
rect -63485 34862 -63165 34890
rect -63485 34238 -63477 34862
rect -63173 34238 -63165 34862
rect -63485 34210 -63165 34238
rect -62485 34862 -62165 34890
rect -62485 34238 -62477 34862
rect -62173 34238 -62165 34862
rect -62485 34210 -62165 34238
rect -61485 34862 -61165 34890
rect -61485 34238 -61477 34862
rect -61173 34238 -61165 34862
rect -61485 34210 -61165 34238
rect -60485 34862 -60165 34890
rect -60485 34238 -60477 34862
rect -60173 34238 -60165 34862
rect -60485 34210 -60165 34238
rect -59485 34862 -59165 34890
rect -59485 34238 -59477 34862
rect -59173 34238 -59165 34862
rect -59485 34210 -59165 34238
rect 9994 34862 10314 34890
rect 9994 34238 10002 34862
rect 10306 34238 10314 34862
rect 9994 34210 10314 34238
rect 10994 34862 11314 34890
rect 10994 34238 11002 34862
rect 11306 34238 11314 34862
rect 10994 34210 11314 34238
rect 11994 34862 12314 34890
rect 11994 34238 12002 34862
rect 12306 34238 12314 34862
rect 11994 34210 12314 34238
rect 12994 34862 13314 34890
rect 12994 34238 13002 34862
rect 13306 34238 13314 34862
rect 12994 34210 13314 34238
rect 13994 34862 14314 34890
rect 13994 34238 14002 34862
rect 14306 34238 14314 34862
rect 13994 34210 14314 34238
rect 14994 34862 15314 34890
rect 14994 34238 15002 34862
rect 15306 34238 15314 34862
rect 14994 34210 15314 34238
rect 15994 34862 16314 34890
rect 15994 34238 16002 34862
rect 16306 34238 16314 34862
rect 15994 34210 16314 34238
rect 16994 34862 17314 34890
rect 16994 34238 17002 34862
rect 17306 34238 17314 34862
rect 16994 34210 17314 34238
rect 17994 34862 18314 34890
rect 17994 34238 18002 34862
rect 18306 34238 18314 34862
rect 17994 34210 18314 34238
rect 18994 34862 19314 34890
rect 18994 34238 19002 34862
rect 19306 34238 19314 34862
rect 18994 34210 19314 34238
rect 19994 34862 20314 34890
rect 19994 34238 20002 34862
rect 20306 34238 20314 34862
rect 19994 34210 20314 34238
rect 20994 34862 21314 34890
rect 20994 34238 21002 34862
rect 21306 34238 21314 34862
rect 20994 34210 21314 34238
rect 21994 34862 22314 34890
rect 21994 34238 22002 34862
rect 22306 34238 22314 34862
rect 21994 34210 22314 34238
rect 22994 34862 23314 34890
rect 22994 34238 23002 34862
rect 23306 34238 23314 34862
rect 22994 34210 23314 34238
rect 23994 34862 24314 34890
rect 23994 34238 24002 34862
rect 24306 34238 24314 34862
rect 23994 34210 24314 34238
rect 24994 34862 25314 34890
rect 24994 34238 25002 34862
rect 25306 34238 25314 34862
rect 24994 34210 25314 34238
rect 25994 34862 26314 34890
rect 25994 34238 26002 34862
rect 26306 34238 26314 34862
rect 25994 34210 26314 34238
rect 26994 34862 27314 34890
rect 26994 34238 27002 34862
rect 27306 34238 27314 34862
rect 26994 34210 27314 34238
rect 27994 34862 28314 34890
rect 27994 34238 28002 34862
rect 28306 34238 28314 34862
rect 27994 34210 28314 34238
rect 28994 34862 29314 34890
rect 28994 34238 29002 34862
rect 29306 34238 29314 34862
rect 28994 34210 29314 34238
rect 29994 34862 30314 34890
rect 29994 34238 30002 34862
rect 30306 34238 30314 34862
rect 29994 34210 30314 34238
rect 30994 34862 31314 34890
rect 30994 34238 31002 34862
rect 31306 34238 31314 34862
rect 30994 34210 31314 34238
rect 31994 34862 32314 34890
rect 31994 34238 32002 34862
rect 32306 34238 32314 34862
rect 31994 34210 32314 34238
rect 32994 34862 33314 34890
rect 32994 34238 33002 34862
rect 33306 34238 33314 34862
rect 32994 34210 33314 34238
rect 33994 34862 34314 34890
rect 33994 34238 34002 34862
rect 34306 34238 34314 34862
rect 33994 34210 34314 34238
rect -74825 34202 -58825 34210
rect -74825 33898 -74817 34202
rect -74513 33898 -74477 34202
rect -74173 33898 -74137 34202
rect -73513 33898 -73477 34202
rect -73173 33898 -73137 34202
rect -72513 33898 -72477 34202
rect -72173 33898 -72137 34202
rect -71513 33898 -71477 34202
rect -71173 33898 -71137 34202
rect -70513 33898 -70477 34202
rect -70173 33898 -70137 34202
rect -69513 33898 -69477 34202
rect -69173 33898 -69137 34202
rect -68513 33898 -68477 34202
rect -68173 33898 -68137 34202
rect -67513 33898 -67477 34202
rect -67173 33898 -67137 34202
rect -66513 33898 -66477 34202
rect -66173 33898 -66137 34202
rect -65513 33898 -65477 34202
rect -65173 33898 -65137 34202
rect -64513 33898 -64477 34202
rect -64173 33898 -64137 34202
rect -63513 33898 -63477 34202
rect -63173 33898 -63137 34202
rect -62513 33898 -62477 34202
rect -62173 33898 -62137 34202
rect -61513 33898 -61477 34202
rect -61173 33898 -61137 34202
rect -60513 33898 -60477 34202
rect -60173 33898 -60137 34202
rect -59513 33898 -59477 34202
rect -59173 33898 -59137 34202
rect -58833 33898 -58825 34202
rect -74825 33890 -58825 33898
rect 9654 34202 34654 34210
rect 9654 33898 9662 34202
rect 9966 33898 10002 34202
rect 10306 33898 10342 34202
rect 10966 33898 11002 34202
rect 11306 33898 11342 34202
rect 11966 33898 12002 34202
rect 12306 33898 12342 34202
rect 12966 33898 13002 34202
rect 13306 33898 13342 34202
rect 13966 33898 14002 34202
rect 14306 33898 14342 34202
rect 14966 33898 15002 34202
rect 15306 33898 15342 34202
rect 15966 33898 16002 34202
rect 16306 33898 16342 34202
rect 16966 33898 17002 34202
rect 17306 33898 17342 34202
rect 17966 33898 18002 34202
rect 18306 33898 18342 34202
rect 18966 33898 19002 34202
rect 19306 33898 19342 34202
rect 19966 33898 20002 34202
rect 20306 33898 20342 34202
rect 20966 33898 21002 34202
rect 21306 33898 21342 34202
rect 21966 33898 22002 34202
rect 22306 33898 22342 34202
rect 22966 33898 23002 34202
rect 23306 33898 23342 34202
rect 23966 33898 24002 34202
rect 24306 33898 24342 34202
rect 24966 33898 25002 34202
rect 25306 33898 25342 34202
rect 25966 33898 26002 34202
rect 26306 33898 26342 34202
rect 26966 33898 27002 34202
rect 27306 33898 27342 34202
rect 27966 33898 28002 34202
rect 28306 33898 28342 34202
rect 28966 33898 29002 34202
rect 29306 33898 29342 34202
rect 29966 33898 30002 34202
rect 30306 33898 30342 34202
rect 30966 33898 31002 34202
rect 31306 33898 31342 34202
rect 31966 33898 32002 34202
rect 32306 33898 32342 34202
rect 32966 33898 33002 34202
rect 33306 33898 33342 34202
rect 33966 33898 34002 34202
rect 34306 33898 34342 34202
rect 34646 33898 34654 34202
rect 9654 33890 34654 33898
rect -74485 33862 -74165 33890
rect -74485 33238 -74477 33862
rect -74173 33238 -74165 33862
rect -74485 33210 -74165 33238
rect -73485 33862 -73165 33890
rect -73485 33238 -73477 33862
rect -73173 33238 -73165 33862
rect -73485 33210 -73165 33238
rect -72485 33862 -72165 33890
rect -72485 33238 -72477 33862
rect -72173 33238 -72165 33862
rect -72485 33210 -72165 33238
rect -71485 33862 -71165 33890
rect -71485 33238 -71477 33862
rect -71173 33238 -71165 33862
rect -71485 33210 -71165 33238
rect -70485 33862 -70165 33890
rect -70485 33238 -70477 33862
rect -70173 33238 -70165 33862
rect -70485 33210 -70165 33238
rect -69485 33862 -69165 33890
rect -69485 33238 -69477 33862
rect -69173 33238 -69165 33862
rect -69485 33210 -69165 33238
rect -68485 33862 -68165 33890
rect -68485 33238 -68477 33862
rect -68173 33238 -68165 33862
rect -68485 33210 -68165 33238
rect -67485 33862 -67165 33890
rect -67485 33238 -67477 33862
rect -67173 33238 -67165 33862
rect -67485 33210 -67165 33238
rect -66485 33862 -66165 33890
rect -66485 33238 -66477 33862
rect -66173 33238 -66165 33862
rect -66485 33210 -66165 33238
rect -65485 33862 -65165 33890
rect -65485 33238 -65477 33862
rect -65173 33238 -65165 33862
rect -65485 33210 -65165 33238
rect -64485 33862 -64165 33890
rect -64485 33238 -64477 33862
rect -64173 33238 -64165 33862
rect -64485 33210 -64165 33238
rect -63485 33862 -63165 33890
rect -63485 33238 -63477 33862
rect -63173 33238 -63165 33862
rect -63485 33210 -63165 33238
rect -62485 33862 -62165 33890
rect -62485 33238 -62477 33862
rect -62173 33238 -62165 33862
rect -62485 33210 -62165 33238
rect -61485 33862 -61165 33890
rect -61485 33238 -61477 33862
rect -61173 33238 -61165 33862
rect -61485 33210 -61165 33238
rect -60485 33862 -60165 33890
rect -60485 33238 -60477 33862
rect -60173 33238 -60165 33862
rect -60485 33210 -60165 33238
rect -59485 33862 -59165 33890
rect -59485 33238 -59477 33862
rect -59173 33238 -59165 33862
rect -59485 33210 -59165 33238
rect 9994 33862 10314 33890
rect 9994 33238 10002 33862
rect 10306 33238 10314 33862
rect 9994 33210 10314 33238
rect 10994 33862 11314 33890
rect 10994 33238 11002 33862
rect 11306 33238 11314 33862
rect 10994 33210 11314 33238
rect 11994 33862 12314 33890
rect 11994 33238 12002 33862
rect 12306 33238 12314 33862
rect 11994 33210 12314 33238
rect 12994 33862 13314 33890
rect 12994 33238 13002 33862
rect 13306 33238 13314 33862
rect 12994 33210 13314 33238
rect 13994 33862 14314 33890
rect 13994 33238 14002 33862
rect 14306 33238 14314 33862
rect 13994 33210 14314 33238
rect 14994 33862 15314 33890
rect 14994 33238 15002 33862
rect 15306 33238 15314 33862
rect 14994 33210 15314 33238
rect 15994 33862 16314 33890
rect 15994 33238 16002 33862
rect 16306 33238 16314 33862
rect 15994 33210 16314 33238
rect 16994 33862 17314 33890
rect 16994 33238 17002 33862
rect 17306 33238 17314 33862
rect 16994 33210 17314 33238
rect 17994 33862 18314 33890
rect 17994 33238 18002 33862
rect 18306 33238 18314 33862
rect 17994 33210 18314 33238
rect 18994 33862 19314 33890
rect 18994 33238 19002 33862
rect 19306 33238 19314 33862
rect 18994 33210 19314 33238
rect 19994 33862 20314 33890
rect 19994 33238 20002 33862
rect 20306 33238 20314 33862
rect 19994 33210 20314 33238
rect 20994 33862 21314 33890
rect 20994 33238 21002 33862
rect 21306 33238 21314 33862
rect 20994 33210 21314 33238
rect 21994 33862 22314 33890
rect 21994 33238 22002 33862
rect 22306 33238 22314 33862
rect 21994 33210 22314 33238
rect 22994 33862 23314 33890
rect 22994 33238 23002 33862
rect 23306 33238 23314 33862
rect 22994 33210 23314 33238
rect 23994 33862 24314 33890
rect 23994 33238 24002 33862
rect 24306 33238 24314 33862
rect 23994 33210 24314 33238
rect 24994 33862 25314 33890
rect 24994 33238 25002 33862
rect 25306 33238 25314 33862
rect 24994 33210 25314 33238
rect 25994 33862 26314 33890
rect 25994 33238 26002 33862
rect 26306 33238 26314 33862
rect 25994 33210 26314 33238
rect 26994 33862 27314 33890
rect 26994 33238 27002 33862
rect 27306 33238 27314 33862
rect 26994 33210 27314 33238
rect 27994 33862 28314 33890
rect 27994 33238 28002 33862
rect 28306 33238 28314 33862
rect 27994 33210 28314 33238
rect 28994 33862 29314 33890
rect 28994 33238 29002 33862
rect 29306 33238 29314 33862
rect 28994 33210 29314 33238
rect 29994 33862 30314 33890
rect 29994 33238 30002 33862
rect 30306 33238 30314 33862
rect 29994 33210 30314 33238
rect 30994 33862 31314 33890
rect 30994 33238 31002 33862
rect 31306 33238 31314 33862
rect 30994 33210 31314 33238
rect 31994 33862 32314 33890
rect 31994 33238 32002 33862
rect 32306 33238 32314 33862
rect 31994 33210 32314 33238
rect 32994 33862 33314 33890
rect 32994 33238 33002 33862
rect 33306 33238 33314 33862
rect 32994 33210 33314 33238
rect 33994 33862 34314 33890
rect 33994 33238 34002 33862
rect 34306 33238 34314 33862
rect 33994 33210 34314 33238
rect -74825 33202 -58825 33210
rect -74825 32898 -74817 33202
rect -74513 32898 -74477 33202
rect -74173 32898 -74137 33202
rect -73513 32898 -73477 33202
rect -73173 32898 -73137 33202
rect -72513 32898 -72477 33202
rect -72173 32898 -72137 33202
rect -71513 32898 -71477 33202
rect -71173 32898 -71137 33202
rect -70513 32898 -70477 33202
rect -70173 32898 -70137 33202
rect -69513 32898 -69477 33202
rect -69173 32898 -69137 33202
rect -68513 32898 -68477 33202
rect -68173 32898 -68137 33202
rect -67513 32898 -67477 33202
rect -67173 32898 -67137 33202
rect -66513 32898 -66477 33202
rect -66173 32898 -66137 33202
rect -65513 32898 -65477 33202
rect -65173 32898 -65137 33202
rect -64513 32898 -64477 33202
rect -64173 32898 -64137 33202
rect -63513 32898 -63477 33202
rect -63173 32898 -63137 33202
rect -62513 32898 -62477 33202
rect -62173 32898 -62137 33202
rect -61513 32898 -61477 33202
rect -61173 32898 -61137 33202
rect -60513 32898 -60477 33202
rect -60173 32898 -60137 33202
rect -59513 32898 -59477 33202
rect -59173 32898 -59137 33202
rect -58833 32898 -58825 33202
rect -74825 32890 -58825 32898
rect 9654 33202 34654 33210
rect 9654 32898 9662 33202
rect 9966 32898 10002 33202
rect 10306 32898 10342 33202
rect 10966 32898 11002 33202
rect 11306 32898 11342 33202
rect 11966 32898 12002 33202
rect 12306 32898 12342 33202
rect 12966 32898 13002 33202
rect 13306 32898 13342 33202
rect 13966 32898 14002 33202
rect 14306 32898 14342 33202
rect 14966 32898 15002 33202
rect 15306 32898 15342 33202
rect 15966 32898 16002 33202
rect 16306 32898 16342 33202
rect 16966 32898 17002 33202
rect 17306 32898 17342 33202
rect 17966 32898 18002 33202
rect 18306 32898 18342 33202
rect 18966 32898 19002 33202
rect 19306 32898 19342 33202
rect 19966 32898 20002 33202
rect 20306 32898 20342 33202
rect 20966 32898 21002 33202
rect 21306 32898 21342 33202
rect 21966 32898 22002 33202
rect 22306 32898 22342 33202
rect 22966 32898 23002 33202
rect 23306 32898 23342 33202
rect 23966 32898 24002 33202
rect 24306 32898 24342 33202
rect 24966 32898 25002 33202
rect 25306 32898 25342 33202
rect 25966 32898 26002 33202
rect 26306 32898 26342 33202
rect 26966 32898 27002 33202
rect 27306 32898 27342 33202
rect 27966 32898 28002 33202
rect 28306 32898 28342 33202
rect 28966 32898 29002 33202
rect 29306 32898 29342 33202
rect 29966 32898 30002 33202
rect 30306 32898 30342 33202
rect 30966 32898 31002 33202
rect 31306 32898 31342 33202
rect 31966 32898 32002 33202
rect 32306 32898 32342 33202
rect 32966 32898 33002 33202
rect 33306 32898 33342 33202
rect 33966 32898 34002 33202
rect 34306 32898 34342 33202
rect 34646 32898 34654 33202
rect 9654 32890 34654 32898
rect -74485 32862 -74165 32890
rect -74485 32238 -74477 32862
rect -74173 32238 -74165 32862
rect -74485 32210 -74165 32238
rect -73485 32862 -73165 32890
rect -73485 32238 -73477 32862
rect -73173 32238 -73165 32862
rect -73485 32210 -73165 32238
rect -72485 32862 -72165 32890
rect -72485 32238 -72477 32862
rect -72173 32238 -72165 32862
rect -72485 32210 -72165 32238
rect -71485 32862 -71165 32890
rect -71485 32238 -71477 32862
rect -71173 32238 -71165 32862
rect -71485 32210 -71165 32238
rect -70485 32862 -70165 32890
rect -70485 32238 -70477 32862
rect -70173 32238 -70165 32862
rect -70485 32210 -70165 32238
rect -69485 32862 -69165 32890
rect -69485 32238 -69477 32862
rect -69173 32238 -69165 32862
rect -69485 32210 -69165 32238
rect -68485 32862 -68165 32890
rect -68485 32238 -68477 32862
rect -68173 32238 -68165 32862
rect -68485 32210 -68165 32238
rect -67485 32862 -67165 32890
rect -67485 32238 -67477 32862
rect -67173 32238 -67165 32862
rect -67485 32210 -67165 32238
rect -66485 32862 -66165 32890
rect -66485 32238 -66477 32862
rect -66173 32238 -66165 32862
rect -66485 32210 -66165 32238
rect -65485 32862 -65165 32890
rect -65485 32238 -65477 32862
rect -65173 32238 -65165 32862
rect -65485 32210 -65165 32238
rect -64485 32862 -64165 32890
rect -64485 32238 -64477 32862
rect -64173 32238 -64165 32862
rect -64485 32210 -64165 32238
rect -63485 32862 -63165 32890
rect -63485 32238 -63477 32862
rect -63173 32238 -63165 32862
rect -63485 32210 -63165 32238
rect -62485 32862 -62165 32890
rect -62485 32238 -62477 32862
rect -62173 32238 -62165 32862
rect -62485 32210 -62165 32238
rect -61485 32862 -61165 32890
rect -61485 32238 -61477 32862
rect -61173 32238 -61165 32862
rect -61485 32210 -61165 32238
rect -60485 32862 -60165 32890
rect -60485 32238 -60477 32862
rect -60173 32238 -60165 32862
rect -60485 32210 -60165 32238
rect -59485 32862 -59165 32890
rect -59485 32238 -59477 32862
rect -59173 32238 -59165 32862
rect -59485 32210 -59165 32238
rect 9994 32862 10314 32890
rect 9994 32238 10002 32862
rect 10306 32238 10314 32862
rect 9994 32210 10314 32238
rect 10994 32862 11314 32890
rect 10994 32238 11002 32862
rect 11306 32238 11314 32862
rect 10994 32210 11314 32238
rect 11994 32862 12314 32890
rect 11994 32238 12002 32862
rect 12306 32238 12314 32862
rect 11994 32210 12314 32238
rect 12994 32862 13314 32890
rect 12994 32238 13002 32862
rect 13306 32238 13314 32862
rect 12994 32210 13314 32238
rect 13994 32862 14314 32890
rect 13994 32238 14002 32862
rect 14306 32238 14314 32862
rect 13994 32210 14314 32238
rect 14994 32862 15314 32890
rect 14994 32238 15002 32862
rect 15306 32238 15314 32862
rect 14994 32210 15314 32238
rect 15994 32862 16314 32890
rect 15994 32238 16002 32862
rect 16306 32238 16314 32862
rect 15994 32210 16314 32238
rect 16994 32862 17314 32890
rect 16994 32238 17002 32862
rect 17306 32238 17314 32862
rect 16994 32210 17314 32238
rect 17994 32862 18314 32890
rect 17994 32238 18002 32862
rect 18306 32238 18314 32862
rect 17994 32210 18314 32238
rect 18994 32862 19314 32890
rect 18994 32238 19002 32862
rect 19306 32238 19314 32862
rect 18994 32210 19314 32238
rect 19994 32862 20314 32890
rect 19994 32238 20002 32862
rect 20306 32238 20314 32862
rect 19994 32210 20314 32238
rect 20994 32862 21314 32890
rect 20994 32238 21002 32862
rect 21306 32238 21314 32862
rect 20994 32210 21314 32238
rect 21994 32862 22314 32890
rect 21994 32238 22002 32862
rect 22306 32238 22314 32862
rect 21994 32210 22314 32238
rect 22994 32862 23314 32890
rect 22994 32238 23002 32862
rect 23306 32238 23314 32862
rect 22994 32210 23314 32238
rect 23994 32862 24314 32890
rect 23994 32238 24002 32862
rect 24306 32238 24314 32862
rect 23994 32210 24314 32238
rect 24994 32862 25314 32890
rect 24994 32238 25002 32862
rect 25306 32238 25314 32862
rect 24994 32210 25314 32238
rect 25994 32862 26314 32890
rect 25994 32238 26002 32862
rect 26306 32238 26314 32862
rect 25994 32210 26314 32238
rect 26994 32862 27314 32890
rect 26994 32238 27002 32862
rect 27306 32238 27314 32862
rect 26994 32210 27314 32238
rect 27994 32862 28314 32890
rect 27994 32238 28002 32862
rect 28306 32238 28314 32862
rect 27994 32210 28314 32238
rect 28994 32862 29314 32890
rect 28994 32238 29002 32862
rect 29306 32238 29314 32862
rect 28994 32210 29314 32238
rect 29994 32862 30314 32890
rect 29994 32238 30002 32862
rect 30306 32238 30314 32862
rect 29994 32210 30314 32238
rect 30994 32862 31314 32890
rect 30994 32238 31002 32862
rect 31306 32238 31314 32862
rect 30994 32210 31314 32238
rect 31994 32862 32314 32890
rect 31994 32238 32002 32862
rect 32306 32238 32314 32862
rect 31994 32210 32314 32238
rect 32994 32862 33314 32890
rect 32994 32238 33002 32862
rect 33306 32238 33314 32862
rect 32994 32210 33314 32238
rect 33994 32862 34314 32890
rect 33994 32238 34002 32862
rect 34306 32238 34314 32862
rect 33994 32210 34314 32238
rect -74825 32202 -58825 32210
rect -74825 31898 -74817 32202
rect -74513 31898 -74477 32202
rect -74173 31898 -74137 32202
rect -73513 31898 -73477 32202
rect -73173 31898 -73137 32202
rect -72513 31898 -72477 32202
rect -72173 31898 -72137 32202
rect -71513 31898 -71477 32202
rect -71173 31898 -71137 32202
rect -70513 31898 -70477 32202
rect -70173 31898 -70137 32202
rect -69513 31898 -69477 32202
rect -69173 31898 -69137 32202
rect -68513 31898 -68477 32202
rect -68173 31898 -68137 32202
rect -67513 31898 -67477 32202
rect -67173 31898 -67137 32202
rect -66513 31898 -66477 32202
rect -66173 31898 -66137 32202
rect -65513 31898 -65477 32202
rect -65173 31898 -65137 32202
rect -64513 31898 -64477 32202
rect -64173 31898 -64137 32202
rect -63513 31898 -63477 32202
rect -63173 31898 -63137 32202
rect -62513 31898 -62477 32202
rect -62173 31898 -62137 32202
rect -61513 31898 -61477 32202
rect -61173 31898 -61137 32202
rect -60513 31898 -60477 32202
rect -60173 31898 -60137 32202
rect -59513 31898 -59477 32202
rect -59173 31898 -59137 32202
rect -58833 31898 -58825 32202
rect -74825 31890 -58825 31898
rect 9654 32202 34654 32210
rect 9654 31898 9662 32202
rect 9966 31898 10002 32202
rect 10306 31898 10342 32202
rect 10966 31898 11002 32202
rect 11306 31898 11342 32202
rect 11966 31898 12002 32202
rect 12306 31898 12342 32202
rect 12966 31898 13002 32202
rect 13306 31898 13342 32202
rect 13966 31898 14002 32202
rect 14306 31898 14342 32202
rect 14966 31898 15002 32202
rect 15306 31898 15342 32202
rect 15966 31898 16002 32202
rect 16306 31898 16342 32202
rect 16966 31898 17002 32202
rect 17306 31898 17342 32202
rect 17966 31898 18002 32202
rect 18306 31898 18342 32202
rect 18966 31898 19002 32202
rect 19306 31898 19342 32202
rect 19966 31898 20002 32202
rect 20306 31898 20342 32202
rect 20966 31898 21002 32202
rect 21306 31898 21342 32202
rect 21966 31898 22002 32202
rect 22306 31898 22342 32202
rect 22966 31898 23002 32202
rect 23306 31898 23342 32202
rect 23966 31898 24002 32202
rect 24306 31898 24342 32202
rect 24966 31898 25002 32202
rect 25306 31898 25342 32202
rect 25966 31898 26002 32202
rect 26306 31898 26342 32202
rect 26966 31898 27002 32202
rect 27306 31898 27342 32202
rect 27966 31898 28002 32202
rect 28306 31898 28342 32202
rect 28966 31898 29002 32202
rect 29306 31898 29342 32202
rect 29966 31898 30002 32202
rect 30306 31898 30342 32202
rect 30966 31898 31002 32202
rect 31306 31898 31342 32202
rect 31966 31898 32002 32202
rect 32306 31898 32342 32202
rect 32966 31898 33002 32202
rect 33306 31898 33342 32202
rect 33966 31898 34002 32202
rect 34306 31898 34342 32202
rect 34646 31898 34654 32202
rect 9654 31890 34654 31898
rect -74485 31862 -74165 31890
rect -74485 31238 -74477 31862
rect -74173 31238 -74165 31862
rect -74485 31210 -74165 31238
rect -73485 31862 -73165 31890
rect -73485 31238 -73477 31862
rect -73173 31238 -73165 31862
rect -73485 31210 -73165 31238
rect -72485 31862 -72165 31890
rect -72485 31238 -72477 31862
rect -72173 31238 -72165 31862
rect -72485 31210 -72165 31238
rect -71485 31862 -71165 31890
rect -71485 31238 -71477 31862
rect -71173 31238 -71165 31862
rect -71485 31210 -71165 31238
rect -70485 31862 -70165 31890
rect -70485 31238 -70477 31862
rect -70173 31238 -70165 31862
rect -70485 31210 -70165 31238
rect -69485 31862 -69165 31890
rect -69485 31238 -69477 31862
rect -69173 31238 -69165 31862
rect -69485 31210 -69165 31238
rect -68485 31862 -68165 31890
rect -68485 31238 -68477 31862
rect -68173 31238 -68165 31862
rect -68485 31210 -68165 31238
rect -67485 31862 -67165 31890
rect -67485 31238 -67477 31862
rect -67173 31238 -67165 31862
rect -67485 31210 -67165 31238
rect -66485 31862 -66165 31890
rect -66485 31238 -66477 31862
rect -66173 31238 -66165 31862
rect -66485 31210 -66165 31238
rect -65485 31862 -65165 31890
rect -65485 31238 -65477 31862
rect -65173 31238 -65165 31862
rect -65485 31210 -65165 31238
rect -64485 31862 -64165 31890
rect -64485 31238 -64477 31862
rect -64173 31238 -64165 31862
rect -64485 31210 -64165 31238
rect -63485 31862 -63165 31890
rect -63485 31238 -63477 31862
rect -63173 31238 -63165 31862
rect -63485 31210 -63165 31238
rect -62485 31862 -62165 31890
rect -62485 31238 -62477 31862
rect -62173 31238 -62165 31862
rect -62485 31210 -62165 31238
rect -61485 31862 -61165 31890
rect -61485 31238 -61477 31862
rect -61173 31238 -61165 31862
rect -61485 31210 -61165 31238
rect -60485 31862 -60165 31890
rect -60485 31238 -60477 31862
rect -60173 31238 -60165 31862
rect -60485 31210 -60165 31238
rect -59485 31862 -59165 31890
rect -59485 31238 -59477 31862
rect -59173 31238 -59165 31862
rect -59485 31210 -59165 31238
rect 9994 31862 10314 31890
rect 9994 31238 10002 31862
rect 10306 31238 10314 31862
rect 9994 31210 10314 31238
rect 10994 31862 11314 31890
rect 10994 31238 11002 31862
rect 11306 31238 11314 31862
rect 10994 31210 11314 31238
rect 11994 31862 12314 31890
rect 11994 31238 12002 31862
rect 12306 31238 12314 31862
rect 11994 31210 12314 31238
rect 12994 31862 13314 31890
rect 12994 31238 13002 31862
rect 13306 31238 13314 31862
rect 12994 31210 13314 31238
rect 13994 31862 14314 31890
rect 13994 31238 14002 31862
rect 14306 31238 14314 31862
rect 13994 31210 14314 31238
rect 14994 31862 15314 31890
rect 14994 31238 15002 31862
rect 15306 31238 15314 31862
rect 14994 31210 15314 31238
rect 15994 31862 16314 31890
rect 15994 31238 16002 31862
rect 16306 31238 16314 31862
rect 15994 31210 16314 31238
rect 16994 31862 17314 31890
rect 16994 31238 17002 31862
rect 17306 31238 17314 31862
rect 16994 31210 17314 31238
rect 17994 31862 18314 31890
rect 17994 31238 18002 31862
rect 18306 31238 18314 31862
rect 17994 31210 18314 31238
rect 18994 31862 19314 31890
rect 18994 31238 19002 31862
rect 19306 31238 19314 31862
rect 18994 31210 19314 31238
rect 19994 31862 20314 31890
rect 19994 31238 20002 31862
rect 20306 31238 20314 31862
rect 19994 31210 20314 31238
rect 20994 31862 21314 31890
rect 20994 31238 21002 31862
rect 21306 31238 21314 31862
rect 20994 31210 21314 31238
rect 21994 31862 22314 31890
rect 21994 31238 22002 31862
rect 22306 31238 22314 31862
rect 21994 31210 22314 31238
rect 22994 31862 23314 31890
rect 22994 31238 23002 31862
rect 23306 31238 23314 31862
rect 22994 31210 23314 31238
rect 23994 31862 24314 31890
rect 23994 31238 24002 31862
rect 24306 31238 24314 31862
rect 23994 31210 24314 31238
rect 24994 31862 25314 31890
rect 24994 31238 25002 31862
rect 25306 31238 25314 31862
rect 24994 31210 25314 31238
rect 25994 31862 26314 31890
rect 25994 31238 26002 31862
rect 26306 31238 26314 31862
rect 25994 31210 26314 31238
rect 26994 31862 27314 31890
rect 26994 31238 27002 31862
rect 27306 31238 27314 31862
rect 26994 31210 27314 31238
rect 27994 31862 28314 31890
rect 27994 31238 28002 31862
rect 28306 31238 28314 31862
rect 27994 31210 28314 31238
rect 28994 31862 29314 31890
rect 28994 31238 29002 31862
rect 29306 31238 29314 31862
rect 28994 31210 29314 31238
rect 29994 31862 30314 31890
rect 29994 31238 30002 31862
rect 30306 31238 30314 31862
rect 29994 31210 30314 31238
rect 30994 31862 31314 31890
rect 30994 31238 31002 31862
rect 31306 31238 31314 31862
rect 30994 31210 31314 31238
rect 31994 31862 32314 31890
rect 31994 31238 32002 31862
rect 32306 31238 32314 31862
rect 31994 31210 32314 31238
rect 32994 31862 33314 31890
rect 32994 31238 33002 31862
rect 33306 31238 33314 31862
rect 32994 31210 33314 31238
rect 33994 31862 34314 31890
rect 33994 31238 34002 31862
rect 34306 31238 34314 31862
rect 33994 31210 34314 31238
rect -74825 31202 -58825 31210
rect -74825 30898 -74817 31202
rect -74513 30898 -74477 31202
rect -74173 30898 -74137 31202
rect -73513 30898 -73477 31202
rect -73173 30898 -73137 31202
rect -72513 30898 -72477 31202
rect -72173 30898 -72137 31202
rect -71513 30898 -71477 31202
rect -71173 30898 -71137 31202
rect -70513 30898 -70477 31202
rect -70173 30898 -70137 31202
rect -69513 30898 -69477 31202
rect -69173 30898 -69137 31202
rect -68513 30898 -68477 31202
rect -68173 30898 -68137 31202
rect -67513 30898 -67477 31202
rect -67173 30898 -67137 31202
rect -66513 30898 -66477 31202
rect -66173 30898 -66137 31202
rect -65513 30898 -65477 31202
rect -65173 30898 -65137 31202
rect -64513 30898 -64477 31202
rect -64173 30898 -64137 31202
rect -63513 30898 -63477 31202
rect -63173 30898 -63137 31202
rect -62513 30898 -62477 31202
rect -62173 30898 -62137 31202
rect -61513 30898 -61477 31202
rect -61173 30898 -61137 31202
rect -60513 30898 -60477 31202
rect -60173 30898 -60137 31202
rect -59513 30898 -59477 31202
rect -59173 30898 -59137 31202
rect -58833 30898 -58825 31202
rect -74825 30890 -58825 30898
rect 9654 31202 34654 31210
rect 9654 30898 9662 31202
rect 9966 30898 10002 31202
rect 10306 30898 10342 31202
rect 10966 30898 11002 31202
rect 11306 30898 11342 31202
rect 11966 30898 12002 31202
rect 12306 30898 12342 31202
rect 12966 30898 13002 31202
rect 13306 30898 13342 31202
rect 13966 30898 14002 31202
rect 14306 30898 14342 31202
rect 14966 30898 15002 31202
rect 15306 30898 15342 31202
rect 15966 30898 16002 31202
rect 16306 30898 16342 31202
rect 16966 30898 17002 31202
rect 17306 30898 17342 31202
rect 17966 30898 18002 31202
rect 18306 30898 18342 31202
rect 18966 30898 19002 31202
rect 19306 30898 19342 31202
rect 19966 30898 20002 31202
rect 20306 30898 20342 31202
rect 20966 30898 21002 31202
rect 21306 30898 21342 31202
rect 21966 30898 22002 31202
rect 22306 30898 22342 31202
rect 22966 30898 23002 31202
rect 23306 30898 23342 31202
rect 23966 30898 24002 31202
rect 24306 30898 24342 31202
rect 24966 30898 25002 31202
rect 25306 30898 25342 31202
rect 25966 30898 26002 31202
rect 26306 30898 26342 31202
rect 26966 30898 27002 31202
rect 27306 30898 27342 31202
rect 27966 30898 28002 31202
rect 28306 30898 28342 31202
rect 28966 30898 29002 31202
rect 29306 30898 29342 31202
rect 29966 30898 30002 31202
rect 30306 30898 30342 31202
rect 30966 30898 31002 31202
rect 31306 30898 31342 31202
rect 31966 30898 32002 31202
rect 32306 30898 32342 31202
rect 32966 30898 33002 31202
rect 33306 30898 33342 31202
rect 33966 30898 34002 31202
rect 34306 30898 34342 31202
rect 34646 30898 34654 31202
rect 9654 30890 34654 30898
rect -74485 30862 -74165 30890
rect -74485 30238 -74477 30862
rect -74173 30238 -74165 30862
rect -74485 30210 -74165 30238
rect -73485 30862 -73165 30890
rect -73485 30238 -73477 30862
rect -73173 30238 -73165 30862
rect -73485 30210 -73165 30238
rect -72485 30862 -72165 30890
rect -72485 30238 -72477 30862
rect -72173 30238 -72165 30862
rect -72485 30210 -72165 30238
rect -71485 30862 -71165 30890
rect -71485 30238 -71477 30862
rect -71173 30238 -71165 30862
rect -71485 30210 -71165 30238
rect -70485 30862 -70165 30890
rect -70485 30238 -70477 30862
rect -70173 30238 -70165 30862
rect -70485 30210 -70165 30238
rect -69485 30862 -69165 30890
rect -69485 30238 -69477 30862
rect -69173 30238 -69165 30862
rect -69485 30210 -69165 30238
rect -68485 30862 -68165 30890
rect -68485 30238 -68477 30862
rect -68173 30238 -68165 30862
rect -68485 30210 -68165 30238
rect -67485 30862 -67165 30890
rect -67485 30238 -67477 30862
rect -67173 30238 -67165 30862
rect -67485 30210 -67165 30238
rect -66485 30862 -66165 30890
rect -66485 30238 -66477 30862
rect -66173 30238 -66165 30862
rect -66485 30210 -66165 30238
rect -65485 30862 -65165 30890
rect -65485 30238 -65477 30862
rect -65173 30238 -65165 30862
rect -65485 30210 -65165 30238
rect -64485 30862 -64165 30890
rect -64485 30238 -64477 30862
rect -64173 30238 -64165 30862
rect -64485 30210 -64165 30238
rect -63485 30862 -63165 30890
rect -63485 30238 -63477 30862
rect -63173 30238 -63165 30862
rect -63485 30210 -63165 30238
rect -62485 30862 -62165 30890
rect -62485 30238 -62477 30862
rect -62173 30238 -62165 30862
rect -62485 30210 -62165 30238
rect -61485 30862 -61165 30890
rect -61485 30238 -61477 30862
rect -61173 30238 -61165 30862
rect -61485 30210 -61165 30238
rect -60485 30862 -60165 30890
rect -60485 30238 -60477 30862
rect -60173 30238 -60165 30862
rect -60485 30210 -60165 30238
rect -59485 30862 -59165 30890
rect -59485 30238 -59477 30862
rect -59173 30238 -59165 30862
rect -59485 30210 -59165 30238
rect 9994 30862 10314 30890
rect 9994 30238 10002 30862
rect 10306 30238 10314 30862
rect 9994 30210 10314 30238
rect 10994 30862 11314 30890
rect 10994 30238 11002 30862
rect 11306 30238 11314 30862
rect 10994 30210 11314 30238
rect 11994 30862 12314 30890
rect 11994 30238 12002 30862
rect 12306 30238 12314 30862
rect 11994 30210 12314 30238
rect 12994 30862 13314 30890
rect 12994 30238 13002 30862
rect 13306 30238 13314 30862
rect 12994 30210 13314 30238
rect 13994 30862 14314 30890
rect 13994 30238 14002 30862
rect 14306 30238 14314 30862
rect 13994 30210 14314 30238
rect 14994 30862 15314 30890
rect 14994 30238 15002 30862
rect 15306 30238 15314 30862
rect 14994 30210 15314 30238
rect 15994 30862 16314 30890
rect 15994 30238 16002 30862
rect 16306 30238 16314 30862
rect 15994 30210 16314 30238
rect 16994 30862 17314 30890
rect 16994 30238 17002 30862
rect 17306 30238 17314 30862
rect 16994 30210 17314 30238
rect 17994 30862 18314 30890
rect 17994 30238 18002 30862
rect 18306 30238 18314 30862
rect 17994 30210 18314 30238
rect 18994 30862 19314 30890
rect 18994 30238 19002 30862
rect 19306 30238 19314 30862
rect 18994 30210 19314 30238
rect 19994 30862 20314 30890
rect 19994 30238 20002 30862
rect 20306 30238 20314 30862
rect 19994 30210 20314 30238
rect 20994 30862 21314 30890
rect 20994 30238 21002 30862
rect 21306 30238 21314 30862
rect 20994 30210 21314 30238
rect 21994 30862 22314 30890
rect 21994 30238 22002 30862
rect 22306 30238 22314 30862
rect 21994 30210 22314 30238
rect 22994 30862 23314 30890
rect 22994 30238 23002 30862
rect 23306 30238 23314 30862
rect 22994 30210 23314 30238
rect 23994 30862 24314 30890
rect 23994 30238 24002 30862
rect 24306 30238 24314 30862
rect 23994 30210 24314 30238
rect 24994 30862 25314 30890
rect 24994 30238 25002 30862
rect 25306 30238 25314 30862
rect 24994 30210 25314 30238
rect 25994 30862 26314 30890
rect 25994 30238 26002 30862
rect 26306 30238 26314 30862
rect 25994 30210 26314 30238
rect 26994 30862 27314 30890
rect 26994 30238 27002 30862
rect 27306 30238 27314 30862
rect 26994 30210 27314 30238
rect 27994 30862 28314 30890
rect 27994 30238 28002 30862
rect 28306 30238 28314 30862
rect 27994 30210 28314 30238
rect 28994 30862 29314 30890
rect 28994 30238 29002 30862
rect 29306 30238 29314 30862
rect 28994 30210 29314 30238
rect 29994 30862 30314 30890
rect 29994 30238 30002 30862
rect 30306 30238 30314 30862
rect 29994 30210 30314 30238
rect 30994 30862 31314 30890
rect 30994 30238 31002 30862
rect 31306 30238 31314 30862
rect 30994 30210 31314 30238
rect 31994 30862 32314 30890
rect 31994 30238 32002 30862
rect 32306 30238 32314 30862
rect 31994 30210 32314 30238
rect 32994 30862 33314 30890
rect 32994 30238 33002 30862
rect 33306 30238 33314 30862
rect 32994 30210 33314 30238
rect 33994 30862 34314 30890
rect 33994 30238 34002 30862
rect 34306 30238 34314 30862
rect 33994 30210 34314 30238
rect -74825 30202 -58825 30210
rect -74825 29898 -74817 30202
rect -74513 29898 -74477 30202
rect -74173 29898 -74137 30202
rect -73513 29898 -73477 30202
rect -73173 29898 -73137 30202
rect -72513 29898 -72477 30202
rect -72173 29898 -72137 30202
rect -71513 29898 -71477 30202
rect -71173 29898 -71137 30202
rect -70513 29898 -70477 30202
rect -70173 29898 -70137 30202
rect -69513 29898 -69477 30202
rect -69173 29898 -69137 30202
rect -68513 29898 -68477 30202
rect -68173 29898 -68137 30202
rect -67513 29898 -67477 30202
rect -67173 29898 -67137 30202
rect -66513 29898 -66477 30202
rect -66173 29898 -66137 30202
rect -65513 29898 -65477 30202
rect -65173 29898 -65137 30202
rect -64513 29898 -64477 30202
rect -64173 29898 -64137 30202
rect -63513 29898 -63477 30202
rect -63173 29898 -63137 30202
rect -62513 29898 -62477 30202
rect -62173 29898 -62137 30202
rect -61513 29898 -61477 30202
rect -61173 29898 -61137 30202
rect -60513 29898 -60477 30202
rect -60173 29898 -60137 30202
rect -59513 29898 -59477 30202
rect -59173 29898 -59137 30202
rect -58833 29898 -58825 30202
rect -74825 29890 -58825 29898
rect 9654 30202 34654 30210
rect 9654 29898 9662 30202
rect 9966 29898 10002 30202
rect 10306 29898 10342 30202
rect 10966 29898 11002 30202
rect 11306 29898 11342 30202
rect 11966 29898 12002 30202
rect 12306 29898 12342 30202
rect 12966 29898 13002 30202
rect 13306 29898 13342 30202
rect 13966 29898 14002 30202
rect 14306 29898 14342 30202
rect 14966 29898 15002 30202
rect 15306 29898 15342 30202
rect 15966 29898 16002 30202
rect 16306 29898 16342 30202
rect 16966 29898 17002 30202
rect 17306 29898 17342 30202
rect 17966 29898 18002 30202
rect 18306 29898 18342 30202
rect 18966 29898 19002 30202
rect 19306 29898 19342 30202
rect 19966 29898 20002 30202
rect 20306 29898 20342 30202
rect 20966 29898 21002 30202
rect 21306 29898 21342 30202
rect 21966 29898 22002 30202
rect 22306 29898 22342 30202
rect 22966 29898 23002 30202
rect 23306 29898 23342 30202
rect 23966 29898 24002 30202
rect 24306 29898 24342 30202
rect 24966 29898 25002 30202
rect 25306 29898 25342 30202
rect 25966 29898 26002 30202
rect 26306 29898 26342 30202
rect 26966 29898 27002 30202
rect 27306 29898 27342 30202
rect 27966 29898 28002 30202
rect 28306 29898 28342 30202
rect 28966 29898 29002 30202
rect 29306 29898 29342 30202
rect 29966 29898 30002 30202
rect 30306 29898 30342 30202
rect 30966 29898 31002 30202
rect 31306 29898 31342 30202
rect 31966 29898 32002 30202
rect 32306 29898 32342 30202
rect 32966 29898 33002 30202
rect 33306 29898 33342 30202
rect 33966 29898 34002 30202
rect 34306 29898 34342 30202
rect 34646 29898 34654 30202
rect 9654 29890 34654 29898
rect -74485 29862 -74165 29890
rect -74485 29238 -74477 29862
rect -74173 29238 -74165 29862
rect -74485 29210 -74165 29238
rect -73485 29862 -73165 29890
rect -73485 29238 -73477 29862
rect -73173 29238 -73165 29862
rect -73485 29210 -73165 29238
rect -72485 29862 -72165 29890
rect -72485 29238 -72477 29862
rect -72173 29238 -72165 29862
rect -72485 29210 -72165 29238
rect -71485 29862 -71165 29890
rect -71485 29238 -71477 29862
rect -71173 29238 -71165 29862
rect -71485 29210 -71165 29238
rect -70485 29862 -70165 29890
rect -70485 29238 -70477 29862
rect -70173 29238 -70165 29862
rect -70485 29210 -70165 29238
rect -69485 29862 -69165 29890
rect -69485 29238 -69477 29862
rect -69173 29238 -69165 29862
rect -69485 29210 -69165 29238
rect -68485 29862 -68165 29890
rect -68485 29238 -68477 29862
rect -68173 29238 -68165 29862
rect -68485 29210 -68165 29238
rect -67485 29862 -67165 29890
rect -67485 29238 -67477 29862
rect -67173 29238 -67165 29862
rect -67485 29210 -67165 29238
rect -66485 29862 -66165 29890
rect -66485 29238 -66477 29862
rect -66173 29238 -66165 29862
rect -66485 29210 -66165 29238
rect -65485 29862 -65165 29890
rect -65485 29238 -65477 29862
rect -65173 29238 -65165 29862
rect -65485 29210 -65165 29238
rect -64485 29862 -64165 29890
rect -64485 29238 -64477 29862
rect -64173 29238 -64165 29862
rect -64485 29210 -64165 29238
rect -63485 29862 -63165 29890
rect -63485 29238 -63477 29862
rect -63173 29238 -63165 29862
rect -63485 29210 -63165 29238
rect -62485 29862 -62165 29890
rect -62485 29238 -62477 29862
rect -62173 29238 -62165 29862
rect -62485 29210 -62165 29238
rect -61485 29862 -61165 29890
rect -61485 29238 -61477 29862
rect -61173 29238 -61165 29862
rect -61485 29210 -61165 29238
rect -60485 29862 -60165 29890
rect -60485 29238 -60477 29862
rect -60173 29238 -60165 29862
rect -60485 29210 -60165 29238
rect -59485 29862 -59165 29890
rect -59485 29238 -59477 29862
rect -59173 29238 -59165 29862
rect -59485 29210 -59165 29238
rect 9994 29862 10314 29890
rect 9994 29238 10002 29862
rect 10306 29238 10314 29862
rect 9994 29210 10314 29238
rect 10994 29862 11314 29890
rect 10994 29238 11002 29862
rect 11306 29238 11314 29862
rect 10994 29210 11314 29238
rect 11994 29862 12314 29890
rect 11994 29238 12002 29862
rect 12306 29238 12314 29862
rect 11994 29210 12314 29238
rect 12994 29862 13314 29890
rect 12994 29238 13002 29862
rect 13306 29238 13314 29862
rect 12994 29210 13314 29238
rect 13994 29862 14314 29890
rect 13994 29238 14002 29862
rect 14306 29238 14314 29862
rect 13994 29210 14314 29238
rect 14994 29862 15314 29890
rect 14994 29238 15002 29862
rect 15306 29238 15314 29862
rect 14994 29210 15314 29238
rect 15994 29862 16314 29890
rect 15994 29238 16002 29862
rect 16306 29238 16314 29862
rect 15994 29210 16314 29238
rect 16994 29862 17314 29890
rect 16994 29238 17002 29862
rect 17306 29238 17314 29862
rect 16994 29210 17314 29238
rect 17994 29862 18314 29890
rect 17994 29238 18002 29862
rect 18306 29238 18314 29862
rect 17994 29210 18314 29238
rect 18994 29862 19314 29890
rect 18994 29238 19002 29862
rect 19306 29238 19314 29862
rect 18994 29210 19314 29238
rect 19994 29862 20314 29890
rect 19994 29238 20002 29862
rect 20306 29238 20314 29862
rect 19994 29210 20314 29238
rect 20994 29862 21314 29890
rect 20994 29238 21002 29862
rect 21306 29238 21314 29862
rect 20994 29210 21314 29238
rect 21994 29862 22314 29890
rect 21994 29238 22002 29862
rect 22306 29238 22314 29862
rect 21994 29210 22314 29238
rect 22994 29862 23314 29890
rect 22994 29238 23002 29862
rect 23306 29238 23314 29862
rect 22994 29210 23314 29238
rect 23994 29862 24314 29890
rect 23994 29238 24002 29862
rect 24306 29238 24314 29862
rect 23994 29210 24314 29238
rect 24994 29862 25314 29890
rect 24994 29238 25002 29862
rect 25306 29238 25314 29862
rect 24994 29210 25314 29238
rect 25994 29862 26314 29890
rect 25994 29238 26002 29862
rect 26306 29238 26314 29862
rect 25994 29210 26314 29238
rect 26994 29862 27314 29890
rect 26994 29238 27002 29862
rect 27306 29238 27314 29862
rect 26994 29210 27314 29238
rect 27994 29862 28314 29890
rect 27994 29238 28002 29862
rect 28306 29238 28314 29862
rect 27994 29210 28314 29238
rect 28994 29862 29314 29890
rect 28994 29238 29002 29862
rect 29306 29238 29314 29862
rect 28994 29210 29314 29238
rect 29994 29862 30314 29890
rect 29994 29238 30002 29862
rect 30306 29238 30314 29862
rect 29994 29210 30314 29238
rect 30994 29862 31314 29890
rect 30994 29238 31002 29862
rect 31306 29238 31314 29862
rect 30994 29210 31314 29238
rect 31994 29862 32314 29890
rect 31994 29238 32002 29862
rect 32306 29238 32314 29862
rect 31994 29210 32314 29238
rect 32994 29862 33314 29890
rect 32994 29238 33002 29862
rect 33306 29238 33314 29862
rect 32994 29210 33314 29238
rect 33994 29862 34314 29890
rect 33994 29238 34002 29862
rect 34306 29238 34314 29862
rect 33994 29210 34314 29238
rect -74825 29202 -58825 29210
rect -74825 28898 -74817 29202
rect -74513 28898 -74477 29202
rect -74173 28898 -74137 29202
rect -73513 28898 -73477 29202
rect -73173 28898 -73137 29202
rect -72513 28898 -72477 29202
rect -72173 28898 -72137 29202
rect -71513 28898 -71477 29202
rect -71173 28898 -71137 29202
rect -70513 28898 -70477 29202
rect -70173 28898 -70137 29202
rect -69513 28898 -69477 29202
rect -69173 28898 -69137 29202
rect -68513 28898 -68477 29202
rect -68173 28898 -68137 29202
rect -67513 28898 -67477 29202
rect -67173 28898 -67137 29202
rect -66513 28898 -66477 29202
rect -66173 28898 -66137 29202
rect -65513 28898 -65477 29202
rect -65173 28898 -65137 29202
rect -64513 28898 -64477 29202
rect -64173 28898 -64137 29202
rect -63513 28898 -63477 29202
rect -63173 28898 -63137 29202
rect -62513 28898 -62477 29202
rect -62173 28898 -62137 29202
rect -61513 28898 -61477 29202
rect -61173 28898 -61137 29202
rect -60513 28898 -60477 29202
rect -60173 28898 -60137 29202
rect -59513 28898 -59477 29202
rect -59173 28898 -59137 29202
rect -58833 28898 -58825 29202
rect -74825 28890 -58825 28898
rect 9654 29202 34654 29210
rect 9654 28898 9662 29202
rect 9966 28898 10002 29202
rect 10306 28898 10342 29202
rect 10966 28898 11002 29202
rect 11306 28898 11342 29202
rect 11966 28898 12002 29202
rect 12306 28898 12342 29202
rect 12966 28898 13002 29202
rect 13306 28898 13342 29202
rect 13966 28898 14002 29202
rect 14306 28898 14342 29202
rect 14966 28898 15002 29202
rect 15306 28898 15342 29202
rect 15966 28898 16002 29202
rect 16306 28898 16342 29202
rect 16966 28898 17002 29202
rect 17306 28898 17342 29202
rect 17966 28898 18002 29202
rect 18306 28898 18342 29202
rect 18966 28898 19002 29202
rect 19306 28898 19342 29202
rect 19966 28898 20002 29202
rect 20306 28898 20342 29202
rect 20966 28898 21002 29202
rect 21306 28898 21342 29202
rect 21966 28898 22002 29202
rect 22306 28898 22342 29202
rect 22966 28898 23002 29202
rect 23306 28898 23342 29202
rect 23966 28898 24002 29202
rect 24306 28898 24342 29202
rect 24966 28898 25002 29202
rect 25306 28898 25342 29202
rect 25966 28898 26002 29202
rect 26306 28898 26342 29202
rect 26966 28898 27002 29202
rect 27306 28898 27342 29202
rect 27966 28898 28002 29202
rect 28306 28898 28342 29202
rect 28966 28898 29002 29202
rect 29306 28898 29342 29202
rect 29966 28898 30002 29202
rect 30306 28898 30342 29202
rect 30966 28898 31002 29202
rect 31306 28898 31342 29202
rect 31966 28898 32002 29202
rect 32306 28898 32342 29202
rect 32966 28898 33002 29202
rect 33306 28898 33342 29202
rect 33966 28898 34002 29202
rect 34306 28898 34342 29202
rect 34646 28898 34654 29202
rect 9654 28890 34654 28898
rect -74485 28862 -74165 28890
rect -74485 28558 -74477 28862
rect -74173 28558 -74165 28862
rect -74485 28550 -74165 28558
rect -73485 28862 -73165 28890
rect -73485 28558 -73477 28862
rect -73173 28558 -73165 28862
rect -73485 28550 -73165 28558
rect -72485 28862 -72165 28890
rect -72485 28558 -72477 28862
rect -72173 28558 -72165 28862
rect -72485 28550 -72165 28558
rect -71485 28862 -71165 28890
rect -71485 28558 -71477 28862
rect -71173 28558 -71165 28862
rect -71485 28550 -71165 28558
rect -70485 28862 -70165 28890
rect -70485 28558 -70477 28862
rect -70173 28558 -70165 28862
rect -70485 28550 -70165 28558
rect -69485 28862 -69165 28890
rect -69485 28558 -69477 28862
rect -69173 28558 -69165 28862
rect -69485 28550 -69165 28558
rect -68485 28862 -68165 28890
rect -68485 28558 -68477 28862
rect -68173 28558 -68165 28862
rect -68485 28550 -68165 28558
rect -67485 28862 -67165 28890
rect -67485 28558 -67477 28862
rect -67173 28558 -67165 28862
rect -67485 28550 -67165 28558
rect -66485 28862 -66165 28890
rect -66485 28558 -66477 28862
rect -66173 28558 -66165 28862
rect -66485 28550 -66165 28558
rect -65485 28862 -65165 28890
rect -65485 28558 -65477 28862
rect -65173 28558 -65165 28862
rect -65485 28550 -65165 28558
rect -64485 28862 -64165 28890
rect -64485 28558 -64477 28862
rect -64173 28558 -64165 28862
rect -64485 28550 -64165 28558
rect -63485 28862 -63165 28890
rect -63485 28558 -63477 28862
rect -63173 28558 -63165 28862
rect -63485 28550 -63165 28558
rect -62485 28862 -62165 28890
rect -62485 28558 -62477 28862
rect -62173 28558 -62165 28862
rect -62485 28550 -62165 28558
rect -61485 28862 -61165 28890
rect -61485 28558 -61477 28862
rect -61173 28558 -61165 28862
rect -61485 28550 -61165 28558
rect -60485 28862 -60165 28890
rect -60485 28558 -60477 28862
rect -60173 28558 -60165 28862
rect -60485 28550 -60165 28558
rect -59485 28862 -59165 28890
rect -59485 28558 -59477 28862
rect -59173 28558 -59165 28862
rect -59485 28550 -59165 28558
rect 9994 28862 10314 28890
rect 9994 28558 10002 28862
rect 10306 28558 10314 28862
rect 9994 28550 10314 28558
rect 10994 28862 11314 28890
rect 10994 28558 11002 28862
rect 11306 28558 11314 28862
rect 10994 28550 11314 28558
rect 11994 28862 12314 28890
rect 11994 28558 12002 28862
rect 12306 28558 12314 28862
rect 11994 28550 12314 28558
rect 12994 28862 13314 28890
rect 12994 28558 13002 28862
rect 13306 28558 13314 28862
rect 12994 28550 13314 28558
rect 13994 28862 14314 28890
rect 13994 28558 14002 28862
rect 14306 28558 14314 28862
rect 13994 28550 14314 28558
rect 14994 28862 15314 28890
rect 14994 28558 15002 28862
rect 15306 28558 15314 28862
rect 14994 28550 15314 28558
rect 15994 28862 16314 28890
rect 15994 28558 16002 28862
rect 16306 28558 16314 28862
rect 15994 28550 16314 28558
rect 16994 28862 17314 28890
rect 16994 28558 17002 28862
rect 17306 28558 17314 28862
rect 16994 28550 17314 28558
rect 17994 28862 18314 28890
rect 17994 28558 18002 28862
rect 18306 28558 18314 28862
rect 17994 28550 18314 28558
rect 18994 28862 19314 28890
rect 18994 28558 19002 28862
rect 19306 28558 19314 28862
rect 18994 28550 19314 28558
rect 19994 28862 20314 28890
rect 19994 28558 20002 28862
rect 20306 28558 20314 28862
rect 19994 28550 20314 28558
rect 20994 28862 21314 28890
rect 20994 28558 21002 28862
rect 21306 28558 21314 28862
rect 20994 28550 21314 28558
rect 21994 28862 22314 28890
rect 21994 28558 22002 28862
rect 22306 28558 22314 28862
rect 21994 28550 22314 28558
rect 22994 28862 23314 28890
rect 22994 28558 23002 28862
rect 23306 28558 23314 28862
rect 22994 28550 23314 28558
rect 23994 28862 24314 28890
rect 23994 28558 24002 28862
rect 24306 28558 24314 28862
rect 23994 28550 24314 28558
rect 24994 28862 25314 28890
rect 24994 28558 25002 28862
rect 25306 28558 25314 28862
rect 24994 28550 25314 28558
rect 25994 28862 26314 28890
rect 25994 28558 26002 28862
rect 26306 28558 26314 28862
rect 25994 28550 26314 28558
rect 26994 28862 27314 28890
rect 26994 28558 27002 28862
rect 27306 28558 27314 28862
rect 26994 28550 27314 28558
rect 27994 28862 28314 28890
rect 27994 28558 28002 28862
rect 28306 28558 28314 28862
rect 27994 28550 28314 28558
rect 28994 28862 29314 28890
rect 28994 28558 29002 28862
rect 29306 28558 29314 28862
rect 28994 28550 29314 28558
rect 29994 28862 30314 28890
rect 29994 28558 30002 28862
rect 30306 28558 30314 28862
rect 29994 28550 30314 28558
rect 30994 28862 31314 28890
rect 30994 28558 31002 28862
rect 31306 28558 31314 28862
rect 30994 28550 31314 28558
rect 31994 28862 32314 28890
rect 31994 28558 32002 28862
rect 32306 28558 32314 28862
rect 31994 28550 32314 28558
rect 32994 28862 33314 28890
rect 32994 28558 33002 28862
rect 33306 28558 33314 28862
rect 32994 28550 33314 28558
rect 33994 28862 34314 28890
rect 33994 28558 34002 28862
rect 34306 28558 34314 28862
rect 33994 28550 34314 28558
rect -72825 25947 -60825 26000
rect -72825 16043 -72782 25947
rect -60878 16043 -60825 25947
rect -72825 16000 -60825 16043
rect 20275 25952 32275 26000
rect 20275 16048 20318 25952
rect 32222 16048 32275 25952
rect 20275 16000 32275 16048
rect -21216 15122 -19300 15128
rect -21216 13858 -21210 15122
rect -19306 13858 -19300 15122
rect -21216 13850 -19300 13858
rect -42440 13802 -40660 13850
rect -42440 7898 -42382 13802
rect -40718 7898 -40660 13802
rect -42440 7850 -40660 7898
rect -24275 13688 -16275 13850
rect -24275 8012 -24233 13688
rect -16317 8012 -16275 13688
rect -42440 2312 -40660 2350
rect -42440 -2312 -42382 2312
rect -40718 -2312 -40660 2312
rect -42440 -2350 -40660 -2312
rect -24275 -7850 -16275 8012
rect 110 13802 1890 13850
rect 110 7898 168 13802
rect 1832 7898 1890 13802
rect 110 7850 1890 7898
rect 110 2312 1890 2350
rect 110 -2312 168 2312
rect 1832 -2312 1890 2312
rect 110 -2350 1890 -2312
rect -42440 -7898 -40660 -7850
rect -42440 -13802 -42382 -7898
rect -40718 -13802 -40660 -7898
rect -42440 -13850 -40660 -13802
rect -29525 -8017 -11025 -7850
rect -29525 -13693 -29423 -8017
rect -28227 -8026 -11025 -8017
rect -28227 -13693 -12323 -8026
rect -29525 -13702 -12323 -13693
rect -11127 -13702 -11025 -8026
rect -29525 -13850 -11025 -13702
rect 110 -7898 1890 -7850
rect 110 -13802 168 -7898
rect 1832 -13802 1890 -7898
rect 110 -13850 1890 -13802
rect -72825 -16048 -60825 -16000
rect -72825 -25952 -72782 -16048
rect -60878 -25952 -60825 -16048
rect -72825 -26000 -60825 -25952
rect 20275 -16048 32275 -16000
rect 20275 -25952 20318 -16048
rect 32222 -25952 32275 -16048
rect 20275 -26000 32275 -25952
rect -74485 -28558 -74165 -28550
rect -74485 -28862 -74477 -28558
rect -74173 -28862 -74165 -28558
rect -74485 -28890 -74165 -28862
rect -73485 -28558 -73165 -28550
rect -73485 -28862 -73477 -28558
rect -73173 -28862 -73165 -28558
rect -73485 -28890 -73165 -28862
rect -72485 -28558 -72165 -28550
rect -72485 -28862 -72477 -28558
rect -72173 -28862 -72165 -28558
rect -72485 -28890 -72165 -28862
rect -71485 -28558 -71165 -28550
rect -71485 -28862 -71477 -28558
rect -71173 -28862 -71165 -28558
rect -71485 -28890 -71165 -28862
rect -70485 -28558 -70165 -28550
rect -70485 -28862 -70477 -28558
rect -70173 -28862 -70165 -28558
rect -70485 -28890 -70165 -28862
rect -69485 -28558 -69165 -28550
rect -69485 -28862 -69477 -28558
rect -69173 -28862 -69165 -28558
rect -69485 -28890 -69165 -28862
rect -68485 -28558 -68165 -28550
rect -68485 -28862 -68477 -28558
rect -68173 -28862 -68165 -28558
rect -68485 -28890 -68165 -28862
rect -67485 -28558 -67165 -28550
rect -67485 -28862 -67477 -28558
rect -67173 -28862 -67165 -28558
rect -67485 -28890 -67165 -28862
rect -66485 -28558 -66165 -28550
rect -66485 -28862 -66477 -28558
rect -66173 -28862 -66165 -28558
rect -66485 -28890 -66165 -28862
rect -65485 -28558 -65165 -28550
rect -65485 -28862 -65477 -28558
rect -65173 -28862 -65165 -28558
rect -65485 -28890 -65165 -28862
rect -64485 -28558 -64165 -28550
rect -64485 -28862 -64477 -28558
rect -64173 -28862 -64165 -28558
rect -64485 -28890 -64165 -28862
rect -63485 -28558 -63165 -28550
rect -63485 -28862 -63477 -28558
rect -63173 -28862 -63165 -28558
rect -63485 -28890 -63165 -28862
rect -62485 -28558 -62165 -28550
rect -62485 -28862 -62477 -28558
rect -62173 -28862 -62165 -28558
rect -62485 -28890 -62165 -28862
rect -61485 -28558 -61165 -28550
rect -61485 -28862 -61477 -28558
rect -61173 -28862 -61165 -28558
rect -61485 -28890 -61165 -28862
rect -60485 -28558 -60165 -28550
rect -60485 -28862 -60477 -28558
rect -60173 -28862 -60165 -28558
rect -60485 -28890 -60165 -28862
rect -59485 -28558 -59165 -28550
rect -59485 -28862 -59477 -28558
rect -59173 -28862 -59165 -28558
rect -59485 -28890 -59165 -28862
rect -58485 -28558 -58165 -28550
rect -58485 -28862 -58477 -28558
rect -58173 -28862 -58165 -28558
rect -58485 -28890 -58165 -28862
rect -57485 -28558 -57165 -28550
rect -57485 -28862 -57477 -28558
rect -57173 -28862 -57165 -28558
rect -57485 -28890 -57165 -28862
rect -56485 -28558 -56165 -28550
rect -56485 -28862 -56477 -28558
rect -56173 -28862 -56165 -28558
rect -56485 -28890 -56165 -28862
rect -55485 -28558 -55165 -28550
rect -55485 -28862 -55477 -28558
rect -55173 -28862 -55165 -28558
rect -55485 -28890 -55165 -28862
rect -54485 -28558 -54165 -28550
rect -54485 -28862 -54477 -28558
rect -54173 -28862 -54165 -28558
rect -54485 -28890 -54165 -28862
rect -53485 -28558 -53165 -28550
rect -53485 -28862 -53477 -28558
rect -53173 -28862 -53165 -28558
rect -53485 -28890 -53165 -28862
rect -52485 -28558 -52165 -28550
rect -52485 -28862 -52477 -28558
rect -52173 -28862 -52165 -28558
rect -52485 -28890 -52165 -28862
rect -51485 -28558 -51165 -28550
rect -51485 -28862 -51477 -28558
rect -51173 -28862 -51165 -28558
rect -51485 -28890 -51165 -28862
rect -50485 -28558 -50165 -28550
rect -50485 -28862 -50477 -28558
rect -50173 -28862 -50165 -28558
rect -50485 -28890 -50165 -28862
rect -49485 -28558 -49165 -28550
rect -49485 -28862 -49477 -28558
rect -49173 -28862 -49165 -28558
rect -49485 -28890 -49165 -28862
rect 8615 -28558 8935 -28550
rect 8615 -28862 8623 -28558
rect 8927 -28862 8935 -28558
rect 8615 -28890 8935 -28862
rect 9615 -28558 9935 -28550
rect 9615 -28862 9623 -28558
rect 9927 -28862 9935 -28558
rect 9615 -28890 9935 -28862
rect 10615 -28558 10935 -28550
rect 10615 -28862 10623 -28558
rect 10927 -28862 10935 -28558
rect 10615 -28890 10935 -28862
rect 11615 -28558 11935 -28550
rect 11615 -28862 11623 -28558
rect 11927 -28862 11935 -28558
rect 11615 -28890 11935 -28862
rect 12615 -28558 12935 -28550
rect 12615 -28862 12623 -28558
rect 12927 -28862 12935 -28558
rect 12615 -28890 12935 -28862
rect 13615 -28558 13935 -28550
rect 13615 -28862 13623 -28558
rect 13927 -28862 13935 -28558
rect 13615 -28890 13935 -28862
rect 14615 -28558 14935 -28550
rect 14615 -28862 14623 -28558
rect 14927 -28862 14935 -28558
rect 14615 -28890 14935 -28862
rect 15615 -28558 15935 -28550
rect 15615 -28862 15623 -28558
rect 15927 -28862 15935 -28558
rect 15615 -28890 15935 -28862
rect 16615 -28558 16935 -28550
rect 16615 -28862 16623 -28558
rect 16927 -28862 16935 -28558
rect 16615 -28890 16935 -28862
rect 17615 -28558 17935 -28550
rect 17615 -28862 17623 -28558
rect 17927 -28862 17935 -28558
rect 17615 -28890 17935 -28862
rect 18615 -28558 18935 -28550
rect 18615 -28862 18623 -28558
rect 18927 -28862 18935 -28558
rect 18615 -28890 18935 -28862
rect 19615 -28558 19935 -28550
rect 19615 -28862 19623 -28558
rect 19927 -28862 19935 -28558
rect 19615 -28890 19935 -28862
rect 20615 -28558 20935 -28550
rect 20615 -28862 20623 -28558
rect 20927 -28862 20935 -28558
rect 20615 -28890 20935 -28862
rect 21615 -28558 21935 -28550
rect 21615 -28862 21623 -28558
rect 21927 -28862 21935 -28558
rect 21615 -28890 21935 -28862
rect 22615 -28558 22935 -28550
rect 22615 -28862 22623 -28558
rect 22927 -28862 22935 -28558
rect 22615 -28890 22935 -28862
rect 23615 -28558 23935 -28550
rect 23615 -28862 23623 -28558
rect 23927 -28862 23935 -28558
rect 23615 -28890 23935 -28862
rect 24615 -28558 24935 -28550
rect 24615 -28862 24623 -28558
rect 24927 -28862 24935 -28558
rect 24615 -28890 24935 -28862
rect 25615 -28558 25935 -28550
rect 25615 -28862 25623 -28558
rect 25927 -28862 25935 -28558
rect 25615 -28890 25935 -28862
rect 26615 -28558 26935 -28550
rect 26615 -28862 26623 -28558
rect 26927 -28862 26935 -28558
rect 26615 -28890 26935 -28862
rect 27615 -28558 27935 -28550
rect 27615 -28862 27623 -28558
rect 27927 -28862 27935 -28558
rect 27615 -28890 27935 -28862
rect 28615 -28558 28935 -28550
rect 28615 -28862 28623 -28558
rect 28927 -28862 28935 -28558
rect 28615 -28890 28935 -28862
rect 29615 -28558 29935 -28550
rect 29615 -28862 29623 -28558
rect 29927 -28862 29935 -28558
rect 29615 -28890 29935 -28862
rect 30615 -28558 30935 -28550
rect 30615 -28862 30623 -28558
rect 30927 -28862 30935 -28558
rect 30615 -28890 30935 -28862
rect 31615 -28558 31935 -28550
rect 31615 -28862 31623 -28558
rect 31927 -28862 31935 -28558
rect 31615 -28890 31935 -28862
rect 32615 -28558 32935 -28550
rect 32615 -28862 32623 -28558
rect 32927 -28862 32935 -28558
rect 32615 -28890 32935 -28862
rect 33615 -28558 33935 -28550
rect 33615 -28862 33623 -28558
rect 33927 -28862 33935 -28558
rect 33615 -28890 33935 -28862
rect -74825 -28898 -48825 -28890
rect -74825 -29202 -74817 -28898
rect -74513 -29202 -74477 -28898
rect -74173 -29202 -74137 -28898
rect -73513 -29202 -73477 -28898
rect -73173 -29202 -73137 -28898
rect -72513 -29202 -72477 -28898
rect -72173 -29202 -72137 -28898
rect -71513 -29202 -71477 -28898
rect -71173 -29202 -71137 -28898
rect -70513 -29202 -70477 -28898
rect -70173 -29202 -70137 -28898
rect -69513 -29202 -69477 -28898
rect -69173 -29202 -69137 -28898
rect -68513 -29202 -68477 -28898
rect -68173 -29202 -68137 -28898
rect -67513 -29202 -67477 -28898
rect -67173 -29202 -67137 -28898
rect -66513 -29202 -66477 -28898
rect -66173 -29202 -66137 -28898
rect -65513 -29202 -65477 -28898
rect -65173 -29202 -65137 -28898
rect -64513 -29202 -64477 -28898
rect -64173 -29202 -64137 -28898
rect -63513 -29202 -63477 -28898
rect -63173 -29202 -63137 -28898
rect -62513 -29202 -62477 -28898
rect -62173 -29202 -62137 -28898
rect -61513 -29202 -61477 -28898
rect -61173 -29202 -61137 -28898
rect -60513 -29202 -60477 -28898
rect -60173 -29202 -60137 -28898
rect -59513 -29202 -59477 -28898
rect -59173 -29202 -59137 -28898
rect -58513 -29202 -58477 -28898
rect -58173 -29202 -58137 -28898
rect -57513 -29202 -57477 -28898
rect -57173 -29202 -57137 -28898
rect -56513 -29202 -56477 -28898
rect -56173 -29202 -56137 -28898
rect -55513 -29202 -55477 -28898
rect -55173 -29202 -55137 -28898
rect -54513 -29202 -54477 -28898
rect -54173 -29202 -54137 -28898
rect -53513 -29202 -53477 -28898
rect -53173 -29202 -53137 -28898
rect -52513 -29202 -52477 -28898
rect -52173 -29202 -52137 -28898
rect -51513 -29202 -51477 -28898
rect -51173 -29202 -51137 -28898
rect -50513 -29202 -50477 -28898
rect -50173 -29202 -50137 -28898
rect -49513 -29202 -49477 -28898
rect -49173 -29202 -49137 -28898
rect -48833 -29202 -48825 -28898
rect -74825 -29210 -48825 -29202
rect 8275 -28898 34275 -28890
rect 8275 -29202 8283 -28898
rect 8587 -29202 8623 -28898
rect 8927 -29202 8963 -28898
rect 9587 -29202 9623 -28898
rect 9927 -29202 9963 -28898
rect 10587 -29202 10623 -28898
rect 10927 -29202 10963 -28898
rect 11587 -29202 11623 -28898
rect 11927 -29202 11963 -28898
rect 12587 -29202 12623 -28898
rect 12927 -29202 12963 -28898
rect 13587 -29202 13623 -28898
rect 13927 -29202 13963 -28898
rect 14587 -29202 14623 -28898
rect 14927 -29202 14963 -28898
rect 15587 -29202 15623 -28898
rect 15927 -29202 15963 -28898
rect 16587 -29202 16623 -28898
rect 16927 -29202 16963 -28898
rect 17587 -29202 17623 -28898
rect 17927 -29202 17963 -28898
rect 18587 -29202 18623 -28898
rect 18927 -29202 18963 -28898
rect 19587 -29202 19623 -28898
rect 19927 -29202 19963 -28898
rect 20587 -29202 20623 -28898
rect 20927 -29202 20963 -28898
rect 21587 -29202 21623 -28898
rect 21927 -29202 21963 -28898
rect 22587 -29202 22623 -28898
rect 22927 -29202 22963 -28898
rect 23587 -29202 23623 -28898
rect 23927 -29202 23963 -28898
rect 24587 -29202 24623 -28898
rect 24927 -29202 24963 -28898
rect 25587 -29202 25623 -28898
rect 25927 -29202 25963 -28898
rect 26587 -29202 26623 -28898
rect 26927 -29202 26963 -28898
rect 27587 -29202 27623 -28898
rect 27927 -29202 27963 -28898
rect 28587 -29202 28623 -28898
rect 28927 -29202 28963 -28898
rect 29587 -29202 29623 -28898
rect 29927 -29202 29963 -28898
rect 30587 -29202 30623 -28898
rect 30927 -29202 30963 -28898
rect 31587 -29202 31623 -28898
rect 31927 -29202 31963 -28898
rect 32587 -29202 32623 -28898
rect 32927 -29202 32963 -28898
rect 33587 -29202 33623 -28898
rect 33927 -29202 33963 -28898
rect 34267 -29202 34275 -28898
rect 8275 -29210 34275 -29202
rect -74485 -29238 -74165 -29210
rect -74485 -29862 -74477 -29238
rect -74173 -29862 -74165 -29238
rect -74485 -29890 -74165 -29862
rect -73485 -29238 -73165 -29210
rect -73485 -29862 -73477 -29238
rect -73173 -29862 -73165 -29238
rect -73485 -29890 -73165 -29862
rect -72485 -29238 -72165 -29210
rect -72485 -29862 -72477 -29238
rect -72173 -29862 -72165 -29238
rect -72485 -29890 -72165 -29862
rect -71485 -29238 -71165 -29210
rect -71485 -29862 -71477 -29238
rect -71173 -29862 -71165 -29238
rect -71485 -29890 -71165 -29862
rect -70485 -29238 -70165 -29210
rect -70485 -29862 -70477 -29238
rect -70173 -29862 -70165 -29238
rect -70485 -29890 -70165 -29862
rect -69485 -29238 -69165 -29210
rect -69485 -29862 -69477 -29238
rect -69173 -29862 -69165 -29238
rect -69485 -29890 -69165 -29862
rect -68485 -29238 -68165 -29210
rect -68485 -29862 -68477 -29238
rect -68173 -29862 -68165 -29238
rect -68485 -29890 -68165 -29862
rect -67485 -29238 -67165 -29210
rect -67485 -29862 -67477 -29238
rect -67173 -29862 -67165 -29238
rect -67485 -29890 -67165 -29862
rect -66485 -29238 -66165 -29210
rect -66485 -29862 -66477 -29238
rect -66173 -29862 -66165 -29238
rect -66485 -29890 -66165 -29862
rect -65485 -29238 -65165 -29210
rect -65485 -29862 -65477 -29238
rect -65173 -29862 -65165 -29238
rect -65485 -29890 -65165 -29862
rect -64485 -29238 -64165 -29210
rect -64485 -29862 -64477 -29238
rect -64173 -29862 -64165 -29238
rect -64485 -29890 -64165 -29862
rect -63485 -29238 -63165 -29210
rect -63485 -29862 -63477 -29238
rect -63173 -29862 -63165 -29238
rect -63485 -29890 -63165 -29862
rect -62485 -29238 -62165 -29210
rect -62485 -29862 -62477 -29238
rect -62173 -29862 -62165 -29238
rect -62485 -29890 -62165 -29862
rect -61485 -29238 -61165 -29210
rect -61485 -29862 -61477 -29238
rect -61173 -29862 -61165 -29238
rect -61485 -29890 -61165 -29862
rect -60485 -29238 -60165 -29210
rect -60485 -29862 -60477 -29238
rect -60173 -29862 -60165 -29238
rect -60485 -29890 -60165 -29862
rect -59485 -29238 -59165 -29210
rect -59485 -29862 -59477 -29238
rect -59173 -29862 -59165 -29238
rect -59485 -29890 -59165 -29862
rect -58485 -29238 -58165 -29210
rect -58485 -29862 -58477 -29238
rect -58173 -29862 -58165 -29238
rect -58485 -29890 -58165 -29862
rect -57485 -29238 -57165 -29210
rect -57485 -29862 -57477 -29238
rect -57173 -29862 -57165 -29238
rect -57485 -29890 -57165 -29862
rect -56485 -29238 -56165 -29210
rect -56485 -29862 -56477 -29238
rect -56173 -29862 -56165 -29238
rect -56485 -29890 -56165 -29862
rect -55485 -29238 -55165 -29210
rect -55485 -29862 -55477 -29238
rect -55173 -29862 -55165 -29238
rect -55485 -29890 -55165 -29862
rect -54485 -29238 -54165 -29210
rect -54485 -29862 -54477 -29238
rect -54173 -29862 -54165 -29238
rect -54485 -29890 -54165 -29862
rect -53485 -29238 -53165 -29210
rect -53485 -29862 -53477 -29238
rect -53173 -29862 -53165 -29238
rect -53485 -29890 -53165 -29862
rect -52485 -29238 -52165 -29210
rect -52485 -29862 -52477 -29238
rect -52173 -29862 -52165 -29238
rect -52485 -29890 -52165 -29862
rect -51485 -29238 -51165 -29210
rect -51485 -29862 -51477 -29238
rect -51173 -29862 -51165 -29238
rect -51485 -29890 -51165 -29862
rect -50485 -29238 -50165 -29210
rect -50485 -29862 -50477 -29238
rect -50173 -29862 -50165 -29238
rect -50485 -29890 -50165 -29862
rect -49485 -29238 -49165 -29210
rect -49485 -29862 -49477 -29238
rect -49173 -29862 -49165 -29238
rect -49485 -29890 -49165 -29862
rect 8615 -29238 8935 -29210
rect 8615 -29862 8623 -29238
rect 8927 -29862 8935 -29238
rect 8615 -29890 8935 -29862
rect 9615 -29238 9935 -29210
rect 9615 -29862 9623 -29238
rect 9927 -29862 9935 -29238
rect 9615 -29890 9935 -29862
rect 10615 -29238 10935 -29210
rect 10615 -29862 10623 -29238
rect 10927 -29862 10935 -29238
rect 10615 -29890 10935 -29862
rect 11615 -29238 11935 -29210
rect 11615 -29862 11623 -29238
rect 11927 -29862 11935 -29238
rect 11615 -29890 11935 -29862
rect 12615 -29238 12935 -29210
rect 12615 -29862 12623 -29238
rect 12927 -29862 12935 -29238
rect 12615 -29890 12935 -29862
rect 13615 -29238 13935 -29210
rect 13615 -29862 13623 -29238
rect 13927 -29862 13935 -29238
rect 13615 -29890 13935 -29862
rect 14615 -29238 14935 -29210
rect 14615 -29862 14623 -29238
rect 14927 -29862 14935 -29238
rect 14615 -29890 14935 -29862
rect 15615 -29238 15935 -29210
rect 15615 -29862 15623 -29238
rect 15927 -29862 15935 -29238
rect 15615 -29890 15935 -29862
rect 16615 -29238 16935 -29210
rect 16615 -29862 16623 -29238
rect 16927 -29862 16935 -29238
rect 16615 -29890 16935 -29862
rect 17615 -29238 17935 -29210
rect 17615 -29862 17623 -29238
rect 17927 -29862 17935 -29238
rect 17615 -29890 17935 -29862
rect 18615 -29238 18935 -29210
rect 18615 -29862 18623 -29238
rect 18927 -29862 18935 -29238
rect 18615 -29890 18935 -29862
rect 19615 -29238 19935 -29210
rect 19615 -29862 19623 -29238
rect 19927 -29862 19935 -29238
rect 19615 -29890 19935 -29862
rect 20615 -29238 20935 -29210
rect 20615 -29862 20623 -29238
rect 20927 -29862 20935 -29238
rect 20615 -29890 20935 -29862
rect 21615 -29238 21935 -29210
rect 21615 -29862 21623 -29238
rect 21927 -29862 21935 -29238
rect 21615 -29890 21935 -29862
rect 22615 -29238 22935 -29210
rect 22615 -29862 22623 -29238
rect 22927 -29862 22935 -29238
rect 22615 -29890 22935 -29862
rect 23615 -29238 23935 -29210
rect 23615 -29862 23623 -29238
rect 23927 -29862 23935 -29238
rect 23615 -29890 23935 -29862
rect 24615 -29238 24935 -29210
rect 24615 -29862 24623 -29238
rect 24927 -29862 24935 -29238
rect 24615 -29890 24935 -29862
rect 25615 -29238 25935 -29210
rect 25615 -29862 25623 -29238
rect 25927 -29862 25935 -29238
rect 25615 -29890 25935 -29862
rect 26615 -29238 26935 -29210
rect 26615 -29862 26623 -29238
rect 26927 -29862 26935 -29238
rect 26615 -29890 26935 -29862
rect 27615 -29238 27935 -29210
rect 27615 -29862 27623 -29238
rect 27927 -29862 27935 -29238
rect 27615 -29890 27935 -29862
rect 28615 -29238 28935 -29210
rect 28615 -29862 28623 -29238
rect 28927 -29862 28935 -29238
rect 28615 -29890 28935 -29862
rect 29615 -29238 29935 -29210
rect 29615 -29862 29623 -29238
rect 29927 -29862 29935 -29238
rect 29615 -29890 29935 -29862
rect 30615 -29238 30935 -29210
rect 30615 -29862 30623 -29238
rect 30927 -29862 30935 -29238
rect 30615 -29890 30935 -29862
rect 31615 -29238 31935 -29210
rect 31615 -29862 31623 -29238
rect 31927 -29862 31935 -29238
rect 31615 -29890 31935 -29862
rect 32615 -29238 32935 -29210
rect 32615 -29862 32623 -29238
rect 32927 -29862 32935 -29238
rect 32615 -29890 32935 -29862
rect 33615 -29238 33935 -29210
rect 33615 -29862 33623 -29238
rect 33927 -29862 33935 -29238
rect 33615 -29890 33935 -29862
rect -74825 -29898 -48825 -29890
rect -74825 -30202 -74817 -29898
rect -74513 -30202 -74477 -29898
rect -74173 -30202 -74137 -29898
rect -73513 -30202 -73477 -29898
rect -73173 -30202 -73137 -29898
rect -72513 -30202 -72477 -29898
rect -72173 -30202 -72137 -29898
rect -71513 -30202 -71477 -29898
rect -71173 -30202 -71137 -29898
rect -70513 -30202 -70477 -29898
rect -70173 -30202 -70137 -29898
rect -69513 -30202 -69477 -29898
rect -69173 -30202 -69137 -29898
rect -68513 -30202 -68477 -29898
rect -68173 -30202 -68137 -29898
rect -67513 -30202 -67477 -29898
rect -67173 -30202 -67137 -29898
rect -66513 -30202 -66477 -29898
rect -66173 -30202 -66137 -29898
rect -65513 -30202 -65477 -29898
rect -65173 -30202 -65137 -29898
rect -64513 -30202 -64477 -29898
rect -64173 -30202 -64137 -29898
rect -63513 -30202 -63477 -29898
rect -63173 -30202 -63137 -29898
rect -62513 -30202 -62477 -29898
rect -62173 -30202 -62137 -29898
rect -61513 -30202 -61477 -29898
rect -61173 -30202 -61137 -29898
rect -60513 -30202 -60477 -29898
rect -60173 -30202 -60137 -29898
rect -59513 -30202 -59477 -29898
rect -59173 -30202 -59137 -29898
rect -58513 -30202 -58477 -29898
rect -58173 -30202 -58137 -29898
rect -57513 -30202 -57477 -29898
rect -57173 -30202 -57137 -29898
rect -56513 -30202 -56477 -29898
rect -56173 -30202 -56137 -29898
rect -55513 -30202 -55477 -29898
rect -55173 -30202 -55137 -29898
rect -54513 -30202 -54477 -29898
rect -54173 -30202 -54137 -29898
rect -53513 -30202 -53477 -29898
rect -53173 -30202 -53137 -29898
rect -52513 -30202 -52477 -29898
rect -52173 -30202 -52137 -29898
rect -51513 -30202 -51477 -29898
rect -51173 -30202 -51137 -29898
rect -50513 -30202 -50477 -29898
rect -50173 -30202 -50137 -29898
rect -49513 -30202 -49477 -29898
rect -49173 -30202 -49137 -29898
rect -48833 -30202 -48825 -29898
rect -74825 -30210 -48825 -30202
rect 8275 -29898 34275 -29890
rect 8275 -30202 8283 -29898
rect 8587 -30202 8623 -29898
rect 8927 -30202 8963 -29898
rect 9587 -30202 9623 -29898
rect 9927 -30202 9963 -29898
rect 10587 -30202 10623 -29898
rect 10927 -30202 10963 -29898
rect 11587 -30202 11623 -29898
rect 11927 -30202 11963 -29898
rect 12587 -30202 12623 -29898
rect 12927 -30202 12963 -29898
rect 13587 -30202 13623 -29898
rect 13927 -30202 13963 -29898
rect 14587 -30202 14623 -29898
rect 14927 -30202 14963 -29898
rect 15587 -30202 15623 -29898
rect 15927 -30202 15963 -29898
rect 16587 -30202 16623 -29898
rect 16927 -30202 16963 -29898
rect 17587 -30202 17623 -29898
rect 17927 -30202 17963 -29898
rect 18587 -30202 18623 -29898
rect 18927 -30202 18963 -29898
rect 19587 -30202 19623 -29898
rect 19927 -30202 19963 -29898
rect 20587 -30202 20623 -29898
rect 20927 -30202 20963 -29898
rect 21587 -30202 21623 -29898
rect 21927 -30202 21963 -29898
rect 22587 -30202 22623 -29898
rect 22927 -30202 22963 -29898
rect 23587 -30202 23623 -29898
rect 23927 -30202 23963 -29898
rect 24587 -30202 24623 -29898
rect 24927 -30202 24963 -29898
rect 25587 -30202 25623 -29898
rect 25927 -30202 25963 -29898
rect 26587 -30202 26623 -29898
rect 26927 -30202 26963 -29898
rect 27587 -30202 27623 -29898
rect 27927 -30202 27963 -29898
rect 28587 -30202 28623 -29898
rect 28927 -30202 28963 -29898
rect 29587 -30202 29623 -29898
rect 29927 -30202 29963 -29898
rect 30587 -30202 30623 -29898
rect 30927 -30202 30963 -29898
rect 31587 -30202 31623 -29898
rect 31927 -30202 31963 -29898
rect 32587 -30202 32623 -29898
rect 32927 -30202 32963 -29898
rect 33587 -30202 33623 -29898
rect 33927 -30202 33963 -29898
rect 34267 -30202 34275 -29898
rect 8275 -30210 34275 -30202
rect -74485 -30238 -74165 -30210
rect -74485 -30862 -74477 -30238
rect -74173 -30862 -74165 -30238
rect -74485 -30890 -74165 -30862
rect -73485 -30238 -73165 -30210
rect -73485 -30862 -73477 -30238
rect -73173 -30862 -73165 -30238
rect -73485 -30890 -73165 -30862
rect -72485 -30238 -72165 -30210
rect -72485 -30862 -72477 -30238
rect -72173 -30862 -72165 -30238
rect -72485 -30890 -72165 -30862
rect -71485 -30238 -71165 -30210
rect -71485 -30862 -71477 -30238
rect -71173 -30862 -71165 -30238
rect -71485 -30890 -71165 -30862
rect -70485 -30238 -70165 -30210
rect -70485 -30862 -70477 -30238
rect -70173 -30862 -70165 -30238
rect -70485 -30890 -70165 -30862
rect -69485 -30238 -69165 -30210
rect -69485 -30862 -69477 -30238
rect -69173 -30862 -69165 -30238
rect -69485 -30890 -69165 -30862
rect -68485 -30238 -68165 -30210
rect -68485 -30862 -68477 -30238
rect -68173 -30862 -68165 -30238
rect -68485 -30890 -68165 -30862
rect -67485 -30238 -67165 -30210
rect -67485 -30862 -67477 -30238
rect -67173 -30862 -67165 -30238
rect -67485 -30890 -67165 -30862
rect -66485 -30238 -66165 -30210
rect -66485 -30862 -66477 -30238
rect -66173 -30862 -66165 -30238
rect -66485 -30890 -66165 -30862
rect -65485 -30238 -65165 -30210
rect -65485 -30862 -65477 -30238
rect -65173 -30862 -65165 -30238
rect -65485 -30890 -65165 -30862
rect -64485 -30238 -64165 -30210
rect -64485 -30862 -64477 -30238
rect -64173 -30862 -64165 -30238
rect -64485 -30890 -64165 -30862
rect -63485 -30238 -63165 -30210
rect -63485 -30862 -63477 -30238
rect -63173 -30862 -63165 -30238
rect -63485 -30890 -63165 -30862
rect -62485 -30238 -62165 -30210
rect -62485 -30862 -62477 -30238
rect -62173 -30862 -62165 -30238
rect -62485 -30890 -62165 -30862
rect -61485 -30238 -61165 -30210
rect -61485 -30862 -61477 -30238
rect -61173 -30862 -61165 -30238
rect -61485 -30890 -61165 -30862
rect -60485 -30238 -60165 -30210
rect -60485 -30862 -60477 -30238
rect -60173 -30862 -60165 -30238
rect -60485 -30890 -60165 -30862
rect -59485 -30238 -59165 -30210
rect -59485 -30862 -59477 -30238
rect -59173 -30862 -59165 -30238
rect -59485 -30890 -59165 -30862
rect -58485 -30238 -58165 -30210
rect -58485 -30862 -58477 -30238
rect -58173 -30862 -58165 -30238
rect -58485 -30890 -58165 -30862
rect -57485 -30238 -57165 -30210
rect -57485 -30862 -57477 -30238
rect -57173 -30862 -57165 -30238
rect -57485 -30890 -57165 -30862
rect -56485 -30238 -56165 -30210
rect -56485 -30862 -56477 -30238
rect -56173 -30862 -56165 -30238
rect -56485 -30890 -56165 -30862
rect -55485 -30238 -55165 -30210
rect -55485 -30862 -55477 -30238
rect -55173 -30862 -55165 -30238
rect -55485 -30890 -55165 -30862
rect -54485 -30238 -54165 -30210
rect -54485 -30862 -54477 -30238
rect -54173 -30862 -54165 -30238
rect -54485 -30890 -54165 -30862
rect -53485 -30238 -53165 -30210
rect -53485 -30862 -53477 -30238
rect -53173 -30862 -53165 -30238
rect -53485 -30890 -53165 -30862
rect -52485 -30238 -52165 -30210
rect -52485 -30862 -52477 -30238
rect -52173 -30862 -52165 -30238
rect -52485 -30890 -52165 -30862
rect -51485 -30238 -51165 -30210
rect -51485 -30862 -51477 -30238
rect -51173 -30862 -51165 -30238
rect -51485 -30890 -51165 -30862
rect -50485 -30238 -50165 -30210
rect -50485 -30862 -50477 -30238
rect -50173 -30862 -50165 -30238
rect -50485 -30890 -50165 -30862
rect -49485 -30238 -49165 -30210
rect -49485 -30862 -49477 -30238
rect -49173 -30862 -49165 -30238
rect -49485 -30890 -49165 -30862
rect 8615 -30238 8935 -30210
rect 8615 -30862 8623 -30238
rect 8927 -30862 8935 -30238
rect 8615 -30890 8935 -30862
rect 9615 -30238 9935 -30210
rect 9615 -30862 9623 -30238
rect 9927 -30862 9935 -30238
rect 9615 -30890 9935 -30862
rect 10615 -30238 10935 -30210
rect 10615 -30862 10623 -30238
rect 10927 -30862 10935 -30238
rect 10615 -30890 10935 -30862
rect 11615 -30238 11935 -30210
rect 11615 -30862 11623 -30238
rect 11927 -30862 11935 -30238
rect 11615 -30890 11935 -30862
rect 12615 -30238 12935 -30210
rect 12615 -30862 12623 -30238
rect 12927 -30862 12935 -30238
rect 12615 -30890 12935 -30862
rect 13615 -30238 13935 -30210
rect 13615 -30862 13623 -30238
rect 13927 -30862 13935 -30238
rect 13615 -30890 13935 -30862
rect 14615 -30238 14935 -30210
rect 14615 -30862 14623 -30238
rect 14927 -30862 14935 -30238
rect 14615 -30890 14935 -30862
rect 15615 -30238 15935 -30210
rect 15615 -30862 15623 -30238
rect 15927 -30862 15935 -30238
rect 15615 -30890 15935 -30862
rect 16615 -30238 16935 -30210
rect 16615 -30862 16623 -30238
rect 16927 -30862 16935 -30238
rect 16615 -30890 16935 -30862
rect 17615 -30238 17935 -30210
rect 17615 -30862 17623 -30238
rect 17927 -30862 17935 -30238
rect 17615 -30890 17935 -30862
rect 18615 -30238 18935 -30210
rect 18615 -30862 18623 -30238
rect 18927 -30862 18935 -30238
rect 18615 -30890 18935 -30862
rect 19615 -30238 19935 -30210
rect 19615 -30862 19623 -30238
rect 19927 -30862 19935 -30238
rect 19615 -30890 19935 -30862
rect 20615 -30238 20935 -30210
rect 20615 -30862 20623 -30238
rect 20927 -30862 20935 -30238
rect 20615 -30890 20935 -30862
rect 21615 -30238 21935 -30210
rect 21615 -30862 21623 -30238
rect 21927 -30862 21935 -30238
rect 21615 -30890 21935 -30862
rect 22615 -30238 22935 -30210
rect 22615 -30862 22623 -30238
rect 22927 -30862 22935 -30238
rect 22615 -30890 22935 -30862
rect 23615 -30238 23935 -30210
rect 23615 -30862 23623 -30238
rect 23927 -30862 23935 -30238
rect 23615 -30890 23935 -30862
rect 24615 -30238 24935 -30210
rect 24615 -30862 24623 -30238
rect 24927 -30862 24935 -30238
rect 24615 -30890 24935 -30862
rect 25615 -30238 25935 -30210
rect 25615 -30862 25623 -30238
rect 25927 -30862 25935 -30238
rect 25615 -30890 25935 -30862
rect 26615 -30238 26935 -30210
rect 26615 -30862 26623 -30238
rect 26927 -30862 26935 -30238
rect 26615 -30890 26935 -30862
rect 27615 -30238 27935 -30210
rect 27615 -30862 27623 -30238
rect 27927 -30862 27935 -30238
rect 27615 -30890 27935 -30862
rect 28615 -30238 28935 -30210
rect 28615 -30862 28623 -30238
rect 28927 -30862 28935 -30238
rect 28615 -30890 28935 -30862
rect 29615 -30238 29935 -30210
rect 29615 -30862 29623 -30238
rect 29927 -30862 29935 -30238
rect 29615 -30890 29935 -30862
rect 30615 -30238 30935 -30210
rect 30615 -30862 30623 -30238
rect 30927 -30862 30935 -30238
rect 30615 -30890 30935 -30862
rect 31615 -30238 31935 -30210
rect 31615 -30862 31623 -30238
rect 31927 -30862 31935 -30238
rect 31615 -30890 31935 -30862
rect 32615 -30238 32935 -30210
rect 32615 -30862 32623 -30238
rect 32927 -30862 32935 -30238
rect 32615 -30890 32935 -30862
rect 33615 -30238 33935 -30210
rect 33615 -30862 33623 -30238
rect 33927 -30862 33935 -30238
rect 33615 -30890 33935 -30862
rect -74825 -30898 -48825 -30890
rect -74825 -31202 -74817 -30898
rect -74513 -31202 -74477 -30898
rect -74173 -31202 -74137 -30898
rect -73513 -31202 -73477 -30898
rect -73173 -31202 -73137 -30898
rect -72513 -31202 -72477 -30898
rect -72173 -31202 -72137 -30898
rect -71513 -31202 -71477 -30898
rect -71173 -31202 -71137 -30898
rect -70513 -31202 -70477 -30898
rect -70173 -31202 -70137 -30898
rect -69513 -31202 -69477 -30898
rect -69173 -31202 -69137 -30898
rect -68513 -31202 -68477 -30898
rect -68173 -31202 -68137 -30898
rect -67513 -31202 -67477 -30898
rect -67173 -31202 -67137 -30898
rect -66513 -31202 -66477 -30898
rect -66173 -31202 -66137 -30898
rect -65513 -31202 -65477 -30898
rect -65173 -31202 -65137 -30898
rect -64513 -31202 -64477 -30898
rect -64173 -31202 -64137 -30898
rect -63513 -31202 -63477 -30898
rect -63173 -31202 -63137 -30898
rect -62513 -31202 -62477 -30898
rect -62173 -31202 -62137 -30898
rect -61513 -31202 -61477 -30898
rect -61173 -31202 -61137 -30898
rect -60513 -31202 -60477 -30898
rect -60173 -31202 -60137 -30898
rect -59513 -31202 -59477 -30898
rect -59173 -31202 -59137 -30898
rect -58513 -31202 -58477 -30898
rect -58173 -31202 -58137 -30898
rect -57513 -31202 -57477 -30898
rect -57173 -31202 -57137 -30898
rect -56513 -31202 -56477 -30898
rect -56173 -31202 -56137 -30898
rect -55513 -31202 -55477 -30898
rect -55173 -31202 -55137 -30898
rect -54513 -31202 -54477 -30898
rect -54173 -31202 -54137 -30898
rect -53513 -31202 -53477 -30898
rect -53173 -31202 -53137 -30898
rect -52513 -31202 -52477 -30898
rect -52173 -31202 -52137 -30898
rect -51513 -31202 -51477 -30898
rect -51173 -31202 -51137 -30898
rect -50513 -31202 -50477 -30898
rect -50173 -31202 -50137 -30898
rect -49513 -31202 -49477 -30898
rect -49173 -31202 -49137 -30898
rect -48833 -31202 -48825 -30898
rect -74825 -31210 -48825 -31202
rect 8275 -30898 34275 -30890
rect 8275 -31202 8283 -30898
rect 8587 -31202 8623 -30898
rect 8927 -31202 8963 -30898
rect 9587 -31202 9623 -30898
rect 9927 -31202 9963 -30898
rect 10587 -31202 10623 -30898
rect 10927 -31202 10963 -30898
rect 11587 -31202 11623 -30898
rect 11927 -31202 11963 -30898
rect 12587 -31202 12623 -30898
rect 12927 -31202 12963 -30898
rect 13587 -31202 13623 -30898
rect 13927 -31202 13963 -30898
rect 14587 -31202 14623 -30898
rect 14927 -31202 14963 -30898
rect 15587 -31202 15623 -30898
rect 15927 -31202 15963 -30898
rect 16587 -31202 16623 -30898
rect 16927 -31202 16963 -30898
rect 17587 -31202 17623 -30898
rect 17927 -31202 17963 -30898
rect 18587 -31202 18623 -30898
rect 18927 -31202 18963 -30898
rect 19587 -31202 19623 -30898
rect 19927 -31202 19963 -30898
rect 20587 -31202 20623 -30898
rect 20927 -31202 20963 -30898
rect 21587 -31202 21623 -30898
rect 21927 -31202 21963 -30898
rect 22587 -31202 22623 -30898
rect 22927 -31202 22963 -30898
rect 23587 -31202 23623 -30898
rect 23927 -31202 23963 -30898
rect 24587 -31202 24623 -30898
rect 24927 -31202 24963 -30898
rect 25587 -31202 25623 -30898
rect 25927 -31202 25963 -30898
rect 26587 -31202 26623 -30898
rect 26927 -31202 26963 -30898
rect 27587 -31202 27623 -30898
rect 27927 -31202 27963 -30898
rect 28587 -31202 28623 -30898
rect 28927 -31202 28963 -30898
rect 29587 -31202 29623 -30898
rect 29927 -31202 29963 -30898
rect 30587 -31202 30623 -30898
rect 30927 -31202 30963 -30898
rect 31587 -31202 31623 -30898
rect 31927 -31202 31963 -30898
rect 32587 -31202 32623 -30898
rect 32927 -31202 32963 -30898
rect 33587 -31202 33623 -30898
rect 33927 -31202 33963 -30898
rect 34267 -31202 34275 -30898
rect 8275 -31210 34275 -31202
rect -74485 -31238 -74165 -31210
rect -74485 -31862 -74477 -31238
rect -74173 -31862 -74165 -31238
rect -74485 -31890 -74165 -31862
rect -73485 -31238 -73165 -31210
rect -73485 -31862 -73477 -31238
rect -73173 -31862 -73165 -31238
rect -73485 -31890 -73165 -31862
rect -72485 -31238 -72165 -31210
rect -72485 -31862 -72477 -31238
rect -72173 -31862 -72165 -31238
rect -72485 -31890 -72165 -31862
rect -71485 -31238 -71165 -31210
rect -71485 -31862 -71477 -31238
rect -71173 -31862 -71165 -31238
rect -71485 -31890 -71165 -31862
rect -70485 -31238 -70165 -31210
rect -70485 -31862 -70477 -31238
rect -70173 -31862 -70165 -31238
rect -70485 -31890 -70165 -31862
rect -69485 -31238 -69165 -31210
rect -69485 -31862 -69477 -31238
rect -69173 -31862 -69165 -31238
rect -69485 -31890 -69165 -31862
rect -68485 -31238 -68165 -31210
rect -68485 -31862 -68477 -31238
rect -68173 -31862 -68165 -31238
rect -68485 -31890 -68165 -31862
rect -67485 -31238 -67165 -31210
rect -67485 -31862 -67477 -31238
rect -67173 -31862 -67165 -31238
rect -67485 -31890 -67165 -31862
rect -66485 -31238 -66165 -31210
rect -66485 -31862 -66477 -31238
rect -66173 -31862 -66165 -31238
rect -66485 -31890 -66165 -31862
rect -65485 -31238 -65165 -31210
rect -65485 -31862 -65477 -31238
rect -65173 -31862 -65165 -31238
rect -65485 -31890 -65165 -31862
rect -64485 -31238 -64165 -31210
rect -64485 -31862 -64477 -31238
rect -64173 -31862 -64165 -31238
rect -64485 -31890 -64165 -31862
rect -63485 -31238 -63165 -31210
rect -63485 -31862 -63477 -31238
rect -63173 -31862 -63165 -31238
rect -63485 -31890 -63165 -31862
rect -62485 -31238 -62165 -31210
rect -62485 -31862 -62477 -31238
rect -62173 -31862 -62165 -31238
rect -62485 -31890 -62165 -31862
rect -61485 -31238 -61165 -31210
rect -61485 -31862 -61477 -31238
rect -61173 -31862 -61165 -31238
rect -61485 -31890 -61165 -31862
rect -60485 -31238 -60165 -31210
rect -60485 -31862 -60477 -31238
rect -60173 -31862 -60165 -31238
rect -60485 -31890 -60165 -31862
rect -59485 -31238 -59165 -31210
rect -59485 -31862 -59477 -31238
rect -59173 -31862 -59165 -31238
rect -59485 -31890 -59165 -31862
rect -58485 -31238 -58165 -31210
rect -58485 -31862 -58477 -31238
rect -58173 -31862 -58165 -31238
rect -58485 -31890 -58165 -31862
rect -57485 -31238 -57165 -31210
rect -57485 -31862 -57477 -31238
rect -57173 -31862 -57165 -31238
rect -57485 -31890 -57165 -31862
rect -56485 -31238 -56165 -31210
rect -56485 -31862 -56477 -31238
rect -56173 -31862 -56165 -31238
rect -56485 -31890 -56165 -31862
rect -55485 -31238 -55165 -31210
rect -55485 -31862 -55477 -31238
rect -55173 -31862 -55165 -31238
rect -55485 -31890 -55165 -31862
rect -54485 -31238 -54165 -31210
rect -54485 -31862 -54477 -31238
rect -54173 -31862 -54165 -31238
rect -54485 -31890 -54165 -31862
rect -53485 -31238 -53165 -31210
rect -53485 -31862 -53477 -31238
rect -53173 -31862 -53165 -31238
rect -53485 -31890 -53165 -31862
rect -52485 -31238 -52165 -31210
rect -52485 -31862 -52477 -31238
rect -52173 -31862 -52165 -31238
rect -52485 -31890 -52165 -31862
rect -51485 -31238 -51165 -31210
rect -51485 -31862 -51477 -31238
rect -51173 -31862 -51165 -31238
rect -51485 -31890 -51165 -31862
rect -50485 -31238 -50165 -31210
rect -50485 -31862 -50477 -31238
rect -50173 -31862 -50165 -31238
rect -50485 -31890 -50165 -31862
rect -49485 -31238 -49165 -31210
rect -49485 -31862 -49477 -31238
rect -49173 -31862 -49165 -31238
rect -49485 -31890 -49165 -31862
rect 8615 -31238 8935 -31210
rect 8615 -31862 8623 -31238
rect 8927 -31862 8935 -31238
rect 8615 -31890 8935 -31862
rect 9615 -31238 9935 -31210
rect 9615 -31862 9623 -31238
rect 9927 -31862 9935 -31238
rect 9615 -31890 9935 -31862
rect 10615 -31238 10935 -31210
rect 10615 -31862 10623 -31238
rect 10927 -31862 10935 -31238
rect 10615 -31890 10935 -31862
rect 11615 -31238 11935 -31210
rect 11615 -31862 11623 -31238
rect 11927 -31862 11935 -31238
rect 11615 -31890 11935 -31862
rect 12615 -31238 12935 -31210
rect 12615 -31862 12623 -31238
rect 12927 -31862 12935 -31238
rect 12615 -31890 12935 -31862
rect 13615 -31238 13935 -31210
rect 13615 -31862 13623 -31238
rect 13927 -31862 13935 -31238
rect 13615 -31890 13935 -31862
rect 14615 -31238 14935 -31210
rect 14615 -31862 14623 -31238
rect 14927 -31862 14935 -31238
rect 14615 -31890 14935 -31862
rect 15615 -31238 15935 -31210
rect 15615 -31862 15623 -31238
rect 15927 -31862 15935 -31238
rect 15615 -31890 15935 -31862
rect 16615 -31238 16935 -31210
rect 16615 -31862 16623 -31238
rect 16927 -31862 16935 -31238
rect 16615 -31890 16935 -31862
rect 17615 -31238 17935 -31210
rect 17615 -31862 17623 -31238
rect 17927 -31862 17935 -31238
rect 17615 -31890 17935 -31862
rect 18615 -31238 18935 -31210
rect 18615 -31862 18623 -31238
rect 18927 -31862 18935 -31238
rect 18615 -31890 18935 -31862
rect 19615 -31238 19935 -31210
rect 19615 -31862 19623 -31238
rect 19927 -31862 19935 -31238
rect 19615 -31890 19935 -31862
rect 20615 -31238 20935 -31210
rect 20615 -31862 20623 -31238
rect 20927 -31862 20935 -31238
rect 20615 -31890 20935 -31862
rect 21615 -31238 21935 -31210
rect 21615 -31862 21623 -31238
rect 21927 -31862 21935 -31238
rect 21615 -31890 21935 -31862
rect 22615 -31238 22935 -31210
rect 22615 -31862 22623 -31238
rect 22927 -31862 22935 -31238
rect 22615 -31890 22935 -31862
rect 23615 -31238 23935 -31210
rect 23615 -31862 23623 -31238
rect 23927 -31862 23935 -31238
rect 23615 -31890 23935 -31862
rect 24615 -31238 24935 -31210
rect 24615 -31862 24623 -31238
rect 24927 -31862 24935 -31238
rect 24615 -31890 24935 -31862
rect 25615 -31238 25935 -31210
rect 25615 -31862 25623 -31238
rect 25927 -31862 25935 -31238
rect 25615 -31890 25935 -31862
rect 26615 -31238 26935 -31210
rect 26615 -31862 26623 -31238
rect 26927 -31862 26935 -31238
rect 26615 -31890 26935 -31862
rect 27615 -31238 27935 -31210
rect 27615 -31862 27623 -31238
rect 27927 -31862 27935 -31238
rect 27615 -31890 27935 -31862
rect 28615 -31238 28935 -31210
rect 28615 -31862 28623 -31238
rect 28927 -31862 28935 -31238
rect 28615 -31890 28935 -31862
rect 29615 -31238 29935 -31210
rect 29615 -31862 29623 -31238
rect 29927 -31862 29935 -31238
rect 29615 -31890 29935 -31862
rect 30615 -31238 30935 -31210
rect 30615 -31862 30623 -31238
rect 30927 -31862 30935 -31238
rect 30615 -31890 30935 -31862
rect 31615 -31238 31935 -31210
rect 31615 -31862 31623 -31238
rect 31927 -31862 31935 -31238
rect 31615 -31890 31935 -31862
rect 32615 -31238 32935 -31210
rect 32615 -31862 32623 -31238
rect 32927 -31862 32935 -31238
rect 32615 -31890 32935 -31862
rect 33615 -31238 33935 -31210
rect 33615 -31862 33623 -31238
rect 33927 -31862 33935 -31238
rect 33615 -31890 33935 -31862
rect -74825 -31898 -48825 -31890
rect -74825 -32202 -74817 -31898
rect -74513 -32202 -74477 -31898
rect -74173 -32202 -74137 -31898
rect -73513 -32202 -73477 -31898
rect -73173 -32202 -73137 -31898
rect -72513 -32202 -72477 -31898
rect -72173 -32202 -72137 -31898
rect -71513 -32202 -71477 -31898
rect -71173 -32202 -71137 -31898
rect -70513 -32202 -70477 -31898
rect -70173 -32202 -70137 -31898
rect -69513 -32202 -69477 -31898
rect -69173 -32202 -69137 -31898
rect -68513 -32202 -68477 -31898
rect -68173 -32202 -68137 -31898
rect -67513 -32202 -67477 -31898
rect -67173 -32202 -67137 -31898
rect -66513 -32202 -66477 -31898
rect -66173 -32202 -66137 -31898
rect -65513 -32202 -65477 -31898
rect -65173 -32202 -65137 -31898
rect -64513 -32202 -64477 -31898
rect -64173 -32202 -64137 -31898
rect -63513 -32202 -63477 -31898
rect -63173 -32202 -63137 -31898
rect -62513 -32202 -62477 -31898
rect -62173 -32202 -62137 -31898
rect -61513 -32202 -61477 -31898
rect -61173 -32202 -61137 -31898
rect -60513 -32202 -60477 -31898
rect -60173 -32202 -60137 -31898
rect -59513 -32202 -59477 -31898
rect -59173 -32202 -59137 -31898
rect -58513 -32202 -58477 -31898
rect -58173 -32202 -58137 -31898
rect -57513 -32202 -57477 -31898
rect -57173 -32202 -57137 -31898
rect -56513 -32202 -56477 -31898
rect -56173 -32202 -56137 -31898
rect -55513 -32202 -55477 -31898
rect -55173 -32202 -55137 -31898
rect -54513 -32202 -54477 -31898
rect -54173 -32202 -54137 -31898
rect -53513 -32202 -53477 -31898
rect -53173 -32202 -53137 -31898
rect -52513 -32202 -52477 -31898
rect -52173 -32202 -52137 -31898
rect -51513 -32202 -51477 -31898
rect -51173 -32202 -51137 -31898
rect -50513 -32202 -50477 -31898
rect -50173 -32202 -50137 -31898
rect -49513 -32202 -49477 -31898
rect -49173 -32202 -49137 -31898
rect -48833 -32202 -48825 -31898
rect -74825 -32210 -48825 -32202
rect 8275 -31898 34275 -31890
rect 8275 -32202 8283 -31898
rect 8587 -32202 8623 -31898
rect 8927 -32202 8963 -31898
rect 9587 -32202 9623 -31898
rect 9927 -32202 9963 -31898
rect 10587 -32202 10623 -31898
rect 10927 -32202 10963 -31898
rect 11587 -32202 11623 -31898
rect 11927 -32202 11963 -31898
rect 12587 -32202 12623 -31898
rect 12927 -32202 12963 -31898
rect 13587 -32202 13623 -31898
rect 13927 -32202 13963 -31898
rect 14587 -32202 14623 -31898
rect 14927 -32202 14963 -31898
rect 15587 -32202 15623 -31898
rect 15927 -32202 15963 -31898
rect 16587 -32202 16623 -31898
rect 16927 -32202 16963 -31898
rect 17587 -32202 17623 -31898
rect 17927 -32202 17963 -31898
rect 18587 -32202 18623 -31898
rect 18927 -32202 18963 -31898
rect 19587 -32202 19623 -31898
rect 19927 -32202 19963 -31898
rect 20587 -32202 20623 -31898
rect 20927 -32202 20963 -31898
rect 21587 -32202 21623 -31898
rect 21927 -32202 21963 -31898
rect 22587 -32202 22623 -31898
rect 22927 -32202 22963 -31898
rect 23587 -32202 23623 -31898
rect 23927 -32202 23963 -31898
rect 24587 -32202 24623 -31898
rect 24927 -32202 24963 -31898
rect 25587 -32202 25623 -31898
rect 25927 -32202 25963 -31898
rect 26587 -32202 26623 -31898
rect 26927 -32202 26963 -31898
rect 27587 -32202 27623 -31898
rect 27927 -32202 27963 -31898
rect 28587 -32202 28623 -31898
rect 28927 -32202 28963 -31898
rect 29587 -32202 29623 -31898
rect 29927 -32202 29963 -31898
rect 30587 -32202 30623 -31898
rect 30927 -32202 30963 -31898
rect 31587 -32202 31623 -31898
rect 31927 -32202 31963 -31898
rect 32587 -32202 32623 -31898
rect 32927 -32202 32963 -31898
rect 33587 -32202 33623 -31898
rect 33927 -32202 33963 -31898
rect 34267 -32202 34275 -31898
rect 8275 -32210 34275 -32202
rect -74485 -32238 -74165 -32210
rect -74485 -32862 -74477 -32238
rect -74173 -32862 -74165 -32238
rect -74485 -32890 -74165 -32862
rect -73485 -32238 -73165 -32210
rect -73485 -32862 -73477 -32238
rect -73173 -32862 -73165 -32238
rect -73485 -32890 -73165 -32862
rect -72485 -32238 -72165 -32210
rect -72485 -32862 -72477 -32238
rect -72173 -32862 -72165 -32238
rect -72485 -32890 -72165 -32862
rect -71485 -32238 -71165 -32210
rect -71485 -32862 -71477 -32238
rect -71173 -32862 -71165 -32238
rect -71485 -32890 -71165 -32862
rect -70485 -32238 -70165 -32210
rect -70485 -32862 -70477 -32238
rect -70173 -32862 -70165 -32238
rect -70485 -32890 -70165 -32862
rect -69485 -32238 -69165 -32210
rect -69485 -32862 -69477 -32238
rect -69173 -32862 -69165 -32238
rect -69485 -32890 -69165 -32862
rect -68485 -32238 -68165 -32210
rect -68485 -32862 -68477 -32238
rect -68173 -32862 -68165 -32238
rect -68485 -32890 -68165 -32862
rect -67485 -32238 -67165 -32210
rect -67485 -32862 -67477 -32238
rect -67173 -32862 -67165 -32238
rect -67485 -32890 -67165 -32862
rect -66485 -32238 -66165 -32210
rect -66485 -32862 -66477 -32238
rect -66173 -32862 -66165 -32238
rect -66485 -32890 -66165 -32862
rect -65485 -32238 -65165 -32210
rect -65485 -32862 -65477 -32238
rect -65173 -32862 -65165 -32238
rect -65485 -32890 -65165 -32862
rect -64485 -32238 -64165 -32210
rect -64485 -32862 -64477 -32238
rect -64173 -32862 -64165 -32238
rect -64485 -32890 -64165 -32862
rect -63485 -32238 -63165 -32210
rect -63485 -32862 -63477 -32238
rect -63173 -32862 -63165 -32238
rect -63485 -32890 -63165 -32862
rect -62485 -32238 -62165 -32210
rect -62485 -32862 -62477 -32238
rect -62173 -32862 -62165 -32238
rect -62485 -32890 -62165 -32862
rect -61485 -32238 -61165 -32210
rect -61485 -32862 -61477 -32238
rect -61173 -32862 -61165 -32238
rect -61485 -32890 -61165 -32862
rect -60485 -32238 -60165 -32210
rect -60485 -32862 -60477 -32238
rect -60173 -32862 -60165 -32238
rect -60485 -32890 -60165 -32862
rect -59485 -32238 -59165 -32210
rect -59485 -32862 -59477 -32238
rect -59173 -32862 -59165 -32238
rect -59485 -32890 -59165 -32862
rect -58485 -32238 -58165 -32210
rect -58485 -32862 -58477 -32238
rect -58173 -32862 -58165 -32238
rect -58485 -32890 -58165 -32862
rect -57485 -32238 -57165 -32210
rect -57485 -32862 -57477 -32238
rect -57173 -32862 -57165 -32238
rect -57485 -32890 -57165 -32862
rect -56485 -32238 -56165 -32210
rect -56485 -32862 -56477 -32238
rect -56173 -32862 -56165 -32238
rect -56485 -32890 -56165 -32862
rect -55485 -32238 -55165 -32210
rect -55485 -32862 -55477 -32238
rect -55173 -32862 -55165 -32238
rect -55485 -32890 -55165 -32862
rect -54485 -32238 -54165 -32210
rect -54485 -32862 -54477 -32238
rect -54173 -32862 -54165 -32238
rect -54485 -32890 -54165 -32862
rect -53485 -32238 -53165 -32210
rect -53485 -32862 -53477 -32238
rect -53173 -32862 -53165 -32238
rect -53485 -32890 -53165 -32862
rect -52485 -32238 -52165 -32210
rect -52485 -32862 -52477 -32238
rect -52173 -32862 -52165 -32238
rect -52485 -32890 -52165 -32862
rect -51485 -32238 -51165 -32210
rect -51485 -32862 -51477 -32238
rect -51173 -32862 -51165 -32238
rect -51485 -32890 -51165 -32862
rect -50485 -32238 -50165 -32210
rect -50485 -32862 -50477 -32238
rect -50173 -32862 -50165 -32238
rect -50485 -32890 -50165 -32862
rect -49485 -32238 -49165 -32210
rect -49485 -32862 -49477 -32238
rect -49173 -32862 -49165 -32238
rect 8615 -32238 8935 -32210
rect -49485 -32890 -49165 -32862
rect -46275 -32598 -36275 -32550
rect -74825 -32898 -48825 -32890
rect -74825 -33202 -74817 -32898
rect -74513 -33202 -74477 -32898
rect -74173 -33202 -74137 -32898
rect -73513 -33202 -73477 -32898
rect -73173 -33202 -73137 -32898
rect -72513 -33202 -72477 -32898
rect -72173 -33202 -72137 -32898
rect -71513 -33202 -71477 -32898
rect -71173 -33202 -71137 -32898
rect -70513 -33202 -70477 -32898
rect -70173 -33202 -70137 -32898
rect -69513 -33202 -69477 -32898
rect -69173 -33202 -69137 -32898
rect -68513 -33202 -68477 -32898
rect -68173 -33202 -68137 -32898
rect -67513 -33202 -67477 -32898
rect -67173 -33202 -67137 -32898
rect -66513 -33202 -66477 -32898
rect -66173 -33202 -66137 -32898
rect -65513 -33202 -65477 -32898
rect -65173 -33202 -65137 -32898
rect -64513 -33202 -64477 -32898
rect -64173 -33202 -64137 -32898
rect -63513 -33202 -63477 -32898
rect -63173 -33202 -63137 -32898
rect -62513 -33202 -62477 -32898
rect -62173 -33202 -62137 -32898
rect -61513 -33202 -61477 -32898
rect -61173 -33202 -61137 -32898
rect -60513 -33202 -60477 -32898
rect -60173 -33202 -60137 -32898
rect -59513 -33202 -59477 -32898
rect -59173 -33202 -59137 -32898
rect -58513 -33202 -58477 -32898
rect -58173 -33202 -58137 -32898
rect -57513 -33202 -57477 -32898
rect -57173 -33202 -57137 -32898
rect -56513 -33202 -56477 -32898
rect -56173 -33202 -56137 -32898
rect -55513 -33202 -55477 -32898
rect -55173 -33202 -55137 -32898
rect -54513 -33202 -54477 -32898
rect -54173 -33202 -54137 -32898
rect -53513 -33202 -53477 -32898
rect -53173 -33202 -53137 -32898
rect -52513 -33202 -52477 -32898
rect -52173 -33202 -52137 -32898
rect -51513 -33202 -51477 -32898
rect -51173 -33202 -51137 -32898
rect -50513 -33202 -50477 -32898
rect -50173 -33202 -50137 -32898
rect -49513 -33202 -49477 -32898
rect -49173 -33202 -49137 -32898
rect -48833 -33202 -48825 -32898
rect -74825 -33210 -48825 -33202
rect -74485 -33238 -74165 -33210
rect -74485 -33862 -74477 -33238
rect -74173 -33862 -74165 -33238
rect -74485 -33890 -74165 -33862
rect -73485 -33238 -73165 -33210
rect -73485 -33862 -73477 -33238
rect -73173 -33862 -73165 -33238
rect -73485 -33890 -73165 -33862
rect -72485 -33238 -72165 -33210
rect -72485 -33862 -72477 -33238
rect -72173 -33862 -72165 -33238
rect -72485 -33890 -72165 -33862
rect -71485 -33238 -71165 -33210
rect -71485 -33862 -71477 -33238
rect -71173 -33862 -71165 -33238
rect -71485 -33890 -71165 -33862
rect -70485 -33238 -70165 -33210
rect -70485 -33862 -70477 -33238
rect -70173 -33862 -70165 -33238
rect -70485 -33890 -70165 -33862
rect -69485 -33238 -69165 -33210
rect -69485 -33862 -69477 -33238
rect -69173 -33862 -69165 -33238
rect -69485 -33890 -69165 -33862
rect -68485 -33238 -68165 -33210
rect -68485 -33862 -68477 -33238
rect -68173 -33862 -68165 -33238
rect -68485 -33890 -68165 -33862
rect -67485 -33238 -67165 -33210
rect -67485 -33862 -67477 -33238
rect -67173 -33862 -67165 -33238
rect -67485 -33890 -67165 -33862
rect -66485 -33238 -66165 -33210
rect -66485 -33862 -66477 -33238
rect -66173 -33862 -66165 -33238
rect -66485 -33890 -66165 -33862
rect -65485 -33238 -65165 -33210
rect -65485 -33862 -65477 -33238
rect -65173 -33862 -65165 -33238
rect -65485 -33890 -65165 -33862
rect -64485 -33238 -64165 -33210
rect -64485 -33862 -64477 -33238
rect -64173 -33862 -64165 -33238
rect -64485 -33890 -64165 -33862
rect -63485 -33238 -63165 -33210
rect -63485 -33862 -63477 -33238
rect -63173 -33862 -63165 -33238
rect -63485 -33890 -63165 -33862
rect -62485 -33238 -62165 -33210
rect -62485 -33862 -62477 -33238
rect -62173 -33862 -62165 -33238
rect -62485 -33890 -62165 -33862
rect -61485 -33238 -61165 -33210
rect -61485 -33862 -61477 -33238
rect -61173 -33862 -61165 -33238
rect -61485 -33890 -61165 -33862
rect -60485 -33238 -60165 -33210
rect -60485 -33862 -60477 -33238
rect -60173 -33862 -60165 -33238
rect -60485 -33890 -60165 -33862
rect -59485 -33238 -59165 -33210
rect -59485 -33862 -59477 -33238
rect -59173 -33862 -59165 -33238
rect -59485 -33890 -59165 -33862
rect -58485 -33238 -58165 -33210
rect -58485 -33862 -58477 -33238
rect -58173 -33862 -58165 -33238
rect -58485 -33890 -58165 -33862
rect -57485 -33238 -57165 -33210
rect -57485 -33862 -57477 -33238
rect -57173 -33862 -57165 -33238
rect -57485 -33890 -57165 -33862
rect -56485 -33238 -56165 -33210
rect -56485 -33862 -56477 -33238
rect -56173 -33862 -56165 -33238
rect -56485 -33890 -56165 -33862
rect -55485 -33238 -55165 -33210
rect -55485 -33862 -55477 -33238
rect -55173 -33862 -55165 -33238
rect -55485 -33890 -55165 -33862
rect -54485 -33238 -54165 -33210
rect -54485 -33862 -54477 -33238
rect -54173 -33862 -54165 -33238
rect -54485 -33890 -54165 -33862
rect -53485 -33238 -53165 -33210
rect -53485 -33862 -53477 -33238
rect -53173 -33862 -53165 -33238
rect -53485 -33890 -53165 -33862
rect -52485 -33238 -52165 -33210
rect -52485 -33862 -52477 -33238
rect -52173 -33862 -52165 -33238
rect -52485 -33890 -52165 -33862
rect -51485 -33238 -51165 -33210
rect -51485 -33862 -51477 -33238
rect -51173 -33862 -51165 -33238
rect -51485 -33890 -51165 -33862
rect -50485 -33238 -50165 -33210
rect -50485 -33862 -50477 -33238
rect -50173 -33862 -50165 -33238
rect -50485 -33890 -50165 -33862
rect -49485 -33238 -49165 -33210
rect -49485 -33862 -49477 -33238
rect -49173 -33862 -49165 -33238
rect -49485 -33890 -49165 -33862
rect -74825 -33898 -48825 -33890
rect -74825 -34202 -74817 -33898
rect -74513 -34202 -74477 -33898
rect -74173 -34202 -74137 -33898
rect -73513 -34202 -73477 -33898
rect -73173 -34202 -73137 -33898
rect -72513 -34202 -72477 -33898
rect -72173 -34202 -72137 -33898
rect -71513 -34202 -71477 -33898
rect -71173 -34202 -71137 -33898
rect -70513 -34202 -70477 -33898
rect -70173 -34202 -70137 -33898
rect -69513 -34202 -69477 -33898
rect -69173 -34202 -69137 -33898
rect -68513 -34202 -68477 -33898
rect -68173 -34202 -68137 -33898
rect -67513 -34202 -67477 -33898
rect -67173 -34202 -67137 -33898
rect -66513 -34202 -66477 -33898
rect -66173 -34202 -66137 -33898
rect -65513 -34202 -65477 -33898
rect -65173 -34202 -65137 -33898
rect -64513 -34202 -64477 -33898
rect -64173 -34202 -64137 -33898
rect -63513 -34202 -63477 -33898
rect -63173 -34202 -63137 -33898
rect -62513 -34202 -62477 -33898
rect -62173 -34202 -62137 -33898
rect -61513 -34202 -61477 -33898
rect -61173 -34202 -61137 -33898
rect -60513 -34202 -60477 -33898
rect -60173 -34202 -60137 -33898
rect -59513 -34202 -59477 -33898
rect -59173 -34202 -59137 -33898
rect -58513 -34202 -58477 -33898
rect -58173 -34202 -58137 -33898
rect -57513 -34202 -57477 -33898
rect -57173 -34202 -57137 -33898
rect -56513 -34202 -56477 -33898
rect -56173 -34202 -56137 -33898
rect -55513 -34202 -55477 -33898
rect -55173 -34202 -55137 -33898
rect -54513 -34202 -54477 -33898
rect -54173 -34202 -54137 -33898
rect -53513 -34202 -53477 -33898
rect -53173 -34202 -53137 -33898
rect -52513 -34202 -52477 -33898
rect -52173 -34202 -52137 -33898
rect -51513 -34202 -51477 -33898
rect -51173 -34202 -51137 -33898
rect -50513 -34202 -50477 -33898
rect -50173 -34202 -50137 -33898
rect -49513 -34202 -49477 -33898
rect -49173 -34202 -49137 -33898
rect -48833 -34202 -48825 -33898
rect -74825 -34210 -48825 -34202
rect -74485 -34238 -74165 -34210
rect -74485 -34862 -74477 -34238
rect -74173 -34862 -74165 -34238
rect -74485 -34890 -74165 -34862
rect -73485 -34238 -73165 -34210
rect -73485 -34862 -73477 -34238
rect -73173 -34862 -73165 -34238
rect -73485 -34890 -73165 -34862
rect -72485 -34238 -72165 -34210
rect -72485 -34862 -72477 -34238
rect -72173 -34862 -72165 -34238
rect -72485 -34890 -72165 -34862
rect -71485 -34238 -71165 -34210
rect -71485 -34862 -71477 -34238
rect -71173 -34862 -71165 -34238
rect -71485 -34890 -71165 -34862
rect -70485 -34238 -70165 -34210
rect -70485 -34862 -70477 -34238
rect -70173 -34862 -70165 -34238
rect -70485 -34890 -70165 -34862
rect -69485 -34238 -69165 -34210
rect -69485 -34862 -69477 -34238
rect -69173 -34862 -69165 -34238
rect -69485 -34890 -69165 -34862
rect -68485 -34238 -68165 -34210
rect -68485 -34862 -68477 -34238
rect -68173 -34862 -68165 -34238
rect -68485 -34890 -68165 -34862
rect -67485 -34238 -67165 -34210
rect -67485 -34862 -67477 -34238
rect -67173 -34862 -67165 -34238
rect -67485 -34890 -67165 -34862
rect -66485 -34238 -66165 -34210
rect -66485 -34862 -66477 -34238
rect -66173 -34862 -66165 -34238
rect -66485 -34890 -66165 -34862
rect -65485 -34238 -65165 -34210
rect -65485 -34862 -65477 -34238
rect -65173 -34862 -65165 -34238
rect -65485 -34890 -65165 -34862
rect -64485 -34238 -64165 -34210
rect -64485 -34862 -64477 -34238
rect -64173 -34862 -64165 -34238
rect -64485 -34890 -64165 -34862
rect -63485 -34238 -63165 -34210
rect -63485 -34862 -63477 -34238
rect -63173 -34862 -63165 -34238
rect -63485 -34890 -63165 -34862
rect -62485 -34238 -62165 -34210
rect -62485 -34862 -62477 -34238
rect -62173 -34862 -62165 -34238
rect -62485 -34890 -62165 -34862
rect -61485 -34238 -61165 -34210
rect -61485 -34862 -61477 -34238
rect -61173 -34862 -61165 -34238
rect -61485 -34890 -61165 -34862
rect -60485 -34238 -60165 -34210
rect -60485 -34862 -60477 -34238
rect -60173 -34862 -60165 -34238
rect -60485 -34890 -60165 -34862
rect -59485 -34238 -59165 -34210
rect -59485 -34862 -59477 -34238
rect -59173 -34862 -59165 -34238
rect -59485 -34890 -59165 -34862
rect -58485 -34238 -58165 -34210
rect -58485 -34862 -58477 -34238
rect -58173 -34862 -58165 -34238
rect -58485 -34890 -58165 -34862
rect -57485 -34238 -57165 -34210
rect -57485 -34862 -57477 -34238
rect -57173 -34862 -57165 -34238
rect -57485 -34890 -57165 -34862
rect -56485 -34238 -56165 -34210
rect -56485 -34862 -56477 -34238
rect -56173 -34862 -56165 -34238
rect -56485 -34890 -56165 -34862
rect -55485 -34238 -55165 -34210
rect -55485 -34862 -55477 -34238
rect -55173 -34862 -55165 -34238
rect -55485 -34890 -55165 -34862
rect -54485 -34238 -54165 -34210
rect -54485 -34862 -54477 -34238
rect -54173 -34862 -54165 -34238
rect -54485 -34890 -54165 -34862
rect -53485 -34238 -53165 -34210
rect -53485 -34862 -53477 -34238
rect -53173 -34862 -53165 -34238
rect -53485 -34890 -53165 -34862
rect -52485 -34238 -52165 -34210
rect -52485 -34862 -52477 -34238
rect -52173 -34862 -52165 -34238
rect -52485 -34890 -52165 -34862
rect -51485 -34238 -51165 -34210
rect -51485 -34862 -51477 -34238
rect -51173 -34862 -51165 -34238
rect -51485 -34890 -51165 -34862
rect -50485 -34238 -50165 -34210
rect -50485 -34862 -50477 -34238
rect -50173 -34862 -50165 -34238
rect -50485 -34890 -50165 -34862
rect -49485 -34238 -49165 -34210
rect -49485 -34862 -49477 -34238
rect -49173 -34862 -49165 -34238
rect -49485 -34890 -49165 -34862
rect -74825 -34898 -48825 -34890
rect -74825 -35202 -74817 -34898
rect -74513 -35202 -74477 -34898
rect -74173 -35202 -74137 -34898
rect -73513 -35202 -73477 -34898
rect -73173 -35202 -73137 -34898
rect -72513 -35202 -72477 -34898
rect -72173 -35202 -72137 -34898
rect -71513 -35202 -71477 -34898
rect -71173 -35202 -71137 -34898
rect -70513 -35202 -70477 -34898
rect -70173 -35202 -70137 -34898
rect -69513 -35202 -69477 -34898
rect -69173 -35202 -69137 -34898
rect -68513 -35202 -68477 -34898
rect -68173 -35202 -68137 -34898
rect -67513 -35202 -67477 -34898
rect -67173 -35202 -67137 -34898
rect -66513 -35202 -66477 -34898
rect -66173 -35202 -66137 -34898
rect -65513 -35202 -65477 -34898
rect -65173 -35202 -65137 -34898
rect -64513 -35202 -64477 -34898
rect -64173 -35202 -64137 -34898
rect -63513 -35202 -63477 -34898
rect -63173 -35202 -63137 -34898
rect -62513 -35202 -62477 -34898
rect -62173 -35202 -62137 -34898
rect -61513 -35202 -61477 -34898
rect -61173 -35202 -61137 -34898
rect -60513 -35202 -60477 -34898
rect -60173 -35202 -60137 -34898
rect -59513 -35202 -59477 -34898
rect -59173 -35202 -59137 -34898
rect -58513 -35202 -58477 -34898
rect -58173 -35202 -58137 -34898
rect -57513 -35202 -57477 -34898
rect -57173 -35202 -57137 -34898
rect -56513 -35202 -56477 -34898
rect -56173 -35202 -56137 -34898
rect -55513 -35202 -55477 -34898
rect -55173 -35202 -55137 -34898
rect -54513 -35202 -54477 -34898
rect -54173 -35202 -54137 -34898
rect -53513 -35202 -53477 -34898
rect -53173 -35202 -53137 -34898
rect -52513 -35202 -52477 -34898
rect -52173 -35202 -52137 -34898
rect -51513 -35202 -51477 -34898
rect -51173 -35202 -51137 -34898
rect -50513 -35202 -50477 -34898
rect -50173 -35202 -50137 -34898
rect -49513 -35202 -49477 -34898
rect -49173 -35202 -49137 -34898
rect -48833 -35202 -48825 -34898
rect -74825 -35210 -48825 -35202
rect -74485 -35238 -74165 -35210
rect -74485 -35862 -74477 -35238
rect -74173 -35862 -74165 -35238
rect -74485 -35890 -74165 -35862
rect -73485 -35238 -73165 -35210
rect -73485 -35862 -73477 -35238
rect -73173 -35862 -73165 -35238
rect -73485 -35890 -73165 -35862
rect -72485 -35238 -72165 -35210
rect -72485 -35862 -72477 -35238
rect -72173 -35862 -72165 -35238
rect -72485 -35890 -72165 -35862
rect -71485 -35238 -71165 -35210
rect -71485 -35862 -71477 -35238
rect -71173 -35862 -71165 -35238
rect -71485 -35890 -71165 -35862
rect -70485 -35238 -70165 -35210
rect -70485 -35862 -70477 -35238
rect -70173 -35862 -70165 -35238
rect -70485 -35890 -70165 -35862
rect -69485 -35238 -69165 -35210
rect -69485 -35862 -69477 -35238
rect -69173 -35862 -69165 -35238
rect -69485 -35890 -69165 -35862
rect -68485 -35238 -68165 -35210
rect -68485 -35862 -68477 -35238
rect -68173 -35862 -68165 -35238
rect -68485 -35890 -68165 -35862
rect -67485 -35238 -67165 -35210
rect -67485 -35862 -67477 -35238
rect -67173 -35862 -67165 -35238
rect -67485 -35890 -67165 -35862
rect -66485 -35238 -66165 -35210
rect -66485 -35862 -66477 -35238
rect -66173 -35862 -66165 -35238
rect -66485 -35890 -66165 -35862
rect -65485 -35238 -65165 -35210
rect -65485 -35862 -65477 -35238
rect -65173 -35862 -65165 -35238
rect -65485 -35890 -65165 -35862
rect -64485 -35238 -64165 -35210
rect -64485 -35862 -64477 -35238
rect -64173 -35862 -64165 -35238
rect -64485 -35890 -64165 -35862
rect -63485 -35238 -63165 -35210
rect -63485 -35862 -63477 -35238
rect -63173 -35862 -63165 -35238
rect -63485 -35890 -63165 -35862
rect -62485 -35238 -62165 -35210
rect -62485 -35862 -62477 -35238
rect -62173 -35862 -62165 -35238
rect -62485 -35890 -62165 -35862
rect -61485 -35238 -61165 -35210
rect -61485 -35862 -61477 -35238
rect -61173 -35862 -61165 -35238
rect -61485 -35890 -61165 -35862
rect -60485 -35238 -60165 -35210
rect -60485 -35862 -60477 -35238
rect -60173 -35862 -60165 -35238
rect -60485 -35890 -60165 -35862
rect -59485 -35238 -59165 -35210
rect -59485 -35862 -59477 -35238
rect -59173 -35862 -59165 -35238
rect -59485 -35890 -59165 -35862
rect -58485 -35238 -58165 -35210
rect -58485 -35862 -58477 -35238
rect -58173 -35862 -58165 -35238
rect -58485 -35890 -58165 -35862
rect -57485 -35238 -57165 -35210
rect -57485 -35862 -57477 -35238
rect -57173 -35862 -57165 -35238
rect -57485 -35890 -57165 -35862
rect -56485 -35238 -56165 -35210
rect -56485 -35862 -56477 -35238
rect -56173 -35862 -56165 -35238
rect -56485 -35890 -56165 -35862
rect -55485 -35238 -55165 -35210
rect -55485 -35862 -55477 -35238
rect -55173 -35862 -55165 -35238
rect -55485 -35890 -55165 -35862
rect -54485 -35238 -54165 -35210
rect -54485 -35862 -54477 -35238
rect -54173 -35862 -54165 -35238
rect -54485 -35890 -54165 -35862
rect -53485 -35238 -53165 -35210
rect -53485 -35862 -53477 -35238
rect -53173 -35862 -53165 -35238
rect -53485 -35890 -53165 -35862
rect -52485 -35238 -52165 -35210
rect -52485 -35862 -52477 -35238
rect -52173 -35862 -52165 -35238
rect -52485 -35890 -52165 -35862
rect -51485 -35238 -51165 -35210
rect -51485 -35862 -51477 -35238
rect -51173 -35862 -51165 -35238
rect -51485 -35890 -51165 -35862
rect -50485 -35238 -50165 -35210
rect -50485 -35862 -50477 -35238
rect -50173 -35862 -50165 -35238
rect -50485 -35890 -50165 -35862
rect -49485 -35238 -49165 -35210
rect -49485 -35862 -49477 -35238
rect -49173 -35862 -49165 -35238
rect -49485 -35890 -49165 -35862
rect -74825 -35898 -48825 -35890
rect -74825 -36202 -74817 -35898
rect -74513 -36202 -74477 -35898
rect -74173 -36202 -74137 -35898
rect -73513 -36202 -73477 -35898
rect -73173 -36202 -73137 -35898
rect -72513 -36202 -72477 -35898
rect -72173 -36202 -72137 -35898
rect -71513 -36202 -71477 -35898
rect -71173 -36202 -71137 -35898
rect -70513 -36202 -70477 -35898
rect -70173 -36202 -70137 -35898
rect -69513 -36202 -69477 -35898
rect -69173 -36202 -69137 -35898
rect -68513 -36202 -68477 -35898
rect -68173 -36202 -68137 -35898
rect -67513 -36202 -67477 -35898
rect -67173 -36202 -67137 -35898
rect -66513 -36202 -66477 -35898
rect -66173 -36202 -66137 -35898
rect -65513 -36202 -65477 -35898
rect -65173 -36202 -65137 -35898
rect -64513 -36202 -64477 -35898
rect -64173 -36202 -64137 -35898
rect -63513 -36202 -63477 -35898
rect -63173 -36202 -63137 -35898
rect -62513 -36202 -62477 -35898
rect -62173 -36202 -62137 -35898
rect -61513 -36202 -61477 -35898
rect -61173 -36202 -61137 -35898
rect -60513 -36202 -60477 -35898
rect -60173 -36202 -60137 -35898
rect -59513 -36202 -59477 -35898
rect -59173 -36202 -59137 -35898
rect -58513 -36202 -58477 -35898
rect -58173 -36202 -58137 -35898
rect -57513 -36202 -57477 -35898
rect -57173 -36202 -57137 -35898
rect -56513 -36202 -56477 -35898
rect -56173 -36202 -56137 -35898
rect -55513 -36202 -55477 -35898
rect -55173 -36202 -55137 -35898
rect -54513 -36202 -54477 -35898
rect -54173 -36202 -54137 -35898
rect -53513 -36202 -53477 -35898
rect -53173 -36202 -53137 -35898
rect -52513 -36202 -52477 -35898
rect -52173 -36202 -52137 -35898
rect -51513 -36202 -51477 -35898
rect -51173 -36202 -51137 -35898
rect -50513 -36202 -50477 -35898
rect -50173 -36202 -50137 -35898
rect -49513 -36202 -49477 -35898
rect -49173 -36202 -49137 -35898
rect -48833 -36202 -48825 -35898
rect -74825 -36210 -48825 -36202
rect -74485 -36238 -74165 -36210
rect -74485 -36862 -74477 -36238
rect -74173 -36862 -74165 -36238
rect -74485 -36890 -74165 -36862
rect -73485 -36238 -73165 -36210
rect -73485 -36862 -73477 -36238
rect -73173 -36862 -73165 -36238
rect -73485 -36890 -73165 -36862
rect -72485 -36238 -72165 -36210
rect -72485 -36862 -72477 -36238
rect -72173 -36862 -72165 -36238
rect -72485 -36890 -72165 -36862
rect -71485 -36238 -71165 -36210
rect -71485 -36862 -71477 -36238
rect -71173 -36862 -71165 -36238
rect -71485 -36890 -71165 -36862
rect -70485 -36238 -70165 -36210
rect -70485 -36862 -70477 -36238
rect -70173 -36862 -70165 -36238
rect -70485 -36890 -70165 -36862
rect -69485 -36238 -69165 -36210
rect -69485 -36862 -69477 -36238
rect -69173 -36862 -69165 -36238
rect -69485 -36890 -69165 -36862
rect -68485 -36238 -68165 -36210
rect -68485 -36862 -68477 -36238
rect -68173 -36862 -68165 -36238
rect -68485 -36890 -68165 -36862
rect -67485 -36238 -67165 -36210
rect -67485 -36862 -67477 -36238
rect -67173 -36862 -67165 -36238
rect -67485 -36890 -67165 -36862
rect -66485 -36238 -66165 -36210
rect -66485 -36862 -66477 -36238
rect -66173 -36862 -66165 -36238
rect -66485 -36890 -66165 -36862
rect -65485 -36238 -65165 -36210
rect -65485 -36862 -65477 -36238
rect -65173 -36862 -65165 -36238
rect -65485 -36890 -65165 -36862
rect -64485 -36238 -64165 -36210
rect -64485 -36862 -64477 -36238
rect -64173 -36862 -64165 -36238
rect -64485 -36890 -64165 -36862
rect -63485 -36238 -63165 -36210
rect -63485 -36862 -63477 -36238
rect -63173 -36862 -63165 -36238
rect -63485 -36890 -63165 -36862
rect -62485 -36238 -62165 -36210
rect -62485 -36862 -62477 -36238
rect -62173 -36862 -62165 -36238
rect -62485 -36890 -62165 -36862
rect -61485 -36238 -61165 -36210
rect -61485 -36862 -61477 -36238
rect -61173 -36862 -61165 -36238
rect -61485 -36890 -61165 -36862
rect -60485 -36238 -60165 -36210
rect -60485 -36862 -60477 -36238
rect -60173 -36862 -60165 -36238
rect -60485 -36890 -60165 -36862
rect -59485 -36238 -59165 -36210
rect -59485 -36862 -59477 -36238
rect -59173 -36862 -59165 -36238
rect -59485 -36890 -59165 -36862
rect -58485 -36238 -58165 -36210
rect -58485 -36862 -58477 -36238
rect -58173 -36862 -58165 -36238
rect -58485 -36890 -58165 -36862
rect -57485 -36238 -57165 -36210
rect -57485 -36862 -57477 -36238
rect -57173 -36862 -57165 -36238
rect -57485 -36890 -57165 -36862
rect -56485 -36238 -56165 -36210
rect -56485 -36862 -56477 -36238
rect -56173 -36862 -56165 -36238
rect -56485 -36890 -56165 -36862
rect -55485 -36238 -55165 -36210
rect -55485 -36862 -55477 -36238
rect -55173 -36862 -55165 -36238
rect -55485 -36890 -55165 -36862
rect -54485 -36238 -54165 -36210
rect -54485 -36862 -54477 -36238
rect -54173 -36862 -54165 -36238
rect -54485 -36890 -54165 -36862
rect -53485 -36238 -53165 -36210
rect -53485 -36862 -53477 -36238
rect -53173 -36862 -53165 -36238
rect -53485 -36890 -53165 -36862
rect -52485 -36238 -52165 -36210
rect -52485 -36862 -52477 -36238
rect -52173 -36862 -52165 -36238
rect -52485 -36890 -52165 -36862
rect -51485 -36238 -51165 -36210
rect -51485 -36862 -51477 -36238
rect -51173 -36862 -51165 -36238
rect -51485 -36890 -51165 -36862
rect -50485 -36238 -50165 -36210
rect -50485 -36862 -50477 -36238
rect -50173 -36862 -50165 -36238
rect -50485 -36890 -50165 -36862
rect -49485 -36238 -49165 -36210
rect -49485 -36862 -49477 -36238
rect -49173 -36862 -49165 -36238
rect -49485 -36890 -49165 -36862
rect -74825 -36898 -48825 -36890
rect -74825 -37202 -74817 -36898
rect -74513 -37202 -74477 -36898
rect -74173 -37202 -74137 -36898
rect -73513 -37202 -73477 -36898
rect -73173 -37202 -73137 -36898
rect -72513 -37202 -72477 -36898
rect -72173 -37202 -72137 -36898
rect -71513 -37202 -71477 -36898
rect -71173 -37202 -71137 -36898
rect -70513 -37202 -70477 -36898
rect -70173 -37202 -70137 -36898
rect -69513 -37202 -69477 -36898
rect -69173 -37202 -69137 -36898
rect -68513 -37202 -68477 -36898
rect -68173 -37202 -68137 -36898
rect -67513 -37202 -67477 -36898
rect -67173 -37202 -67137 -36898
rect -66513 -37202 -66477 -36898
rect -66173 -37202 -66137 -36898
rect -65513 -37202 -65477 -36898
rect -65173 -37202 -65137 -36898
rect -64513 -37202 -64477 -36898
rect -64173 -37202 -64137 -36898
rect -63513 -37202 -63477 -36898
rect -63173 -37202 -63137 -36898
rect -62513 -37202 -62477 -36898
rect -62173 -37202 -62137 -36898
rect -61513 -37202 -61477 -36898
rect -61173 -37202 -61137 -36898
rect -60513 -37202 -60477 -36898
rect -60173 -37202 -60137 -36898
rect -59513 -37202 -59477 -36898
rect -59173 -37202 -59137 -36898
rect -58513 -37202 -58477 -36898
rect -58173 -37202 -58137 -36898
rect -57513 -37202 -57477 -36898
rect -57173 -37202 -57137 -36898
rect -56513 -37202 -56477 -36898
rect -56173 -37202 -56137 -36898
rect -55513 -37202 -55477 -36898
rect -55173 -37202 -55137 -36898
rect -54513 -37202 -54477 -36898
rect -54173 -37202 -54137 -36898
rect -53513 -37202 -53477 -36898
rect -53173 -37202 -53137 -36898
rect -52513 -37202 -52477 -36898
rect -52173 -37202 -52137 -36898
rect -51513 -37202 -51477 -36898
rect -51173 -37202 -51137 -36898
rect -50513 -37202 -50477 -36898
rect -50173 -37202 -50137 -36898
rect -49513 -37202 -49477 -36898
rect -49173 -37202 -49137 -36898
rect -48833 -37202 -48825 -36898
rect -74825 -37210 -48825 -37202
rect -74485 -37238 -74165 -37210
rect -74485 -37862 -74477 -37238
rect -74173 -37862 -74165 -37238
rect -74485 -37890 -74165 -37862
rect -73485 -37238 -73165 -37210
rect -73485 -37862 -73477 -37238
rect -73173 -37862 -73165 -37238
rect -73485 -37890 -73165 -37862
rect -72485 -37238 -72165 -37210
rect -72485 -37862 -72477 -37238
rect -72173 -37862 -72165 -37238
rect -72485 -37890 -72165 -37862
rect -71485 -37238 -71165 -37210
rect -71485 -37862 -71477 -37238
rect -71173 -37862 -71165 -37238
rect -71485 -37890 -71165 -37862
rect -70485 -37238 -70165 -37210
rect -70485 -37862 -70477 -37238
rect -70173 -37862 -70165 -37238
rect -70485 -37890 -70165 -37862
rect -69485 -37238 -69165 -37210
rect -69485 -37862 -69477 -37238
rect -69173 -37862 -69165 -37238
rect -69485 -37890 -69165 -37862
rect -68485 -37238 -68165 -37210
rect -68485 -37862 -68477 -37238
rect -68173 -37862 -68165 -37238
rect -68485 -37890 -68165 -37862
rect -67485 -37238 -67165 -37210
rect -67485 -37862 -67477 -37238
rect -67173 -37862 -67165 -37238
rect -67485 -37890 -67165 -37862
rect -66485 -37238 -66165 -37210
rect -66485 -37862 -66477 -37238
rect -66173 -37862 -66165 -37238
rect -66485 -37890 -66165 -37862
rect -65485 -37238 -65165 -37210
rect -65485 -37862 -65477 -37238
rect -65173 -37862 -65165 -37238
rect -65485 -37890 -65165 -37862
rect -64485 -37238 -64165 -37210
rect -64485 -37862 -64477 -37238
rect -64173 -37862 -64165 -37238
rect -64485 -37890 -64165 -37862
rect -63485 -37238 -63165 -37210
rect -63485 -37862 -63477 -37238
rect -63173 -37862 -63165 -37238
rect -63485 -37890 -63165 -37862
rect -62485 -37238 -62165 -37210
rect -62485 -37862 -62477 -37238
rect -62173 -37862 -62165 -37238
rect -62485 -37890 -62165 -37862
rect -61485 -37238 -61165 -37210
rect -61485 -37862 -61477 -37238
rect -61173 -37862 -61165 -37238
rect -61485 -37890 -61165 -37862
rect -60485 -37238 -60165 -37210
rect -60485 -37862 -60477 -37238
rect -60173 -37862 -60165 -37238
rect -60485 -37890 -60165 -37862
rect -59485 -37238 -59165 -37210
rect -59485 -37862 -59477 -37238
rect -59173 -37862 -59165 -37238
rect -59485 -37890 -59165 -37862
rect -58485 -37238 -58165 -37210
rect -58485 -37862 -58477 -37238
rect -58173 -37862 -58165 -37238
rect -58485 -37890 -58165 -37862
rect -57485 -37238 -57165 -37210
rect -57485 -37862 -57477 -37238
rect -57173 -37862 -57165 -37238
rect -57485 -37890 -57165 -37862
rect -56485 -37238 -56165 -37210
rect -56485 -37862 -56477 -37238
rect -56173 -37862 -56165 -37238
rect -56485 -37890 -56165 -37862
rect -55485 -37238 -55165 -37210
rect -55485 -37862 -55477 -37238
rect -55173 -37862 -55165 -37238
rect -55485 -37890 -55165 -37862
rect -54485 -37238 -54165 -37210
rect -54485 -37862 -54477 -37238
rect -54173 -37862 -54165 -37238
rect -54485 -37890 -54165 -37862
rect -53485 -37238 -53165 -37210
rect -53485 -37862 -53477 -37238
rect -53173 -37862 -53165 -37238
rect -53485 -37890 -53165 -37862
rect -52485 -37238 -52165 -37210
rect -52485 -37862 -52477 -37238
rect -52173 -37862 -52165 -37238
rect -52485 -37890 -52165 -37862
rect -51485 -37238 -51165 -37210
rect -51485 -37862 -51477 -37238
rect -51173 -37862 -51165 -37238
rect -51485 -37890 -51165 -37862
rect -50485 -37238 -50165 -37210
rect -50485 -37862 -50477 -37238
rect -50173 -37862 -50165 -37238
rect -50485 -37890 -50165 -37862
rect -49485 -37238 -49165 -37210
rect -49485 -37862 -49477 -37238
rect -49173 -37862 -49165 -37238
rect -49485 -37890 -49165 -37862
rect -74825 -37898 -48825 -37890
rect -74825 -38202 -74817 -37898
rect -74513 -38202 -74477 -37898
rect -74173 -38202 -74137 -37898
rect -73513 -38202 -73477 -37898
rect -73173 -38202 -73137 -37898
rect -72513 -38202 -72477 -37898
rect -72173 -38202 -72137 -37898
rect -71513 -38202 -71477 -37898
rect -71173 -38202 -71137 -37898
rect -70513 -38202 -70477 -37898
rect -70173 -38202 -70137 -37898
rect -69513 -38202 -69477 -37898
rect -69173 -38202 -69137 -37898
rect -68513 -38202 -68477 -37898
rect -68173 -38202 -68137 -37898
rect -67513 -38202 -67477 -37898
rect -67173 -38202 -67137 -37898
rect -66513 -38202 -66477 -37898
rect -66173 -38202 -66137 -37898
rect -65513 -38202 -65477 -37898
rect -65173 -38202 -65137 -37898
rect -64513 -38202 -64477 -37898
rect -64173 -38202 -64137 -37898
rect -63513 -38202 -63477 -37898
rect -63173 -38202 -63137 -37898
rect -62513 -38202 -62477 -37898
rect -62173 -38202 -62137 -37898
rect -61513 -38202 -61477 -37898
rect -61173 -38202 -61137 -37898
rect -60513 -38202 -60477 -37898
rect -60173 -38202 -60137 -37898
rect -59513 -38202 -59477 -37898
rect -59173 -38202 -59137 -37898
rect -58513 -38202 -58477 -37898
rect -58173 -38202 -58137 -37898
rect -57513 -38202 -57477 -37898
rect -57173 -38202 -57137 -37898
rect -56513 -38202 -56477 -37898
rect -56173 -38202 -56137 -37898
rect -55513 -38202 -55477 -37898
rect -55173 -38202 -55137 -37898
rect -54513 -38202 -54477 -37898
rect -54173 -38202 -54137 -37898
rect -53513 -38202 -53477 -37898
rect -53173 -38202 -53137 -37898
rect -52513 -38202 -52477 -37898
rect -52173 -38202 -52137 -37898
rect -51513 -38202 -51477 -37898
rect -51173 -38202 -51137 -37898
rect -50513 -38202 -50477 -37898
rect -50173 -38202 -50137 -37898
rect -49513 -38202 -49477 -37898
rect -49173 -38202 -49137 -37898
rect -48833 -38202 -48825 -37898
rect -74825 -38210 -48825 -38202
rect -74485 -38238 -74165 -38210
rect -74485 -38862 -74477 -38238
rect -74173 -38862 -74165 -38238
rect -74485 -38890 -74165 -38862
rect -73485 -38238 -73165 -38210
rect -73485 -38862 -73477 -38238
rect -73173 -38862 -73165 -38238
rect -73485 -38890 -73165 -38862
rect -72485 -38238 -72165 -38210
rect -72485 -38862 -72477 -38238
rect -72173 -38862 -72165 -38238
rect -72485 -38890 -72165 -38862
rect -71485 -38238 -71165 -38210
rect -71485 -38862 -71477 -38238
rect -71173 -38862 -71165 -38238
rect -71485 -38890 -71165 -38862
rect -70485 -38238 -70165 -38210
rect -70485 -38862 -70477 -38238
rect -70173 -38862 -70165 -38238
rect -70485 -38890 -70165 -38862
rect -69485 -38238 -69165 -38210
rect -69485 -38862 -69477 -38238
rect -69173 -38862 -69165 -38238
rect -69485 -38890 -69165 -38862
rect -68485 -38238 -68165 -38210
rect -68485 -38862 -68477 -38238
rect -68173 -38862 -68165 -38238
rect -68485 -38890 -68165 -38862
rect -67485 -38238 -67165 -38210
rect -67485 -38862 -67477 -38238
rect -67173 -38862 -67165 -38238
rect -67485 -38890 -67165 -38862
rect -66485 -38238 -66165 -38210
rect -66485 -38862 -66477 -38238
rect -66173 -38862 -66165 -38238
rect -66485 -38890 -66165 -38862
rect -65485 -38238 -65165 -38210
rect -65485 -38862 -65477 -38238
rect -65173 -38862 -65165 -38238
rect -65485 -38890 -65165 -38862
rect -64485 -38238 -64165 -38210
rect -64485 -38862 -64477 -38238
rect -64173 -38862 -64165 -38238
rect -64485 -38890 -64165 -38862
rect -63485 -38238 -63165 -38210
rect -63485 -38862 -63477 -38238
rect -63173 -38862 -63165 -38238
rect -63485 -38890 -63165 -38862
rect -62485 -38238 -62165 -38210
rect -62485 -38862 -62477 -38238
rect -62173 -38862 -62165 -38238
rect -62485 -38890 -62165 -38862
rect -61485 -38238 -61165 -38210
rect -61485 -38862 -61477 -38238
rect -61173 -38862 -61165 -38238
rect -61485 -38890 -61165 -38862
rect -60485 -38238 -60165 -38210
rect -60485 -38862 -60477 -38238
rect -60173 -38862 -60165 -38238
rect -60485 -38890 -60165 -38862
rect -59485 -38238 -59165 -38210
rect -59485 -38862 -59477 -38238
rect -59173 -38862 -59165 -38238
rect -59485 -38890 -59165 -38862
rect -58485 -38238 -58165 -38210
rect -58485 -38862 -58477 -38238
rect -58173 -38862 -58165 -38238
rect -58485 -38890 -58165 -38862
rect -57485 -38238 -57165 -38210
rect -57485 -38862 -57477 -38238
rect -57173 -38862 -57165 -38238
rect -57485 -38890 -57165 -38862
rect -56485 -38238 -56165 -38210
rect -56485 -38862 -56477 -38238
rect -56173 -38862 -56165 -38238
rect -56485 -38890 -56165 -38862
rect -55485 -38238 -55165 -38210
rect -55485 -38862 -55477 -38238
rect -55173 -38862 -55165 -38238
rect -55485 -38890 -55165 -38862
rect -54485 -38238 -54165 -38210
rect -54485 -38862 -54477 -38238
rect -54173 -38862 -54165 -38238
rect -54485 -38890 -54165 -38862
rect -53485 -38238 -53165 -38210
rect -53485 -38862 -53477 -38238
rect -53173 -38862 -53165 -38238
rect -53485 -38890 -53165 -38862
rect -52485 -38238 -52165 -38210
rect -52485 -38862 -52477 -38238
rect -52173 -38862 -52165 -38238
rect -52485 -38890 -52165 -38862
rect -51485 -38238 -51165 -38210
rect -51485 -38862 -51477 -38238
rect -51173 -38862 -51165 -38238
rect -51485 -38890 -51165 -38862
rect -50485 -38238 -50165 -38210
rect -50485 -38862 -50477 -38238
rect -50173 -38862 -50165 -38238
rect -50485 -38890 -50165 -38862
rect -49485 -38238 -49165 -38210
rect -49485 -38862 -49477 -38238
rect -49173 -38862 -49165 -38238
rect -49485 -38890 -49165 -38862
rect -74825 -38898 -48825 -38890
rect -74825 -39202 -74817 -38898
rect -74513 -39202 -74477 -38898
rect -74173 -39202 -74137 -38898
rect -73513 -39202 -73477 -38898
rect -73173 -39202 -73137 -38898
rect -72513 -39202 -72477 -38898
rect -72173 -39202 -72137 -38898
rect -71513 -39202 -71477 -38898
rect -71173 -39202 -71137 -38898
rect -70513 -39202 -70477 -38898
rect -70173 -39202 -70137 -38898
rect -69513 -39202 -69477 -38898
rect -69173 -39202 -69137 -38898
rect -68513 -39202 -68477 -38898
rect -68173 -39202 -68137 -38898
rect -67513 -39202 -67477 -38898
rect -67173 -39202 -67137 -38898
rect -66513 -39202 -66477 -38898
rect -66173 -39202 -66137 -38898
rect -65513 -39202 -65477 -38898
rect -65173 -39202 -65137 -38898
rect -64513 -39202 -64477 -38898
rect -64173 -39202 -64137 -38898
rect -63513 -39202 -63477 -38898
rect -63173 -39202 -63137 -38898
rect -62513 -39202 -62477 -38898
rect -62173 -39202 -62137 -38898
rect -61513 -39202 -61477 -38898
rect -61173 -39202 -61137 -38898
rect -60513 -39202 -60477 -38898
rect -60173 -39202 -60137 -38898
rect -59513 -39202 -59477 -38898
rect -59173 -39202 -59137 -38898
rect -58513 -39202 -58477 -38898
rect -58173 -39202 -58137 -38898
rect -57513 -39202 -57477 -38898
rect -57173 -39202 -57137 -38898
rect -56513 -39202 -56477 -38898
rect -56173 -39202 -56137 -38898
rect -55513 -39202 -55477 -38898
rect -55173 -39202 -55137 -38898
rect -54513 -39202 -54477 -38898
rect -54173 -39202 -54137 -38898
rect -53513 -39202 -53477 -38898
rect -53173 -39202 -53137 -38898
rect -52513 -39202 -52477 -38898
rect -52173 -39202 -52137 -38898
rect -51513 -39202 -51477 -38898
rect -51173 -39202 -51137 -38898
rect -50513 -39202 -50477 -38898
rect -50173 -39202 -50137 -38898
rect -49513 -39202 -49477 -38898
rect -49173 -39202 -49137 -38898
rect -48833 -39202 -48825 -38898
rect -74825 -39210 -48825 -39202
rect -74485 -39238 -74165 -39210
rect -74485 -39862 -74477 -39238
rect -74173 -39862 -74165 -39238
rect -74485 -39890 -74165 -39862
rect -73485 -39238 -73165 -39210
rect -73485 -39862 -73477 -39238
rect -73173 -39862 -73165 -39238
rect -73485 -39890 -73165 -39862
rect -72485 -39238 -72165 -39210
rect -72485 -39862 -72477 -39238
rect -72173 -39862 -72165 -39238
rect -72485 -39890 -72165 -39862
rect -71485 -39238 -71165 -39210
rect -71485 -39862 -71477 -39238
rect -71173 -39862 -71165 -39238
rect -71485 -39890 -71165 -39862
rect -70485 -39238 -70165 -39210
rect -70485 -39862 -70477 -39238
rect -70173 -39862 -70165 -39238
rect -70485 -39890 -70165 -39862
rect -69485 -39238 -69165 -39210
rect -69485 -39862 -69477 -39238
rect -69173 -39862 -69165 -39238
rect -69485 -39890 -69165 -39862
rect -68485 -39238 -68165 -39210
rect -68485 -39862 -68477 -39238
rect -68173 -39862 -68165 -39238
rect -68485 -39890 -68165 -39862
rect -67485 -39238 -67165 -39210
rect -67485 -39862 -67477 -39238
rect -67173 -39862 -67165 -39238
rect -67485 -39890 -67165 -39862
rect -66485 -39238 -66165 -39210
rect -66485 -39862 -66477 -39238
rect -66173 -39862 -66165 -39238
rect -66485 -39890 -66165 -39862
rect -65485 -39238 -65165 -39210
rect -65485 -39862 -65477 -39238
rect -65173 -39862 -65165 -39238
rect -65485 -39890 -65165 -39862
rect -64485 -39238 -64165 -39210
rect -64485 -39862 -64477 -39238
rect -64173 -39862 -64165 -39238
rect -64485 -39890 -64165 -39862
rect -63485 -39238 -63165 -39210
rect -63485 -39862 -63477 -39238
rect -63173 -39862 -63165 -39238
rect -63485 -39890 -63165 -39862
rect -62485 -39238 -62165 -39210
rect -62485 -39862 -62477 -39238
rect -62173 -39862 -62165 -39238
rect -62485 -39890 -62165 -39862
rect -61485 -39238 -61165 -39210
rect -61485 -39862 -61477 -39238
rect -61173 -39862 -61165 -39238
rect -61485 -39890 -61165 -39862
rect -60485 -39238 -60165 -39210
rect -60485 -39862 -60477 -39238
rect -60173 -39862 -60165 -39238
rect -60485 -39890 -60165 -39862
rect -59485 -39238 -59165 -39210
rect -59485 -39862 -59477 -39238
rect -59173 -39862 -59165 -39238
rect -59485 -39890 -59165 -39862
rect -58485 -39238 -58165 -39210
rect -58485 -39862 -58477 -39238
rect -58173 -39862 -58165 -39238
rect -58485 -39890 -58165 -39862
rect -57485 -39238 -57165 -39210
rect -57485 -39862 -57477 -39238
rect -57173 -39862 -57165 -39238
rect -57485 -39890 -57165 -39862
rect -56485 -39238 -56165 -39210
rect -56485 -39862 -56477 -39238
rect -56173 -39862 -56165 -39238
rect -56485 -39890 -56165 -39862
rect -55485 -39238 -55165 -39210
rect -55485 -39862 -55477 -39238
rect -55173 -39862 -55165 -39238
rect -55485 -39890 -55165 -39862
rect -54485 -39238 -54165 -39210
rect -54485 -39862 -54477 -39238
rect -54173 -39862 -54165 -39238
rect -54485 -39890 -54165 -39862
rect -53485 -39238 -53165 -39210
rect -53485 -39862 -53477 -39238
rect -53173 -39862 -53165 -39238
rect -53485 -39890 -53165 -39862
rect -52485 -39238 -52165 -39210
rect -52485 -39862 -52477 -39238
rect -52173 -39862 -52165 -39238
rect -52485 -39890 -52165 -39862
rect -51485 -39238 -51165 -39210
rect -51485 -39862 -51477 -39238
rect -51173 -39862 -51165 -39238
rect -51485 -39890 -51165 -39862
rect -50485 -39238 -50165 -39210
rect -50485 -39862 -50477 -39238
rect -50173 -39862 -50165 -39238
rect -50485 -39890 -50165 -39862
rect -49485 -39238 -49165 -39210
rect -49485 -39862 -49477 -39238
rect -49173 -39862 -49165 -39238
rect -49485 -39890 -49165 -39862
rect -74825 -39898 -48825 -39890
rect -74825 -40202 -74817 -39898
rect -74513 -40202 -74477 -39898
rect -74173 -40202 -74137 -39898
rect -73513 -40202 -73477 -39898
rect -73173 -40202 -73137 -39898
rect -72513 -40202 -72477 -39898
rect -72173 -40202 -72137 -39898
rect -71513 -40202 -71477 -39898
rect -71173 -40202 -71137 -39898
rect -70513 -40202 -70477 -39898
rect -70173 -40202 -70137 -39898
rect -69513 -40202 -69477 -39898
rect -69173 -40202 -69137 -39898
rect -68513 -40202 -68477 -39898
rect -68173 -40202 -68137 -39898
rect -67513 -40202 -67477 -39898
rect -67173 -40202 -67137 -39898
rect -66513 -40202 -66477 -39898
rect -66173 -40202 -66137 -39898
rect -65513 -40202 -65477 -39898
rect -65173 -40202 -65137 -39898
rect -64513 -40202 -64477 -39898
rect -64173 -40202 -64137 -39898
rect -63513 -40202 -63477 -39898
rect -63173 -40202 -63137 -39898
rect -62513 -40202 -62477 -39898
rect -62173 -40202 -62137 -39898
rect -61513 -40202 -61477 -39898
rect -61173 -40202 -61137 -39898
rect -60513 -40202 -60477 -39898
rect -60173 -40202 -60137 -39898
rect -59513 -40202 -59477 -39898
rect -59173 -40202 -59137 -39898
rect -58513 -40202 -58477 -39898
rect -58173 -40202 -58137 -39898
rect -57513 -40202 -57477 -39898
rect -57173 -40202 -57137 -39898
rect -56513 -40202 -56477 -39898
rect -56173 -40202 -56137 -39898
rect -55513 -40202 -55477 -39898
rect -55173 -40202 -55137 -39898
rect -54513 -40202 -54477 -39898
rect -54173 -40202 -54137 -39898
rect -53513 -40202 -53477 -39898
rect -53173 -40202 -53137 -39898
rect -52513 -40202 -52477 -39898
rect -52173 -40202 -52137 -39898
rect -51513 -40202 -51477 -39898
rect -51173 -40202 -51137 -39898
rect -50513 -40202 -50477 -39898
rect -50173 -40202 -50137 -39898
rect -49513 -40202 -49477 -39898
rect -49173 -40202 -49137 -39898
rect -48833 -40202 -48825 -39898
rect -74825 -40210 -48825 -40202
rect -74485 -40238 -74165 -40210
rect -74485 -40862 -74477 -40238
rect -74173 -40862 -74165 -40238
rect -74485 -40890 -74165 -40862
rect -73485 -40238 -73165 -40210
rect -73485 -40862 -73477 -40238
rect -73173 -40862 -73165 -40238
rect -73485 -40890 -73165 -40862
rect -72485 -40238 -72165 -40210
rect -72485 -40862 -72477 -40238
rect -72173 -40862 -72165 -40238
rect -72485 -40890 -72165 -40862
rect -71485 -40238 -71165 -40210
rect -71485 -40862 -71477 -40238
rect -71173 -40862 -71165 -40238
rect -71485 -40890 -71165 -40862
rect -70485 -40238 -70165 -40210
rect -70485 -40862 -70477 -40238
rect -70173 -40862 -70165 -40238
rect -70485 -40890 -70165 -40862
rect -69485 -40238 -69165 -40210
rect -69485 -40862 -69477 -40238
rect -69173 -40862 -69165 -40238
rect -69485 -40890 -69165 -40862
rect -68485 -40238 -68165 -40210
rect -68485 -40862 -68477 -40238
rect -68173 -40862 -68165 -40238
rect -68485 -40890 -68165 -40862
rect -67485 -40238 -67165 -40210
rect -67485 -40862 -67477 -40238
rect -67173 -40862 -67165 -40238
rect -67485 -40890 -67165 -40862
rect -66485 -40238 -66165 -40210
rect -66485 -40862 -66477 -40238
rect -66173 -40862 -66165 -40238
rect -66485 -40890 -66165 -40862
rect -65485 -40238 -65165 -40210
rect -65485 -40862 -65477 -40238
rect -65173 -40862 -65165 -40238
rect -65485 -40890 -65165 -40862
rect -64485 -40238 -64165 -40210
rect -64485 -40862 -64477 -40238
rect -64173 -40862 -64165 -40238
rect -64485 -40890 -64165 -40862
rect -63485 -40238 -63165 -40210
rect -63485 -40862 -63477 -40238
rect -63173 -40862 -63165 -40238
rect -63485 -40890 -63165 -40862
rect -62485 -40238 -62165 -40210
rect -62485 -40862 -62477 -40238
rect -62173 -40862 -62165 -40238
rect -62485 -40890 -62165 -40862
rect -61485 -40238 -61165 -40210
rect -61485 -40862 -61477 -40238
rect -61173 -40862 -61165 -40238
rect -61485 -40890 -61165 -40862
rect -60485 -40238 -60165 -40210
rect -60485 -40862 -60477 -40238
rect -60173 -40862 -60165 -40238
rect -60485 -40890 -60165 -40862
rect -59485 -40238 -59165 -40210
rect -59485 -40862 -59477 -40238
rect -59173 -40862 -59165 -40238
rect -59485 -40890 -59165 -40862
rect -58485 -40238 -58165 -40210
rect -58485 -40862 -58477 -40238
rect -58173 -40862 -58165 -40238
rect -58485 -40890 -58165 -40862
rect -57485 -40238 -57165 -40210
rect -57485 -40862 -57477 -40238
rect -57173 -40862 -57165 -40238
rect -57485 -40890 -57165 -40862
rect -56485 -40238 -56165 -40210
rect -56485 -40862 -56477 -40238
rect -56173 -40862 -56165 -40238
rect -56485 -40890 -56165 -40862
rect -55485 -40238 -55165 -40210
rect -55485 -40862 -55477 -40238
rect -55173 -40862 -55165 -40238
rect -55485 -40890 -55165 -40862
rect -54485 -40238 -54165 -40210
rect -54485 -40862 -54477 -40238
rect -54173 -40862 -54165 -40238
rect -54485 -40890 -54165 -40862
rect -53485 -40238 -53165 -40210
rect -53485 -40862 -53477 -40238
rect -53173 -40862 -53165 -40238
rect -53485 -40890 -53165 -40862
rect -52485 -40238 -52165 -40210
rect -52485 -40862 -52477 -40238
rect -52173 -40862 -52165 -40238
rect -52485 -40890 -52165 -40862
rect -51485 -40238 -51165 -40210
rect -51485 -40862 -51477 -40238
rect -51173 -40862 -51165 -40238
rect -51485 -40890 -51165 -40862
rect -50485 -40238 -50165 -40210
rect -50485 -40862 -50477 -40238
rect -50173 -40862 -50165 -40238
rect -50485 -40890 -50165 -40862
rect -49485 -40238 -49165 -40210
rect -49485 -40862 -49477 -40238
rect -49173 -40862 -49165 -40238
rect -49485 -40890 -49165 -40862
rect -74825 -40898 -48825 -40890
rect -74825 -41202 -74817 -40898
rect -74513 -41202 -74477 -40898
rect -74173 -41202 -74137 -40898
rect -73513 -41202 -73477 -40898
rect -73173 -41202 -73137 -40898
rect -72513 -41202 -72477 -40898
rect -72173 -41202 -72137 -40898
rect -71513 -41202 -71477 -40898
rect -71173 -41202 -71137 -40898
rect -70513 -41202 -70477 -40898
rect -70173 -41202 -70137 -40898
rect -69513 -41202 -69477 -40898
rect -69173 -41202 -69137 -40898
rect -68513 -41202 -68477 -40898
rect -68173 -41202 -68137 -40898
rect -67513 -41202 -67477 -40898
rect -67173 -41202 -67137 -40898
rect -66513 -41202 -66477 -40898
rect -66173 -41202 -66137 -40898
rect -65513 -41202 -65477 -40898
rect -65173 -41202 -65137 -40898
rect -64513 -41202 -64477 -40898
rect -64173 -41202 -64137 -40898
rect -63513 -41202 -63477 -40898
rect -63173 -41202 -63137 -40898
rect -62513 -41202 -62477 -40898
rect -62173 -41202 -62137 -40898
rect -61513 -41202 -61477 -40898
rect -61173 -41202 -61137 -40898
rect -60513 -41202 -60477 -40898
rect -60173 -41202 -60137 -40898
rect -59513 -41202 -59477 -40898
rect -59173 -41202 -59137 -40898
rect -58513 -41202 -58477 -40898
rect -58173 -41202 -58137 -40898
rect -57513 -41202 -57477 -40898
rect -57173 -41202 -57137 -40898
rect -56513 -41202 -56477 -40898
rect -56173 -41202 -56137 -40898
rect -55513 -41202 -55477 -40898
rect -55173 -41202 -55137 -40898
rect -54513 -41202 -54477 -40898
rect -54173 -41202 -54137 -40898
rect -53513 -41202 -53477 -40898
rect -53173 -41202 -53137 -40898
rect -52513 -41202 -52477 -40898
rect -52173 -41202 -52137 -40898
rect -51513 -41202 -51477 -40898
rect -51173 -41202 -51137 -40898
rect -50513 -41202 -50477 -40898
rect -50173 -41202 -50137 -40898
rect -49513 -41202 -49477 -40898
rect -49173 -41202 -49137 -40898
rect -48833 -41202 -48825 -40898
rect -74825 -41210 -48825 -41202
rect -74485 -41238 -74165 -41210
rect -74485 -41862 -74477 -41238
rect -74173 -41862 -74165 -41238
rect -74485 -41890 -74165 -41862
rect -73485 -41238 -73165 -41210
rect -73485 -41862 -73477 -41238
rect -73173 -41862 -73165 -41238
rect -73485 -41890 -73165 -41862
rect -72485 -41238 -72165 -41210
rect -72485 -41862 -72477 -41238
rect -72173 -41862 -72165 -41238
rect -72485 -41890 -72165 -41862
rect -71485 -41238 -71165 -41210
rect -71485 -41862 -71477 -41238
rect -71173 -41862 -71165 -41238
rect -71485 -41890 -71165 -41862
rect -70485 -41238 -70165 -41210
rect -70485 -41862 -70477 -41238
rect -70173 -41862 -70165 -41238
rect -70485 -41890 -70165 -41862
rect -69485 -41238 -69165 -41210
rect -69485 -41862 -69477 -41238
rect -69173 -41862 -69165 -41238
rect -69485 -41890 -69165 -41862
rect -68485 -41238 -68165 -41210
rect -68485 -41862 -68477 -41238
rect -68173 -41862 -68165 -41238
rect -68485 -41890 -68165 -41862
rect -67485 -41238 -67165 -41210
rect -67485 -41862 -67477 -41238
rect -67173 -41862 -67165 -41238
rect -67485 -41890 -67165 -41862
rect -66485 -41238 -66165 -41210
rect -66485 -41862 -66477 -41238
rect -66173 -41862 -66165 -41238
rect -66485 -41890 -66165 -41862
rect -65485 -41238 -65165 -41210
rect -65485 -41862 -65477 -41238
rect -65173 -41862 -65165 -41238
rect -65485 -41890 -65165 -41862
rect -64485 -41238 -64165 -41210
rect -64485 -41862 -64477 -41238
rect -64173 -41862 -64165 -41238
rect -64485 -41890 -64165 -41862
rect -63485 -41238 -63165 -41210
rect -63485 -41862 -63477 -41238
rect -63173 -41862 -63165 -41238
rect -63485 -41890 -63165 -41862
rect -62485 -41238 -62165 -41210
rect -62485 -41862 -62477 -41238
rect -62173 -41862 -62165 -41238
rect -62485 -41890 -62165 -41862
rect -61485 -41238 -61165 -41210
rect -61485 -41862 -61477 -41238
rect -61173 -41862 -61165 -41238
rect -61485 -41890 -61165 -41862
rect -60485 -41238 -60165 -41210
rect -60485 -41862 -60477 -41238
rect -60173 -41862 -60165 -41238
rect -60485 -41890 -60165 -41862
rect -59485 -41238 -59165 -41210
rect -59485 -41862 -59477 -41238
rect -59173 -41862 -59165 -41238
rect -59485 -41890 -59165 -41862
rect -58485 -41238 -58165 -41210
rect -58485 -41862 -58477 -41238
rect -58173 -41862 -58165 -41238
rect -58485 -41890 -58165 -41862
rect -57485 -41238 -57165 -41210
rect -57485 -41862 -57477 -41238
rect -57173 -41862 -57165 -41238
rect -57485 -41890 -57165 -41862
rect -56485 -41238 -56165 -41210
rect -56485 -41862 -56477 -41238
rect -56173 -41862 -56165 -41238
rect -56485 -41890 -56165 -41862
rect -55485 -41238 -55165 -41210
rect -55485 -41862 -55477 -41238
rect -55173 -41862 -55165 -41238
rect -55485 -41890 -55165 -41862
rect -54485 -41238 -54165 -41210
rect -54485 -41862 -54477 -41238
rect -54173 -41862 -54165 -41238
rect -54485 -41890 -54165 -41862
rect -53485 -41238 -53165 -41210
rect -53485 -41862 -53477 -41238
rect -53173 -41862 -53165 -41238
rect -53485 -41890 -53165 -41862
rect -52485 -41238 -52165 -41210
rect -52485 -41862 -52477 -41238
rect -52173 -41862 -52165 -41238
rect -52485 -41890 -52165 -41862
rect -51485 -41238 -51165 -41210
rect -51485 -41862 -51477 -41238
rect -51173 -41862 -51165 -41238
rect -51485 -41890 -51165 -41862
rect -50485 -41238 -50165 -41210
rect -50485 -41862 -50477 -41238
rect -50173 -41862 -50165 -41238
rect -50485 -41890 -50165 -41862
rect -49485 -41238 -49165 -41210
rect -49485 -41862 -49477 -41238
rect -49173 -41862 -49165 -41238
rect -49485 -41890 -49165 -41862
rect -74825 -41898 -48825 -41890
rect -74825 -42202 -74817 -41898
rect -74513 -42202 -74477 -41898
rect -74173 -42202 -74137 -41898
rect -73513 -42202 -73477 -41898
rect -73173 -42202 -73137 -41898
rect -72513 -42202 -72477 -41898
rect -72173 -42202 -72137 -41898
rect -71513 -42202 -71477 -41898
rect -71173 -42202 -71137 -41898
rect -70513 -42202 -70477 -41898
rect -70173 -42202 -70137 -41898
rect -69513 -42202 -69477 -41898
rect -69173 -42202 -69137 -41898
rect -68513 -42202 -68477 -41898
rect -68173 -42202 -68137 -41898
rect -67513 -42202 -67477 -41898
rect -67173 -42202 -67137 -41898
rect -66513 -42202 -66477 -41898
rect -66173 -42202 -66137 -41898
rect -65513 -42202 -65477 -41898
rect -65173 -42202 -65137 -41898
rect -64513 -42202 -64477 -41898
rect -64173 -42202 -64137 -41898
rect -63513 -42202 -63477 -41898
rect -63173 -42202 -63137 -41898
rect -62513 -42202 -62477 -41898
rect -62173 -42202 -62137 -41898
rect -61513 -42202 -61477 -41898
rect -61173 -42202 -61137 -41898
rect -60513 -42202 -60477 -41898
rect -60173 -42202 -60137 -41898
rect -59513 -42202 -59477 -41898
rect -59173 -42202 -59137 -41898
rect -58513 -42202 -58477 -41898
rect -58173 -42202 -58137 -41898
rect -57513 -42202 -57477 -41898
rect -57173 -42202 -57137 -41898
rect -56513 -42202 -56477 -41898
rect -56173 -42202 -56137 -41898
rect -55513 -42202 -55477 -41898
rect -55173 -42202 -55137 -41898
rect -54513 -42202 -54477 -41898
rect -54173 -42202 -54137 -41898
rect -53513 -42202 -53477 -41898
rect -53173 -42202 -53137 -41898
rect -52513 -42202 -52477 -41898
rect -52173 -42202 -52137 -41898
rect -51513 -42202 -51477 -41898
rect -51173 -42202 -51137 -41898
rect -50513 -42202 -50477 -41898
rect -50173 -42202 -50137 -41898
rect -49513 -42202 -49477 -41898
rect -49173 -42202 -49137 -41898
rect -48833 -42202 -48825 -41898
rect -74825 -42210 -48825 -42202
rect -74485 -42238 -74165 -42210
rect -74485 -42862 -74477 -42238
rect -74173 -42862 -74165 -42238
rect -74485 -42890 -74165 -42862
rect -73485 -42238 -73165 -42210
rect -73485 -42862 -73477 -42238
rect -73173 -42862 -73165 -42238
rect -73485 -42890 -73165 -42862
rect -72485 -42238 -72165 -42210
rect -72485 -42862 -72477 -42238
rect -72173 -42862 -72165 -42238
rect -72485 -42890 -72165 -42862
rect -71485 -42238 -71165 -42210
rect -71485 -42862 -71477 -42238
rect -71173 -42862 -71165 -42238
rect -71485 -42890 -71165 -42862
rect -70485 -42238 -70165 -42210
rect -70485 -42862 -70477 -42238
rect -70173 -42862 -70165 -42238
rect -70485 -42890 -70165 -42862
rect -69485 -42238 -69165 -42210
rect -69485 -42862 -69477 -42238
rect -69173 -42862 -69165 -42238
rect -69485 -42890 -69165 -42862
rect -68485 -42238 -68165 -42210
rect -68485 -42862 -68477 -42238
rect -68173 -42862 -68165 -42238
rect -68485 -42890 -68165 -42862
rect -67485 -42238 -67165 -42210
rect -67485 -42862 -67477 -42238
rect -67173 -42862 -67165 -42238
rect -67485 -42890 -67165 -42862
rect -66485 -42238 -66165 -42210
rect -66485 -42862 -66477 -42238
rect -66173 -42862 -66165 -42238
rect -66485 -42890 -66165 -42862
rect -65485 -42238 -65165 -42210
rect -65485 -42862 -65477 -42238
rect -65173 -42862 -65165 -42238
rect -65485 -42890 -65165 -42862
rect -64485 -42238 -64165 -42210
rect -64485 -42862 -64477 -42238
rect -64173 -42862 -64165 -42238
rect -64485 -42890 -64165 -42862
rect -63485 -42238 -63165 -42210
rect -63485 -42862 -63477 -42238
rect -63173 -42862 -63165 -42238
rect -63485 -42890 -63165 -42862
rect -62485 -42238 -62165 -42210
rect -62485 -42862 -62477 -42238
rect -62173 -42862 -62165 -42238
rect -62485 -42890 -62165 -42862
rect -61485 -42238 -61165 -42210
rect -61485 -42862 -61477 -42238
rect -61173 -42862 -61165 -42238
rect -61485 -42890 -61165 -42862
rect -60485 -42238 -60165 -42210
rect -60485 -42862 -60477 -42238
rect -60173 -42862 -60165 -42238
rect -60485 -42890 -60165 -42862
rect -59485 -42238 -59165 -42210
rect -59485 -42862 -59477 -42238
rect -59173 -42862 -59165 -42238
rect -59485 -42890 -59165 -42862
rect -58485 -42238 -58165 -42210
rect -58485 -42862 -58477 -42238
rect -58173 -42862 -58165 -42238
rect -58485 -42890 -58165 -42862
rect -57485 -42238 -57165 -42210
rect -57485 -42862 -57477 -42238
rect -57173 -42862 -57165 -42238
rect -57485 -42890 -57165 -42862
rect -56485 -42238 -56165 -42210
rect -56485 -42862 -56477 -42238
rect -56173 -42862 -56165 -42238
rect -56485 -42890 -56165 -42862
rect -55485 -42238 -55165 -42210
rect -55485 -42862 -55477 -42238
rect -55173 -42862 -55165 -42238
rect -55485 -42890 -55165 -42862
rect -54485 -42238 -54165 -42210
rect -54485 -42862 -54477 -42238
rect -54173 -42862 -54165 -42238
rect -54485 -42890 -54165 -42862
rect -53485 -42238 -53165 -42210
rect -53485 -42862 -53477 -42238
rect -53173 -42862 -53165 -42238
rect -53485 -42890 -53165 -42862
rect -52485 -42238 -52165 -42210
rect -52485 -42862 -52477 -42238
rect -52173 -42862 -52165 -42238
rect -52485 -42890 -52165 -42862
rect -51485 -42238 -51165 -42210
rect -51485 -42862 -51477 -42238
rect -51173 -42862 -51165 -42238
rect -51485 -42890 -51165 -42862
rect -50485 -42238 -50165 -42210
rect -50485 -42862 -50477 -42238
rect -50173 -42862 -50165 -42238
rect -50485 -42890 -50165 -42862
rect -49485 -42238 -49165 -42210
rect -49485 -42862 -49477 -42238
rect -49173 -42862 -49165 -42238
rect -49485 -42890 -49165 -42862
rect -74825 -42898 -48825 -42890
rect -74825 -43202 -74817 -42898
rect -74513 -43202 -74477 -42898
rect -74173 -43202 -74137 -42898
rect -73513 -43202 -73477 -42898
rect -73173 -43202 -73137 -42898
rect -72513 -43202 -72477 -42898
rect -72173 -43202 -72137 -42898
rect -71513 -43202 -71477 -42898
rect -71173 -43202 -71137 -42898
rect -70513 -43202 -70477 -42898
rect -70173 -43202 -70137 -42898
rect -69513 -43202 -69477 -42898
rect -69173 -43202 -69137 -42898
rect -68513 -43202 -68477 -42898
rect -68173 -43202 -68137 -42898
rect -67513 -43202 -67477 -42898
rect -67173 -43202 -67137 -42898
rect -66513 -43202 -66477 -42898
rect -66173 -43202 -66137 -42898
rect -65513 -43202 -65477 -42898
rect -65173 -43202 -65137 -42898
rect -64513 -43202 -64477 -42898
rect -64173 -43202 -64137 -42898
rect -63513 -43202 -63477 -42898
rect -63173 -43202 -63137 -42898
rect -62513 -43202 -62477 -42898
rect -62173 -43202 -62137 -42898
rect -61513 -43202 -61477 -42898
rect -61173 -43202 -61137 -42898
rect -60513 -43202 -60477 -42898
rect -60173 -43202 -60137 -42898
rect -59513 -43202 -59477 -42898
rect -59173 -43202 -59137 -42898
rect -58513 -43202 -58477 -42898
rect -58173 -43202 -58137 -42898
rect -57513 -43202 -57477 -42898
rect -57173 -43202 -57137 -42898
rect -56513 -43202 -56477 -42898
rect -56173 -43202 -56137 -42898
rect -55513 -43202 -55477 -42898
rect -55173 -43202 -55137 -42898
rect -54513 -43202 -54477 -42898
rect -54173 -43202 -54137 -42898
rect -53513 -43202 -53477 -42898
rect -53173 -43202 -53137 -42898
rect -52513 -43202 -52477 -42898
rect -52173 -43202 -52137 -42898
rect -51513 -43202 -51477 -42898
rect -51173 -43202 -51137 -42898
rect -50513 -43202 -50477 -42898
rect -50173 -43202 -50137 -42898
rect -49513 -43202 -49477 -42898
rect -49173 -43202 -49137 -42898
rect -48833 -43202 -48825 -42898
rect -74825 -43210 -48825 -43202
rect -74485 -43238 -74165 -43210
rect -74485 -43862 -74477 -43238
rect -74173 -43862 -74165 -43238
rect -74485 -43890 -74165 -43862
rect -73485 -43238 -73165 -43210
rect -73485 -43862 -73477 -43238
rect -73173 -43862 -73165 -43238
rect -73485 -43890 -73165 -43862
rect -72485 -43238 -72165 -43210
rect -72485 -43862 -72477 -43238
rect -72173 -43862 -72165 -43238
rect -72485 -43890 -72165 -43862
rect -71485 -43238 -71165 -43210
rect -71485 -43862 -71477 -43238
rect -71173 -43862 -71165 -43238
rect -71485 -43890 -71165 -43862
rect -70485 -43238 -70165 -43210
rect -70485 -43862 -70477 -43238
rect -70173 -43862 -70165 -43238
rect -70485 -43890 -70165 -43862
rect -69485 -43238 -69165 -43210
rect -69485 -43862 -69477 -43238
rect -69173 -43862 -69165 -43238
rect -69485 -43890 -69165 -43862
rect -68485 -43238 -68165 -43210
rect -68485 -43862 -68477 -43238
rect -68173 -43862 -68165 -43238
rect -68485 -43890 -68165 -43862
rect -67485 -43238 -67165 -43210
rect -67485 -43862 -67477 -43238
rect -67173 -43862 -67165 -43238
rect -67485 -43890 -67165 -43862
rect -66485 -43238 -66165 -43210
rect -66485 -43862 -66477 -43238
rect -66173 -43862 -66165 -43238
rect -66485 -43890 -66165 -43862
rect -65485 -43238 -65165 -43210
rect -65485 -43862 -65477 -43238
rect -65173 -43862 -65165 -43238
rect -65485 -43890 -65165 -43862
rect -64485 -43238 -64165 -43210
rect -64485 -43862 -64477 -43238
rect -64173 -43862 -64165 -43238
rect -64485 -43890 -64165 -43862
rect -63485 -43238 -63165 -43210
rect -63485 -43862 -63477 -43238
rect -63173 -43862 -63165 -43238
rect -63485 -43890 -63165 -43862
rect -62485 -43238 -62165 -43210
rect -62485 -43862 -62477 -43238
rect -62173 -43862 -62165 -43238
rect -62485 -43890 -62165 -43862
rect -61485 -43238 -61165 -43210
rect -61485 -43862 -61477 -43238
rect -61173 -43862 -61165 -43238
rect -61485 -43890 -61165 -43862
rect -60485 -43238 -60165 -43210
rect -60485 -43862 -60477 -43238
rect -60173 -43862 -60165 -43238
rect -60485 -43890 -60165 -43862
rect -59485 -43238 -59165 -43210
rect -59485 -43862 -59477 -43238
rect -59173 -43862 -59165 -43238
rect -59485 -43890 -59165 -43862
rect -58485 -43238 -58165 -43210
rect -58485 -43862 -58477 -43238
rect -58173 -43862 -58165 -43238
rect -58485 -43890 -58165 -43862
rect -57485 -43238 -57165 -43210
rect -57485 -43862 -57477 -43238
rect -57173 -43862 -57165 -43238
rect -57485 -43890 -57165 -43862
rect -56485 -43238 -56165 -43210
rect -56485 -43862 -56477 -43238
rect -56173 -43862 -56165 -43238
rect -56485 -43890 -56165 -43862
rect -55485 -43238 -55165 -43210
rect -55485 -43862 -55477 -43238
rect -55173 -43862 -55165 -43238
rect -55485 -43890 -55165 -43862
rect -54485 -43238 -54165 -43210
rect -54485 -43862 -54477 -43238
rect -54173 -43862 -54165 -43238
rect -54485 -43890 -54165 -43862
rect -53485 -43238 -53165 -43210
rect -53485 -43862 -53477 -43238
rect -53173 -43862 -53165 -43238
rect -53485 -43890 -53165 -43862
rect -52485 -43238 -52165 -43210
rect -52485 -43862 -52477 -43238
rect -52173 -43862 -52165 -43238
rect -52485 -43890 -52165 -43862
rect -51485 -43238 -51165 -43210
rect -51485 -43862 -51477 -43238
rect -51173 -43862 -51165 -43238
rect -51485 -43890 -51165 -43862
rect -50485 -43238 -50165 -43210
rect -50485 -43862 -50477 -43238
rect -50173 -43862 -50165 -43238
rect -50485 -43890 -50165 -43862
rect -49485 -43238 -49165 -43210
rect -49485 -43862 -49477 -43238
rect -49173 -43862 -49165 -43238
rect -49485 -43890 -49165 -43862
rect -74825 -43898 -48825 -43890
rect -74825 -44202 -74817 -43898
rect -74513 -44202 -74477 -43898
rect -74173 -44202 -74137 -43898
rect -73513 -44202 -73477 -43898
rect -73173 -44202 -73137 -43898
rect -72513 -44202 -72477 -43898
rect -72173 -44202 -72137 -43898
rect -71513 -44202 -71477 -43898
rect -71173 -44202 -71137 -43898
rect -70513 -44202 -70477 -43898
rect -70173 -44202 -70137 -43898
rect -69513 -44202 -69477 -43898
rect -69173 -44202 -69137 -43898
rect -68513 -44202 -68477 -43898
rect -68173 -44202 -68137 -43898
rect -67513 -44202 -67477 -43898
rect -67173 -44202 -67137 -43898
rect -66513 -44202 -66477 -43898
rect -66173 -44202 -66137 -43898
rect -65513 -44202 -65477 -43898
rect -65173 -44202 -65137 -43898
rect -64513 -44202 -64477 -43898
rect -64173 -44202 -64137 -43898
rect -63513 -44202 -63477 -43898
rect -63173 -44202 -63137 -43898
rect -62513 -44202 -62477 -43898
rect -62173 -44202 -62137 -43898
rect -61513 -44202 -61477 -43898
rect -61173 -44202 -61137 -43898
rect -60513 -44202 -60477 -43898
rect -60173 -44202 -60137 -43898
rect -59513 -44202 -59477 -43898
rect -59173 -44202 -59137 -43898
rect -58513 -44202 -58477 -43898
rect -58173 -44202 -58137 -43898
rect -57513 -44202 -57477 -43898
rect -57173 -44202 -57137 -43898
rect -56513 -44202 -56477 -43898
rect -56173 -44202 -56137 -43898
rect -55513 -44202 -55477 -43898
rect -55173 -44202 -55137 -43898
rect -54513 -44202 -54477 -43898
rect -54173 -44202 -54137 -43898
rect -53513 -44202 -53477 -43898
rect -53173 -44202 -53137 -43898
rect -52513 -44202 -52477 -43898
rect -52173 -44202 -52137 -43898
rect -51513 -44202 -51477 -43898
rect -51173 -44202 -51137 -43898
rect -50513 -44202 -50477 -43898
rect -50173 -44202 -50137 -43898
rect -49513 -44202 -49477 -43898
rect -49173 -44202 -49137 -43898
rect -48833 -44202 -48825 -43898
rect -74825 -44210 -48825 -44202
rect -74485 -44238 -74165 -44210
rect -74485 -44862 -74477 -44238
rect -74173 -44862 -74165 -44238
rect -74485 -44890 -74165 -44862
rect -73485 -44238 -73165 -44210
rect -73485 -44862 -73477 -44238
rect -73173 -44862 -73165 -44238
rect -73485 -44890 -73165 -44862
rect -72485 -44238 -72165 -44210
rect -72485 -44862 -72477 -44238
rect -72173 -44862 -72165 -44238
rect -72485 -44890 -72165 -44862
rect -71485 -44238 -71165 -44210
rect -71485 -44862 -71477 -44238
rect -71173 -44862 -71165 -44238
rect -71485 -44890 -71165 -44862
rect -70485 -44238 -70165 -44210
rect -70485 -44862 -70477 -44238
rect -70173 -44862 -70165 -44238
rect -70485 -44890 -70165 -44862
rect -69485 -44238 -69165 -44210
rect -69485 -44862 -69477 -44238
rect -69173 -44862 -69165 -44238
rect -69485 -44890 -69165 -44862
rect -68485 -44238 -68165 -44210
rect -68485 -44862 -68477 -44238
rect -68173 -44862 -68165 -44238
rect -68485 -44890 -68165 -44862
rect -67485 -44238 -67165 -44210
rect -67485 -44862 -67477 -44238
rect -67173 -44862 -67165 -44238
rect -67485 -44890 -67165 -44862
rect -66485 -44238 -66165 -44210
rect -66485 -44862 -66477 -44238
rect -66173 -44862 -66165 -44238
rect -66485 -44890 -66165 -44862
rect -65485 -44238 -65165 -44210
rect -65485 -44862 -65477 -44238
rect -65173 -44862 -65165 -44238
rect -65485 -44890 -65165 -44862
rect -64485 -44238 -64165 -44210
rect -64485 -44862 -64477 -44238
rect -64173 -44862 -64165 -44238
rect -64485 -44890 -64165 -44862
rect -63485 -44238 -63165 -44210
rect -63485 -44862 -63477 -44238
rect -63173 -44862 -63165 -44238
rect -63485 -44890 -63165 -44862
rect -62485 -44238 -62165 -44210
rect -62485 -44862 -62477 -44238
rect -62173 -44862 -62165 -44238
rect -62485 -44890 -62165 -44862
rect -61485 -44238 -61165 -44210
rect -61485 -44862 -61477 -44238
rect -61173 -44862 -61165 -44238
rect -61485 -44890 -61165 -44862
rect -60485 -44238 -60165 -44210
rect -60485 -44862 -60477 -44238
rect -60173 -44862 -60165 -44238
rect -60485 -44890 -60165 -44862
rect -59485 -44238 -59165 -44210
rect -59485 -44862 -59477 -44238
rect -59173 -44862 -59165 -44238
rect -59485 -44890 -59165 -44862
rect -58485 -44238 -58165 -44210
rect -58485 -44862 -58477 -44238
rect -58173 -44862 -58165 -44238
rect -58485 -44890 -58165 -44862
rect -57485 -44238 -57165 -44210
rect -57485 -44862 -57477 -44238
rect -57173 -44862 -57165 -44238
rect -57485 -44890 -57165 -44862
rect -56485 -44238 -56165 -44210
rect -56485 -44862 -56477 -44238
rect -56173 -44862 -56165 -44238
rect -56485 -44890 -56165 -44862
rect -55485 -44238 -55165 -44210
rect -55485 -44862 -55477 -44238
rect -55173 -44862 -55165 -44238
rect -55485 -44890 -55165 -44862
rect -54485 -44238 -54165 -44210
rect -54485 -44862 -54477 -44238
rect -54173 -44862 -54165 -44238
rect -54485 -44890 -54165 -44862
rect -53485 -44238 -53165 -44210
rect -53485 -44862 -53477 -44238
rect -53173 -44862 -53165 -44238
rect -53485 -44890 -53165 -44862
rect -52485 -44238 -52165 -44210
rect -52485 -44862 -52477 -44238
rect -52173 -44862 -52165 -44238
rect -52485 -44890 -52165 -44862
rect -51485 -44238 -51165 -44210
rect -51485 -44862 -51477 -44238
rect -51173 -44862 -51165 -44238
rect -51485 -44890 -51165 -44862
rect -50485 -44238 -50165 -44210
rect -50485 -44862 -50477 -44238
rect -50173 -44862 -50165 -44238
rect -50485 -44890 -50165 -44862
rect -49485 -44238 -49165 -44210
rect -49485 -44862 -49477 -44238
rect -49173 -44862 -49165 -44238
rect -46275 -44502 -46232 -32598
rect -36328 -44502 -36275 -32598
rect -46275 -44550 -36275 -44502
rect -4275 -32598 5725 -32550
rect -4275 -44502 -4232 -32598
rect 5672 -44502 5725 -32598
rect 8615 -32862 8623 -32238
rect 8927 -32862 8935 -32238
rect 8615 -32890 8935 -32862
rect 9615 -32238 9935 -32210
rect 9615 -32862 9623 -32238
rect 9927 -32862 9935 -32238
rect 9615 -32890 9935 -32862
rect 10615 -32238 10935 -32210
rect 10615 -32862 10623 -32238
rect 10927 -32862 10935 -32238
rect 10615 -32890 10935 -32862
rect 11615 -32238 11935 -32210
rect 11615 -32862 11623 -32238
rect 11927 -32862 11935 -32238
rect 11615 -32890 11935 -32862
rect 12615 -32238 12935 -32210
rect 12615 -32862 12623 -32238
rect 12927 -32862 12935 -32238
rect 12615 -32890 12935 -32862
rect 13615 -32238 13935 -32210
rect 13615 -32862 13623 -32238
rect 13927 -32862 13935 -32238
rect 13615 -32890 13935 -32862
rect 14615 -32238 14935 -32210
rect 14615 -32862 14623 -32238
rect 14927 -32862 14935 -32238
rect 14615 -32890 14935 -32862
rect 15615 -32238 15935 -32210
rect 15615 -32862 15623 -32238
rect 15927 -32862 15935 -32238
rect 15615 -32890 15935 -32862
rect 16615 -32238 16935 -32210
rect 16615 -32862 16623 -32238
rect 16927 -32862 16935 -32238
rect 16615 -32890 16935 -32862
rect 17615 -32238 17935 -32210
rect 17615 -32862 17623 -32238
rect 17927 -32862 17935 -32238
rect 17615 -32890 17935 -32862
rect 18615 -32238 18935 -32210
rect 18615 -32862 18623 -32238
rect 18927 -32862 18935 -32238
rect 18615 -32890 18935 -32862
rect 19615 -32238 19935 -32210
rect 19615 -32862 19623 -32238
rect 19927 -32862 19935 -32238
rect 19615 -32890 19935 -32862
rect 20615 -32238 20935 -32210
rect 20615 -32862 20623 -32238
rect 20927 -32862 20935 -32238
rect 20615 -32890 20935 -32862
rect 21615 -32238 21935 -32210
rect 21615 -32862 21623 -32238
rect 21927 -32862 21935 -32238
rect 21615 -32890 21935 -32862
rect 22615 -32238 22935 -32210
rect 22615 -32862 22623 -32238
rect 22927 -32862 22935 -32238
rect 22615 -32890 22935 -32862
rect 23615 -32238 23935 -32210
rect 23615 -32862 23623 -32238
rect 23927 -32862 23935 -32238
rect 23615 -32890 23935 -32862
rect 24615 -32238 24935 -32210
rect 24615 -32862 24623 -32238
rect 24927 -32862 24935 -32238
rect 24615 -32890 24935 -32862
rect 25615 -32238 25935 -32210
rect 25615 -32862 25623 -32238
rect 25927 -32862 25935 -32238
rect 25615 -32890 25935 -32862
rect 26615 -32238 26935 -32210
rect 26615 -32862 26623 -32238
rect 26927 -32862 26935 -32238
rect 26615 -32890 26935 -32862
rect 27615 -32238 27935 -32210
rect 27615 -32862 27623 -32238
rect 27927 -32862 27935 -32238
rect 27615 -32890 27935 -32862
rect 28615 -32238 28935 -32210
rect 28615 -32862 28623 -32238
rect 28927 -32862 28935 -32238
rect 28615 -32890 28935 -32862
rect 29615 -32238 29935 -32210
rect 29615 -32862 29623 -32238
rect 29927 -32862 29935 -32238
rect 29615 -32890 29935 -32862
rect 30615 -32238 30935 -32210
rect 30615 -32862 30623 -32238
rect 30927 -32862 30935 -32238
rect 30615 -32890 30935 -32862
rect 31615 -32238 31935 -32210
rect 31615 -32862 31623 -32238
rect 31927 -32862 31935 -32238
rect 31615 -32890 31935 -32862
rect 32615 -32238 32935 -32210
rect 32615 -32862 32623 -32238
rect 32927 -32862 32935 -32238
rect 32615 -32890 32935 -32862
rect 33615 -32238 33935 -32210
rect 33615 -32862 33623 -32238
rect 33927 -32862 33935 -32238
rect 33615 -32890 33935 -32862
rect 8275 -32898 34275 -32890
rect 8275 -33202 8283 -32898
rect 8587 -33202 8623 -32898
rect 8927 -33202 8963 -32898
rect 9587 -33202 9623 -32898
rect 9927 -33202 9963 -32898
rect 10587 -33202 10623 -32898
rect 10927 -33202 10963 -32898
rect 11587 -33202 11623 -32898
rect 11927 -33202 11963 -32898
rect 12587 -33202 12623 -32898
rect 12927 -33202 12963 -32898
rect 13587 -33202 13623 -32898
rect 13927 -33202 13963 -32898
rect 14587 -33202 14623 -32898
rect 14927 -33202 14963 -32898
rect 15587 -33202 15623 -32898
rect 15927 -33202 15963 -32898
rect 16587 -33202 16623 -32898
rect 16927 -33202 16963 -32898
rect 17587 -33202 17623 -32898
rect 17927 -33202 17963 -32898
rect 18587 -33202 18623 -32898
rect 18927 -33202 18963 -32898
rect 19587 -33202 19623 -32898
rect 19927 -33202 19963 -32898
rect 20587 -33202 20623 -32898
rect 20927 -33202 20963 -32898
rect 21587 -33202 21623 -32898
rect 21927 -33202 21963 -32898
rect 22587 -33202 22623 -32898
rect 22927 -33202 22963 -32898
rect 23587 -33202 23623 -32898
rect 23927 -33202 23963 -32898
rect 24587 -33202 24623 -32898
rect 24927 -33202 24963 -32898
rect 25587 -33202 25623 -32898
rect 25927 -33202 25963 -32898
rect 26587 -33202 26623 -32898
rect 26927 -33202 26963 -32898
rect 27587 -33202 27623 -32898
rect 27927 -33202 27963 -32898
rect 28587 -33202 28623 -32898
rect 28927 -33202 28963 -32898
rect 29587 -33202 29623 -32898
rect 29927 -33202 29963 -32898
rect 30587 -33202 30623 -32898
rect 30927 -33202 30963 -32898
rect 31587 -33202 31623 -32898
rect 31927 -33202 31963 -32898
rect 32587 -33202 32623 -32898
rect 32927 -33202 32963 -32898
rect 33587 -33202 33623 -32898
rect 33927 -33202 33963 -32898
rect 34267 -33202 34275 -32898
rect 8275 -33210 34275 -33202
rect 8615 -33238 8935 -33210
rect 8615 -33862 8623 -33238
rect 8927 -33862 8935 -33238
rect 8615 -33890 8935 -33862
rect 9615 -33238 9935 -33210
rect 9615 -33862 9623 -33238
rect 9927 -33862 9935 -33238
rect 9615 -33890 9935 -33862
rect 10615 -33238 10935 -33210
rect 10615 -33862 10623 -33238
rect 10927 -33862 10935 -33238
rect 10615 -33890 10935 -33862
rect 11615 -33238 11935 -33210
rect 11615 -33862 11623 -33238
rect 11927 -33862 11935 -33238
rect 11615 -33890 11935 -33862
rect 12615 -33238 12935 -33210
rect 12615 -33862 12623 -33238
rect 12927 -33862 12935 -33238
rect 12615 -33890 12935 -33862
rect 13615 -33238 13935 -33210
rect 13615 -33862 13623 -33238
rect 13927 -33862 13935 -33238
rect 13615 -33890 13935 -33862
rect 14615 -33238 14935 -33210
rect 14615 -33862 14623 -33238
rect 14927 -33862 14935 -33238
rect 14615 -33890 14935 -33862
rect 15615 -33238 15935 -33210
rect 15615 -33862 15623 -33238
rect 15927 -33862 15935 -33238
rect 15615 -33890 15935 -33862
rect 16615 -33238 16935 -33210
rect 16615 -33862 16623 -33238
rect 16927 -33862 16935 -33238
rect 16615 -33890 16935 -33862
rect 17615 -33238 17935 -33210
rect 17615 -33862 17623 -33238
rect 17927 -33862 17935 -33238
rect 17615 -33890 17935 -33862
rect 18615 -33238 18935 -33210
rect 18615 -33862 18623 -33238
rect 18927 -33862 18935 -33238
rect 18615 -33890 18935 -33862
rect 19615 -33238 19935 -33210
rect 19615 -33862 19623 -33238
rect 19927 -33862 19935 -33238
rect 19615 -33890 19935 -33862
rect 20615 -33238 20935 -33210
rect 20615 -33862 20623 -33238
rect 20927 -33862 20935 -33238
rect 20615 -33890 20935 -33862
rect 21615 -33238 21935 -33210
rect 21615 -33862 21623 -33238
rect 21927 -33862 21935 -33238
rect 21615 -33890 21935 -33862
rect 22615 -33238 22935 -33210
rect 22615 -33862 22623 -33238
rect 22927 -33862 22935 -33238
rect 22615 -33890 22935 -33862
rect 23615 -33238 23935 -33210
rect 23615 -33862 23623 -33238
rect 23927 -33862 23935 -33238
rect 23615 -33890 23935 -33862
rect 24615 -33238 24935 -33210
rect 24615 -33862 24623 -33238
rect 24927 -33862 24935 -33238
rect 24615 -33890 24935 -33862
rect 25615 -33238 25935 -33210
rect 25615 -33862 25623 -33238
rect 25927 -33862 25935 -33238
rect 25615 -33890 25935 -33862
rect 26615 -33238 26935 -33210
rect 26615 -33862 26623 -33238
rect 26927 -33862 26935 -33238
rect 26615 -33890 26935 -33862
rect 27615 -33238 27935 -33210
rect 27615 -33862 27623 -33238
rect 27927 -33862 27935 -33238
rect 27615 -33890 27935 -33862
rect 28615 -33238 28935 -33210
rect 28615 -33862 28623 -33238
rect 28927 -33862 28935 -33238
rect 28615 -33890 28935 -33862
rect 29615 -33238 29935 -33210
rect 29615 -33862 29623 -33238
rect 29927 -33862 29935 -33238
rect 29615 -33890 29935 -33862
rect 30615 -33238 30935 -33210
rect 30615 -33862 30623 -33238
rect 30927 -33862 30935 -33238
rect 30615 -33890 30935 -33862
rect 31615 -33238 31935 -33210
rect 31615 -33862 31623 -33238
rect 31927 -33862 31935 -33238
rect 31615 -33890 31935 -33862
rect 32615 -33238 32935 -33210
rect 32615 -33862 32623 -33238
rect 32927 -33862 32935 -33238
rect 32615 -33890 32935 -33862
rect 33615 -33238 33935 -33210
rect 33615 -33862 33623 -33238
rect 33927 -33862 33935 -33238
rect 33615 -33890 33935 -33862
rect 8275 -33898 34275 -33890
rect 8275 -34202 8283 -33898
rect 8587 -34202 8623 -33898
rect 8927 -34202 8963 -33898
rect 9587 -34202 9623 -33898
rect 9927 -34202 9963 -33898
rect 10587 -34202 10623 -33898
rect 10927 -34202 10963 -33898
rect 11587 -34202 11623 -33898
rect 11927 -34202 11963 -33898
rect 12587 -34202 12623 -33898
rect 12927 -34202 12963 -33898
rect 13587 -34202 13623 -33898
rect 13927 -34202 13963 -33898
rect 14587 -34202 14623 -33898
rect 14927 -34202 14963 -33898
rect 15587 -34202 15623 -33898
rect 15927 -34202 15963 -33898
rect 16587 -34202 16623 -33898
rect 16927 -34202 16963 -33898
rect 17587 -34202 17623 -33898
rect 17927 -34202 17963 -33898
rect 18587 -34202 18623 -33898
rect 18927 -34202 18963 -33898
rect 19587 -34202 19623 -33898
rect 19927 -34202 19963 -33898
rect 20587 -34202 20623 -33898
rect 20927 -34202 20963 -33898
rect 21587 -34202 21623 -33898
rect 21927 -34202 21963 -33898
rect 22587 -34202 22623 -33898
rect 22927 -34202 22963 -33898
rect 23587 -34202 23623 -33898
rect 23927 -34202 23963 -33898
rect 24587 -34202 24623 -33898
rect 24927 -34202 24963 -33898
rect 25587 -34202 25623 -33898
rect 25927 -34202 25963 -33898
rect 26587 -34202 26623 -33898
rect 26927 -34202 26963 -33898
rect 27587 -34202 27623 -33898
rect 27927 -34202 27963 -33898
rect 28587 -34202 28623 -33898
rect 28927 -34202 28963 -33898
rect 29587 -34202 29623 -33898
rect 29927 -34202 29963 -33898
rect 30587 -34202 30623 -33898
rect 30927 -34202 30963 -33898
rect 31587 -34202 31623 -33898
rect 31927 -34202 31963 -33898
rect 32587 -34202 32623 -33898
rect 32927 -34202 32963 -33898
rect 33587 -34202 33623 -33898
rect 33927 -34202 33963 -33898
rect 34267 -34202 34275 -33898
rect 8275 -34210 34275 -34202
rect 8615 -34238 8935 -34210
rect 8615 -34862 8623 -34238
rect 8927 -34862 8935 -34238
rect 8615 -34890 8935 -34862
rect 9615 -34238 9935 -34210
rect 9615 -34862 9623 -34238
rect 9927 -34862 9935 -34238
rect 9615 -34890 9935 -34862
rect 10615 -34238 10935 -34210
rect 10615 -34862 10623 -34238
rect 10927 -34862 10935 -34238
rect 10615 -34890 10935 -34862
rect 11615 -34238 11935 -34210
rect 11615 -34862 11623 -34238
rect 11927 -34862 11935 -34238
rect 11615 -34890 11935 -34862
rect 12615 -34238 12935 -34210
rect 12615 -34862 12623 -34238
rect 12927 -34862 12935 -34238
rect 12615 -34890 12935 -34862
rect 13615 -34238 13935 -34210
rect 13615 -34862 13623 -34238
rect 13927 -34862 13935 -34238
rect 13615 -34890 13935 -34862
rect 14615 -34238 14935 -34210
rect 14615 -34862 14623 -34238
rect 14927 -34862 14935 -34238
rect 14615 -34890 14935 -34862
rect 15615 -34238 15935 -34210
rect 15615 -34862 15623 -34238
rect 15927 -34862 15935 -34238
rect 15615 -34890 15935 -34862
rect 16615 -34238 16935 -34210
rect 16615 -34862 16623 -34238
rect 16927 -34862 16935 -34238
rect 16615 -34890 16935 -34862
rect 17615 -34238 17935 -34210
rect 17615 -34862 17623 -34238
rect 17927 -34862 17935 -34238
rect 17615 -34890 17935 -34862
rect 18615 -34238 18935 -34210
rect 18615 -34862 18623 -34238
rect 18927 -34862 18935 -34238
rect 18615 -34890 18935 -34862
rect 19615 -34238 19935 -34210
rect 19615 -34862 19623 -34238
rect 19927 -34862 19935 -34238
rect 19615 -34890 19935 -34862
rect 20615 -34238 20935 -34210
rect 20615 -34862 20623 -34238
rect 20927 -34862 20935 -34238
rect 20615 -34890 20935 -34862
rect 21615 -34238 21935 -34210
rect 21615 -34862 21623 -34238
rect 21927 -34862 21935 -34238
rect 21615 -34890 21935 -34862
rect 22615 -34238 22935 -34210
rect 22615 -34862 22623 -34238
rect 22927 -34862 22935 -34238
rect 22615 -34890 22935 -34862
rect 23615 -34238 23935 -34210
rect 23615 -34862 23623 -34238
rect 23927 -34862 23935 -34238
rect 23615 -34890 23935 -34862
rect 24615 -34238 24935 -34210
rect 24615 -34862 24623 -34238
rect 24927 -34862 24935 -34238
rect 24615 -34890 24935 -34862
rect 25615 -34238 25935 -34210
rect 25615 -34862 25623 -34238
rect 25927 -34862 25935 -34238
rect 25615 -34890 25935 -34862
rect 26615 -34238 26935 -34210
rect 26615 -34862 26623 -34238
rect 26927 -34862 26935 -34238
rect 26615 -34890 26935 -34862
rect 27615 -34238 27935 -34210
rect 27615 -34862 27623 -34238
rect 27927 -34862 27935 -34238
rect 27615 -34890 27935 -34862
rect 28615 -34238 28935 -34210
rect 28615 -34862 28623 -34238
rect 28927 -34862 28935 -34238
rect 28615 -34890 28935 -34862
rect 29615 -34238 29935 -34210
rect 29615 -34862 29623 -34238
rect 29927 -34862 29935 -34238
rect 29615 -34890 29935 -34862
rect 30615 -34238 30935 -34210
rect 30615 -34862 30623 -34238
rect 30927 -34862 30935 -34238
rect 30615 -34890 30935 -34862
rect 31615 -34238 31935 -34210
rect 31615 -34862 31623 -34238
rect 31927 -34862 31935 -34238
rect 31615 -34890 31935 -34862
rect 32615 -34238 32935 -34210
rect 32615 -34862 32623 -34238
rect 32927 -34862 32935 -34238
rect 32615 -34890 32935 -34862
rect 33615 -34238 33935 -34210
rect 33615 -34862 33623 -34238
rect 33927 -34862 33935 -34238
rect 33615 -34890 33935 -34862
rect 8275 -34898 34275 -34890
rect 8275 -35202 8283 -34898
rect 8587 -35202 8623 -34898
rect 8927 -35202 8963 -34898
rect 9587 -35202 9623 -34898
rect 9927 -35202 9963 -34898
rect 10587 -35202 10623 -34898
rect 10927 -35202 10963 -34898
rect 11587 -35202 11623 -34898
rect 11927 -35202 11963 -34898
rect 12587 -35202 12623 -34898
rect 12927 -35202 12963 -34898
rect 13587 -35202 13623 -34898
rect 13927 -35202 13963 -34898
rect 14587 -35202 14623 -34898
rect 14927 -35202 14963 -34898
rect 15587 -35202 15623 -34898
rect 15927 -35202 15963 -34898
rect 16587 -35202 16623 -34898
rect 16927 -35202 16963 -34898
rect 17587 -35202 17623 -34898
rect 17927 -35202 17963 -34898
rect 18587 -35202 18623 -34898
rect 18927 -35202 18963 -34898
rect 19587 -35202 19623 -34898
rect 19927 -35202 19963 -34898
rect 20587 -35202 20623 -34898
rect 20927 -35202 20963 -34898
rect 21587 -35202 21623 -34898
rect 21927 -35202 21963 -34898
rect 22587 -35202 22623 -34898
rect 22927 -35202 22963 -34898
rect 23587 -35202 23623 -34898
rect 23927 -35202 23963 -34898
rect 24587 -35202 24623 -34898
rect 24927 -35202 24963 -34898
rect 25587 -35202 25623 -34898
rect 25927 -35202 25963 -34898
rect 26587 -35202 26623 -34898
rect 26927 -35202 26963 -34898
rect 27587 -35202 27623 -34898
rect 27927 -35202 27963 -34898
rect 28587 -35202 28623 -34898
rect 28927 -35202 28963 -34898
rect 29587 -35202 29623 -34898
rect 29927 -35202 29963 -34898
rect 30587 -35202 30623 -34898
rect 30927 -35202 30963 -34898
rect 31587 -35202 31623 -34898
rect 31927 -35202 31963 -34898
rect 32587 -35202 32623 -34898
rect 32927 -35202 32963 -34898
rect 33587 -35202 33623 -34898
rect 33927 -35202 33963 -34898
rect 34267 -35202 34275 -34898
rect 8275 -35210 34275 -35202
rect 8615 -35238 8935 -35210
rect 8615 -35862 8623 -35238
rect 8927 -35862 8935 -35238
rect 8615 -35890 8935 -35862
rect 9615 -35238 9935 -35210
rect 9615 -35862 9623 -35238
rect 9927 -35862 9935 -35238
rect 9615 -35890 9935 -35862
rect 10615 -35238 10935 -35210
rect 10615 -35862 10623 -35238
rect 10927 -35862 10935 -35238
rect 10615 -35890 10935 -35862
rect 11615 -35238 11935 -35210
rect 11615 -35862 11623 -35238
rect 11927 -35862 11935 -35238
rect 11615 -35890 11935 -35862
rect 12615 -35238 12935 -35210
rect 12615 -35862 12623 -35238
rect 12927 -35862 12935 -35238
rect 12615 -35890 12935 -35862
rect 13615 -35238 13935 -35210
rect 13615 -35862 13623 -35238
rect 13927 -35862 13935 -35238
rect 13615 -35890 13935 -35862
rect 14615 -35238 14935 -35210
rect 14615 -35862 14623 -35238
rect 14927 -35862 14935 -35238
rect 14615 -35890 14935 -35862
rect 15615 -35238 15935 -35210
rect 15615 -35862 15623 -35238
rect 15927 -35862 15935 -35238
rect 15615 -35890 15935 -35862
rect 16615 -35238 16935 -35210
rect 16615 -35862 16623 -35238
rect 16927 -35862 16935 -35238
rect 16615 -35890 16935 -35862
rect 17615 -35238 17935 -35210
rect 17615 -35862 17623 -35238
rect 17927 -35862 17935 -35238
rect 17615 -35890 17935 -35862
rect 18615 -35238 18935 -35210
rect 18615 -35862 18623 -35238
rect 18927 -35862 18935 -35238
rect 18615 -35890 18935 -35862
rect 19615 -35238 19935 -35210
rect 19615 -35862 19623 -35238
rect 19927 -35862 19935 -35238
rect 19615 -35890 19935 -35862
rect 20615 -35238 20935 -35210
rect 20615 -35862 20623 -35238
rect 20927 -35862 20935 -35238
rect 20615 -35890 20935 -35862
rect 21615 -35238 21935 -35210
rect 21615 -35862 21623 -35238
rect 21927 -35862 21935 -35238
rect 21615 -35890 21935 -35862
rect 22615 -35238 22935 -35210
rect 22615 -35862 22623 -35238
rect 22927 -35862 22935 -35238
rect 22615 -35890 22935 -35862
rect 23615 -35238 23935 -35210
rect 23615 -35862 23623 -35238
rect 23927 -35862 23935 -35238
rect 23615 -35890 23935 -35862
rect 24615 -35238 24935 -35210
rect 24615 -35862 24623 -35238
rect 24927 -35862 24935 -35238
rect 24615 -35890 24935 -35862
rect 25615 -35238 25935 -35210
rect 25615 -35862 25623 -35238
rect 25927 -35862 25935 -35238
rect 25615 -35890 25935 -35862
rect 26615 -35238 26935 -35210
rect 26615 -35862 26623 -35238
rect 26927 -35862 26935 -35238
rect 26615 -35890 26935 -35862
rect 27615 -35238 27935 -35210
rect 27615 -35862 27623 -35238
rect 27927 -35862 27935 -35238
rect 27615 -35890 27935 -35862
rect 28615 -35238 28935 -35210
rect 28615 -35862 28623 -35238
rect 28927 -35862 28935 -35238
rect 28615 -35890 28935 -35862
rect 29615 -35238 29935 -35210
rect 29615 -35862 29623 -35238
rect 29927 -35862 29935 -35238
rect 29615 -35890 29935 -35862
rect 30615 -35238 30935 -35210
rect 30615 -35862 30623 -35238
rect 30927 -35862 30935 -35238
rect 30615 -35890 30935 -35862
rect 31615 -35238 31935 -35210
rect 31615 -35862 31623 -35238
rect 31927 -35862 31935 -35238
rect 31615 -35890 31935 -35862
rect 32615 -35238 32935 -35210
rect 32615 -35862 32623 -35238
rect 32927 -35862 32935 -35238
rect 32615 -35890 32935 -35862
rect 33615 -35238 33935 -35210
rect 33615 -35862 33623 -35238
rect 33927 -35862 33935 -35238
rect 33615 -35890 33935 -35862
rect 8275 -35898 34275 -35890
rect 8275 -36202 8283 -35898
rect 8587 -36202 8623 -35898
rect 8927 -36202 8963 -35898
rect 9587 -36202 9623 -35898
rect 9927 -36202 9963 -35898
rect 10587 -36202 10623 -35898
rect 10927 -36202 10963 -35898
rect 11587 -36202 11623 -35898
rect 11927 -36202 11963 -35898
rect 12587 -36202 12623 -35898
rect 12927 -36202 12963 -35898
rect 13587 -36202 13623 -35898
rect 13927 -36202 13963 -35898
rect 14587 -36202 14623 -35898
rect 14927 -36202 14963 -35898
rect 15587 -36202 15623 -35898
rect 15927 -36202 15963 -35898
rect 16587 -36202 16623 -35898
rect 16927 -36202 16963 -35898
rect 17587 -36202 17623 -35898
rect 17927 -36202 17963 -35898
rect 18587 -36202 18623 -35898
rect 18927 -36202 18963 -35898
rect 19587 -36202 19623 -35898
rect 19927 -36202 19963 -35898
rect 20587 -36202 20623 -35898
rect 20927 -36202 20963 -35898
rect 21587 -36202 21623 -35898
rect 21927 -36202 21963 -35898
rect 22587 -36202 22623 -35898
rect 22927 -36202 22963 -35898
rect 23587 -36202 23623 -35898
rect 23927 -36202 23963 -35898
rect 24587 -36202 24623 -35898
rect 24927 -36202 24963 -35898
rect 25587 -36202 25623 -35898
rect 25927 -36202 25963 -35898
rect 26587 -36202 26623 -35898
rect 26927 -36202 26963 -35898
rect 27587 -36202 27623 -35898
rect 27927 -36202 27963 -35898
rect 28587 -36202 28623 -35898
rect 28927 -36202 28963 -35898
rect 29587 -36202 29623 -35898
rect 29927 -36202 29963 -35898
rect 30587 -36202 30623 -35898
rect 30927 -36202 30963 -35898
rect 31587 -36202 31623 -35898
rect 31927 -36202 31963 -35898
rect 32587 -36202 32623 -35898
rect 32927 -36202 32963 -35898
rect 33587 -36202 33623 -35898
rect 33927 -36202 33963 -35898
rect 34267 -36202 34275 -35898
rect 8275 -36210 34275 -36202
rect 8615 -36238 8935 -36210
rect 8615 -36862 8623 -36238
rect 8927 -36862 8935 -36238
rect 8615 -36890 8935 -36862
rect 9615 -36238 9935 -36210
rect 9615 -36862 9623 -36238
rect 9927 -36862 9935 -36238
rect 9615 -36890 9935 -36862
rect 10615 -36238 10935 -36210
rect 10615 -36862 10623 -36238
rect 10927 -36862 10935 -36238
rect 10615 -36890 10935 -36862
rect 11615 -36238 11935 -36210
rect 11615 -36862 11623 -36238
rect 11927 -36862 11935 -36238
rect 11615 -36890 11935 -36862
rect 12615 -36238 12935 -36210
rect 12615 -36862 12623 -36238
rect 12927 -36862 12935 -36238
rect 12615 -36890 12935 -36862
rect 13615 -36238 13935 -36210
rect 13615 -36862 13623 -36238
rect 13927 -36862 13935 -36238
rect 13615 -36890 13935 -36862
rect 14615 -36238 14935 -36210
rect 14615 -36862 14623 -36238
rect 14927 -36862 14935 -36238
rect 14615 -36890 14935 -36862
rect 15615 -36238 15935 -36210
rect 15615 -36862 15623 -36238
rect 15927 -36862 15935 -36238
rect 15615 -36890 15935 -36862
rect 16615 -36238 16935 -36210
rect 16615 -36862 16623 -36238
rect 16927 -36862 16935 -36238
rect 16615 -36890 16935 -36862
rect 17615 -36238 17935 -36210
rect 17615 -36862 17623 -36238
rect 17927 -36862 17935 -36238
rect 17615 -36890 17935 -36862
rect 18615 -36238 18935 -36210
rect 18615 -36862 18623 -36238
rect 18927 -36862 18935 -36238
rect 18615 -36890 18935 -36862
rect 19615 -36238 19935 -36210
rect 19615 -36862 19623 -36238
rect 19927 -36862 19935 -36238
rect 19615 -36890 19935 -36862
rect 20615 -36238 20935 -36210
rect 20615 -36862 20623 -36238
rect 20927 -36862 20935 -36238
rect 20615 -36890 20935 -36862
rect 21615 -36238 21935 -36210
rect 21615 -36862 21623 -36238
rect 21927 -36862 21935 -36238
rect 21615 -36890 21935 -36862
rect 22615 -36238 22935 -36210
rect 22615 -36862 22623 -36238
rect 22927 -36862 22935 -36238
rect 22615 -36890 22935 -36862
rect 23615 -36238 23935 -36210
rect 23615 -36862 23623 -36238
rect 23927 -36862 23935 -36238
rect 23615 -36890 23935 -36862
rect 24615 -36238 24935 -36210
rect 24615 -36862 24623 -36238
rect 24927 -36862 24935 -36238
rect 24615 -36890 24935 -36862
rect 25615 -36238 25935 -36210
rect 25615 -36862 25623 -36238
rect 25927 -36862 25935 -36238
rect 25615 -36890 25935 -36862
rect 26615 -36238 26935 -36210
rect 26615 -36862 26623 -36238
rect 26927 -36862 26935 -36238
rect 26615 -36890 26935 -36862
rect 27615 -36238 27935 -36210
rect 27615 -36862 27623 -36238
rect 27927 -36862 27935 -36238
rect 27615 -36890 27935 -36862
rect 28615 -36238 28935 -36210
rect 28615 -36862 28623 -36238
rect 28927 -36862 28935 -36238
rect 28615 -36890 28935 -36862
rect 29615 -36238 29935 -36210
rect 29615 -36862 29623 -36238
rect 29927 -36862 29935 -36238
rect 29615 -36890 29935 -36862
rect 30615 -36238 30935 -36210
rect 30615 -36862 30623 -36238
rect 30927 -36862 30935 -36238
rect 30615 -36890 30935 -36862
rect 31615 -36238 31935 -36210
rect 31615 -36862 31623 -36238
rect 31927 -36862 31935 -36238
rect 31615 -36890 31935 -36862
rect 32615 -36238 32935 -36210
rect 32615 -36862 32623 -36238
rect 32927 -36862 32935 -36238
rect 32615 -36890 32935 -36862
rect 33615 -36238 33935 -36210
rect 33615 -36862 33623 -36238
rect 33927 -36862 33935 -36238
rect 33615 -36890 33935 -36862
rect 8275 -36898 34275 -36890
rect 8275 -37202 8283 -36898
rect 8587 -37202 8623 -36898
rect 8927 -37202 8963 -36898
rect 9587 -37202 9623 -36898
rect 9927 -37202 9963 -36898
rect 10587 -37202 10623 -36898
rect 10927 -37202 10963 -36898
rect 11587 -37202 11623 -36898
rect 11927 -37202 11963 -36898
rect 12587 -37202 12623 -36898
rect 12927 -37202 12963 -36898
rect 13587 -37202 13623 -36898
rect 13927 -37202 13963 -36898
rect 14587 -37202 14623 -36898
rect 14927 -37202 14963 -36898
rect 15587 -37202 15623 -36898
rect 15927 -37202 15963 -36898
rect 16587 -37202 16623 -36898
rect 16927 -37202 16963 -36898
rect 17587 -37202 17623 -36898
rect 17927 -37202 17963 -36898
rect 18587 -37202 18623 -36898
rect 18927 -37202 18963 -36898
rect 19587 -37202 19623 -36898
rect 19927 -37202 19963 -36898
rect 20587 -37202 20623 -36898
rect 20927 -37202 20963 -36898
rect 21587 -37202 21623 -36898
rect 21927 -37202 21963 -36898
rect 22587 -37202 22623 -36898
rect 22927 -37202 22963 -36898
rect 23587 -37202 23623 -36898
rect 23927 -37202 23963 -36898
rect 24587 -37202 24623 -36898
rect 24927 -37202 24963 -36898
rect 25587 -37202 25623 -36898
rect 25927 -37202 25963 -36898
rect 26587 -37202 26623 -36898
rect 26927 -37202 26963 -36898
rect 27587 -37202 27623 -36898
rect 27927 -37202 27963 -36898
rect 28587 -37202 28623 -36898
rect 28927 -37202 28963 -36898
rect 29587 -37202 29623 -36898
rect 29927 -37202 29963 -36898
rect 30587 -37202 30623 -36898
rect 30927 -37202 30963 -36898
rect 31587 -37202 31623 -36898
rect 31927 -37202 31963 -36898
rect 32587 -37202 32623 -36898
rect 32927 -37202 32963 -36898
rect 33587 -37202 33623 -36898
rect 33927 -37202 33963 -36898
rect 34267 -37202 34275 -36898
rect 8275 -37210 34275 -37202
rect 8615 -37238 8935 -37210
rect 8615 -37862 8623 -37238
rect 8927 -37862 8935 -37238
rect 8615 -37890 8935 -37862
rect 9615 -37238 9935 -37210
rect 9615 -37862 9623 -37238
rect 9927 -37862 9935 -37238
rect 9615 -37890 9935 -37862
rect 10615 -37238 10935 -37210
rect 10615 -37862 10623 -37238
rect 10927 -37862 10935 -37238
rect 10615 -37890 10935 -37862
rect 11615 -37238 11935 -37210
rect 11615 -37862 11623 -37238
rect 11927 -37862 11935 -37238
rect 11615 -37890 11935 -37862
rect 12615 -37238 12935 -37210
rect 12615 -37862 12623 -37238
rect 12927 -37862 12935 -37238
rect 12615 -37890 12935 -37862
rect 13615 -37238 13935 -37210
rect 13615 -37862 13623 -37238
rect 13927 -37862 13935 -37238
rect 13615 -37890 13935 -37862
rect 14615 -37238 14935 -37210
rect 14615 -37862 14623 -37238
rect 14927 -37862 14935 -37238
rect 14615 -37890 14935 -37862
rect 15615 -37238 15935 -37210
rect 15615 -37862 15623 -37238
rect 15927 -37862 15935 -37238
rect 15615 -37890 15935 -37862
rect 16615 -37238 16935 -37210
rect 16615 -37862 16623 -37238
rect 16927 -37862 16935 -37238
rect 16615 -37890 16935 -37862
rect 17615 -37238 17935 -37210
rect 17615 -37862 17623 -37238
rect 17927 -37862 17935 -37238
rect 17615 -37890 17935 -37862
rect 18615 -37238 18935 -37210
rect 18615 -37862 18623 -37238
rect 18927 -37862 18935 -37238
rect 18615 -37890 18935 -37862
rect 19615 -37238 19935 -37210
rect 19615 -37862 19623 -37238
rect 19927 -37862 19935 -37238
rect 19615 -37890 19935 -37862
rect 20615 -37238 20935 -37210
rect 20615 -37862 20623 -37238
rect 20927 -37862 20935 -37238
rect 20615 -37890 20935 -37862
rect 21615 -37238 21935 -37210
rect 21615 -37862 21623 -37238
rect 21927 -37862 21935 -37238
rect 21615 -37890 21935 -37862
rect 22615 -37238 22935 -37210
rect 22615 -37862 22623 -37238
rect 22927 -37862 22935 -37238
rect 22615 -37890 22935 -37862
rect 23615 -37238 23935 -37210
rect 23615 -37862 23623 -37238
rect 23927 -37862 23935 -37238
rect 23615 -37890 23935 -37862
rect 24615 -37238 24935 -37210
rect 24615 -37862 24623 -37238
rect 24927 -37862 24935 -37238
rect 24615 -37890 24935 -37862
rect 25615 -37238 25935 -37210
rect 25615 -37862 25623 -37238
rect 25927 -37862 25935 -37238
rect 25615 -37890 25935 -37862
rect 26615 -37238 26935 -37210
rect 26615 -37862 26623 -37238
rect 26927 -37862 26935 -37238
rect 26615 -37890 26935 -37862
rect 27615 -37238 27935 -37210
rect 27615 -37862 27623 -37238
rect 27927 -37862 27935 -37238
rect 27615 -37890 27935 -37862
rect 28615 -37238 28935 -37210
rect 28615 -37862 28623 -37238
rect 28927 -37862 28935 -37238
rect 28615 -37890 28935 -37862
rect 29615 -37238 29935 -37210
rect 29615 -37862 29623 -37238
rect 29927 -37862 29935 -37238
rect 29615 -37890 29935 -37862
rect 30615 -37238 30935 -37210
rect 30615 -37862 30623 -37238
rect 30927 -37862 30935 -37238
rect 30615 -37890 30935 -37862
rect 31615 -37238 31935 -37210
rect 31615 -37862 31623 -37238
rect 31927 -37862 31935 -37238
rect 31615 -37890 31935 -37862
rect 32615 -37238 32935 -37210
rect 32615 -37862 32623 -37238
rect 32927 -37862 32935 -37238
rect 32615 -37890 32935 -37862
rect 33615 -37238 33935 -37210
rect 33615 -37862 33623 -37238
rect 33927 -37862 33935 -37238
rect 33615 -37890 33935 -37862
rect 8275 -37898 34275 -37890
rect 8275 -38202 8283 -37898
rect 8587 -38202 8623 -37898
rect 8927 -38202 8963 -37898
rect 9587 -38202 9623 -37898
rect 9927 -38202 9963 -37898
rect 10587 -38202 10623 -37898
rect 10927 -38202 10963 -37898
rect 11587 -38202 11623 -37898
rect 11927 -38202 11963 -37898
rect 12587 -38202 12623 -37898
rect 12927 -38202 12963 -37898
rect 13587 -38202 13623 -37898
rect 13927 -38202 13963 -37898
rect 14587 -38202 14623 -37898
rect 14927 -38202 14963 -37898
rect 15587 -38202 15623 -37898
rect 15927 -38202 15963 -37898
rect 16587 -38202 16623 -37898
rect 16927 -38202 16963 -37898
rect 17587 -38202 17623 -37898
rect 17927 -38202 17963 -37898
rect 18587 -38202 18623 -37898
rect 18927 -38202 18963 -37898
rect 19587 -38202 19623 -37898
rect 19927 -38202 19963 -37898
rect 20587 -38202 20623 -37898
rect 20927 -38202 20963 -37898
rect 21587 -38202 21623 -37898
rect 21927 -38202 21963 -37898
rect 22587 -38202 22623 -37898
rect 22927 -38202 22963 -37898
rect 23587 -38202 23623 -37898
rect 23927 -38202 23963 -37898
rect 24587 -38202 24623 -37898
rect 24927 -38202 24963 -37898
rect 25587 -38202 25623 -37898
rect 25927 -38202 25963 -37898
rect 26587 -38202 26623 -37898
rect 26927 -38202 26963 -37898
rect 27587 -38202 27623 -37898
rect 27927 -38202 27963 -37898
rect 28587 -38202 28623 -37898
rect 28927 -38202 28963 -37898
rect 29587 -38202 29623 -37898
rect 29927 -38202 29963 -37898
rect 30587 -38202 30623 -37898
rect 30927 -38202 30963 -37898
rect 31587 -38202 31623 -37898
rect 31927 -38202 31963 -37898
rect 32587 -38202 32623 -37898
rect 32927 -38202 32963 -37898
rect 33587 -38202 33623 -37898
rect 33927 -38202 33963 -37898
rect 34267 -38202 34275 -37898
rect 8275 -38210 34275 -38202
rect 8615 -38238 8935 -38210
rect 8615 -38862 8623 -38238
rect 8927 -38862 8935 -38238
rect 8615 -38890 8935 -38862
rect 9615 -38238 9935 -38210
rect 9615 -38862 9623 -38238
rect 9927 -38862 9935 -38238
rect 9615 -38890 9935 -38862
rect 10615 -38238 10935 -38210
rect 10615 -38862 10623 -38238
rect 10927 -38862 10935 -38238
rect 10615 -38890 10935 -38862
rect 11615 -38238 11935 -38210
rect 11615 -38862 11623 -38238
rect 11927 -38862 11935 -38238
rect 11615 -38890 11935 -38862
rect 12615 -38238 12935 -38210
rect 12615 -38862 12623 -38238
rect 12927 -38862 12935 -38238
rect 12615 -38890 12935 -38862
rect 13615 -38238 13935 -38210
rect 13615 -38862 13623 -38238
rect 13927 -38862 13935 -38238
rect 13615 -38890 13935 -38862
rect 14615 -38238 14935 -38210
rect 14615 -38862 14623 -38238
rect 14927 -38862 14935 -38238
rect 14615 -38890 14935 -38862
rect 15615 -38238 15935 -38210
rect 15615 -38862 15623 -38238
rect 15927 -38862 15935 -38238
rect 15615 -38890 15935 -38862
rect 16615 -38238 16935 -38210
rect 16615 -38862 16623 -38238
rect 16927 -38862 16935 -38238
rect 16615 -38890 16935 -38862
rect 17615 -38238 17935 -38210
rect 17615 -38862 17623 -38238
rect 17927 -38862 17935 -38238
rect 17615 -38890 17935 -38862
rect 18615 -38238 18935 -38210
rect 18615 -38862 18623 -38238
rect 18927 -38862 18935 -38238
rect 18615 -38890 18935 -38862
rect 19615 -38238 19935 -38210
rect 19615 -38862 19623 -38238
rect 19927 -38862 19935 -38238
rect 19615 -38890 19935 -38862
rect 20615 -38238 20935 -38210
rect 20615 -38862 20623 -38238
rect 20927 -38862 20935 -38238
rect 20615 -38890 20935 -38862
rect 21615 -38238 21935 -38210
rect 21615 -38862 21623 -38238
rect 21927 -38862 21935 -38238
rect 21615 -38890 21935 -38862
rect 22615 -38238 22935 -38210
rect 22615 -38862 22623 -38238
rect 22927 -38862 22935 -38238
rect 22615 -38890 22935 -38862
rect 23615 -38238 23935 -38210
rect 23615 -38862 23623 -38238
rect 23927 -38862 23935 -38238
rect 23615 -38890 23935 -38862
rect 24615 -38238 24935 -38210
rect 24615 -38862 24623 -38238
rect 24927 -38862 24935 -38238
rect 24615 -38890 24935 -38862
rect 25615 -38238 25935 -38210
rect 25615 -38862 25623 -38238
rect 25927 -38862 25935 -38238
rect 25615 -38890 25935 -38862
rect 26615 -38238 26935 -38210
rect 26615 -38862 26623 -38238
rect 26927 -38862 26935 -38238
rect 26615 -38890 26935 -38862
rect 27615 -38238 27935 -38210
rect 27615 -38862 27623 -38238
rect 27927 -38862 27935 -38238
rect 27615 -38890 27935 -38862
rect 28615 -38238 28935 -38210
rect 28615 -38862 28623 -38238
rect 28927 -38862 28935 -38238
rect 28615 -38890 28935 -38862
rect 29615 -38238 29935 -38210
rect 29615 -38862 29623 -38238
rect 29927 -38862 29935 -38238
rect 29615 -38890 29935 -38862
rect 30615 -38238 30935 -38210
rect 30615 -38862 30623 -38238
rect 30927 -38862 30935 -38238
rect 30615 -38890 30935 -38862
rect 31615 -38238 31935 -38210
rect 31615 -38862 31623 -38238
rect 31927 -38862 31935 -38238
rect 31615 -38890 31935 -38862
rect 32615 -38238 32935 -38210
rect 32615 -38862 32623 -38238
rect 32927 -38862 32935 -38238
rect 32615 -38890 32935 -38862
rect 33615 -38238 33935 -38210
rect 33615 -38862 33623 -38238
rect 33927 -38862 33935 -38238
rect 33615 -38890 33935 -38862
rect 8275 -38898 34275 -38890
rect 8275 -39202 8283 -38898
rect 8587 -39202 8623 -38898
rect 8927 -39202 8963 -38898
rect 9587 -39202 9623 -38898
rect 9927 -39202 9963 -38898
rect 10587 -39202 10623 -38898
rect 10927 -39202 10963 -38898
rect 11587 -39202 11623 -38898
rect 11927 -39202 11963 -38898
rect 12587 -39202 12623 -38898
rect 12927 -39202 12963 -38898
rect 13587 -39202 13623 -38898
rect 13927 -39202 13963 -38898
rect 14587 -39202 14623 -38898
rect 14927 -39202 14963 -38898
rect 15587 -39202 15623 -38898
rect 15927 -39202 15963 -38898
rect 16587 -39202 16623 -38898
rect 16927 -39202 16963 -38898
rect 17587 -39202 17623 -38898
rect 17927 -39202 17963 -38898
rect 18587 -39202 18623 -38898
rect 18927 -39202 18963 -38898
rect 19587 -39202 19623 -38898
rect 19927 -39202 19963 -38898
rect 20587 -39202 20623 -38898
rect 20927 -39202 20963 -38898
rect 21587 -39202 21623 -38898
rect 21927 -39202 21963 -38898
rect 22587 -39202 22623 -38898
rect 22927 -39202 22963 -38898
rect 23587 -39202 23623 -38898
rect 23927 -39202 23963 -38898
rect 24587 -39202 24623 -38898
rect 24927 -39202 24963 -38898
rect 25587 -39202 25623 -38898
rect 25927 -39202 25963 -38898
rect 26587 -39202 26623 -38898
rect 26927 -39202 26963 -38898
rect 27587 -39202 27623 -38898
rect 27927 -39202 27963 -38898
rect 28587 -39202 28623 -38898
rect 28927 -39202 28963 -38898
rect 29587 -39202 29623 -38898
rect 29927 -39202 29963 -38898
rect 30587 -39202 30623 -38898
rect 30927 -39202 30963 -38898
rect 31587 -39202 31623 -38898
rect 31927 -39202 31963 -38898
rect 32587 -39202 32623 -38898
rect 32927 -39202 32963 -38898
rect 33587 -39202 33623 -38898
rect 33927 -39202 33963 -38898
rect 34267 -39202 34275 -38898
rect 8275 -39210 34275 -39202
rect 8615 -39238 8935 -39210
rect 8615 -39862 8623 -39238
rect 8927 -39862 8935 -39238
rect 8615 -39890 8935 -39862
rect 9615 -39238 9935 -39210
rect 9615 -39862 9623 -39238
rect 9927 -39862 9935 -39238
rect 9615 -39890 9935 -39862
rect 10615 -39238 10935 -39210
rect 10615 -39862 10623 -39238
rect 10927 -39862 10935 -39238
rect 10615 -39890 10935 -39862
rect 11615 -39238 11935 -39210
rect 11615 -39862 11623 -39238
rect 11927 -39862 11935 -39238
rect 11615 -39890 11935 -39862
rect 12615 -39238 12935 -39210
rect 12615 -39862 12623 -39238
rect 12927 -39862 12935 -39238
rect 12615 -39890 12935 -39862
rect 13615 -39238 13935 -39210
rect 13615 -39862 13623 -39238
rect 13927 -39862 13935 -39238
rect 13615 -39890 13935 -39862
rect 14615 -39238 14935 -39210
rect 14615 -39862 14623 -39238
rect 14927 -39862 14935 -39238
rect 14615 -39890 14935 -39862
rect 15615 -39238 15935 -39210
rect 15615 -39862 15623 -39238
rect 15927 -39862 15935 -39238
rect 15615 -39890 15935 -39862
rect 16615 -39238 16935 -39210
rect 16615 -39862 16623 -39238
rect 16927 -39862 16935 -39238
rect 16615 -39890 16935 -39862
rect 17615 -39238 17935 -39210
rect 17615 -39862 17623 -39238
rect 17927 -39862 17935 -39238
rect 17615 -39890 17935 -39862
rect 18615 -39238 18935 -39210
rect 18615 -39862 18623 -39238
rect 18927 -39862 18935 -39238
rect 18615 -39890 18935 -39862
rect 19615 -39238 19935 -39210
rect 19615 -39862 19623 -39238
rect 19927 -39862 19935 -39238
rect 19615 -39890 19935 -39862
rect 20615 -39238 20935 -39210
rect 20615 -39862 20623 -39238
rect 20927 -39862 20935 -39238
rect 20615 -39890 20935 -39862
rect 21615 -39238 21935 -39210
rect 21615 -39862 21623 -39238
rect 21927 -39862 21935 -39238
rect 21615 -39890 21935 -39862
rect 22615 -39238 22935 -39210
rect 22615 -39862 22623 -39238
rect 22927 -39862 22935 -39238
rect 22615 -39890 22935 -39862
rect 23615 -39238 23935 -39210
rect 23615 -39862 23623 -39238
rect 23927 -39862 23935 -39238
rect 23615 -39890 23935 -39862
rect 24615 -39238 24935 -39210
rect 24615 -39862 24623 -39238
rect 24927 -39862 24935 -39238
rect 24615 -39890 24935 -39862
rect 25615 -39238 25935 -39210
rect 25615 -39862 25623 -39238
rect 25927 -39862 25935 -39238
rect 25615 -39890 25935 -39862
rect 26615 -39238 26935 -39210
rect 26615 -39862 26623 -39238
rect 26927 -39862 26935 -39238
rect 26615 -39890 26935 -39862
rect 27615 -39238 27935 -39210
rect 27615 -39862 27623 -39238
rect 27927 -39862 27935 -39238
rect 27615 -39890 27935 -39862
rect 28615 -39238 28935 -39210
rect 28615 -39862 28623 -39238
rect 28927 -39862 28935 -39238
rect 28615 -39890 28935 -39862
rect 29615 -39238 29935 -39210
rect 29615 -39862 29623 -39238
rect 29927 -39862 29935 -39238
rect 29615 -39890 29935 -39862
rect 30615 -39238 30935 -39210
rect 30615 -39862 30623 -39238
rect 30927 -39862 30935 -39238
rect 30615 -39890 30935 -39862
rect 31615 -39238 31935 -39210
rect 31615 -39862 31623 -39238
rect 31927 -39862 31935 -39238
rect 31615 -39890 31935 -39862
rect 32615 -39238 32935 -39210
rect 32615 -39862 32623 -39238
rect 32927 -39862 32935 -39238
rect 32615 -39890 32935 -39862
rect 33615 -39238 33935 -39210
rect 33615 -39862 33623 -39238
rect 33927 -39862 33935 -39238
rect 33615 -39890 33935 -39862
rect 8275 -39898 34275 -39890
rect 8275 -40202 8283 -39898
rect 8587 -40202 8623 -39898
rect 8927 -40202 8963 -39898
rect 9587 -40202 9623 -39898
rect 9927 -40202 9963 -39898
rect 10587 -40202 10623 -39898
rect 10927 -40202 10963 -39898
rect 11587 -40202 11623 -39898
rect 11927 -40202 11963 -39898
rect 12587 -40202 12623 -39898
rect 12927 -40202 12963 -39898
rect 13587 -40202 13623 -39898
rect 13927 -40202 13963 -39898
rect 14587 -40202 14623 -39898
rect 14927 -40202 14963 -39898
rect 15587 -40202 15623 -39898
rect 15927 -40202 15963 -39898
rect 16587 -40202 16623 -39898
rect 16927 -40202 16963 -39898
rect 17587 -40202 17623 -39898
rect 17927 -40202 17963 -39898
rect 18587 -40202 18623 -39898
rect 18927 -40202 18963 -39898
rect 19587 -40202 19623 -39898
rect 19927 -40202 19963 -39898
rect 20587 -40202 20623 -39898
rect 20927 -40202 20963 -39898
rect 21587 -40202 21623 -39898
rect 21927 -40202 21963 -39898
rect 22587 -40202 22623 -39898
rect 22927 -40202 22963 -39898
rect 23587 -40202 23623 -39898
rect 23927 -40202 23963 -39898
rect 24587 -40202 24623 -39898
rect 24927 -40202 24963 -39898
rect 25587 -40202 25623 -39898
rect 25927 -40202 25963 -39898
rect 26587 -40202 26623 -39898
rect 26927 -40202 26963 -39898
rect 27587 -40202 27623 -39898
rect 27927 -40202 27963 -39898
rect 28587 -40202 28623 -39898
rect 28927 -40202 28963 -39898
rect 29587 -40202 29623 -39898
rect 29927 -40202 29963 -39898
rect 30587 -40202 30623 -39898
rect 30927 -40202 30963 -39898
rect 31587 -40202 31623 -39898
rect 31927 -40202 31963 -39898
rect 32587 -40202 32623 -39898
rect 32927 -40202 32963 -39898
rect 33587 -40202 33623 -39898
rect 33927 -40202 33963 -39898
rect 34267 -40202 34275 -39898
rect 8275 -40210 34275 -40202
rect 8615 -40238 8935 -40210
rect 8615 -40862 8623 -40238
rect 8927 -40862 8935 -40238
rect 8615 -40890 8935 -40862
rect 9615 -40238 9935 -40210
rect 9615 -40862 9623 -40238
rect 9927 -40862 9935 -40238
rect 9615 -40890 9935 -40862
rect 10615 -40238 10935 -40210
rect 10615 -40862 10623 -40238
rect 10927 -40862 10935 -40238
rect 10615 -40890 10935 -40862
rect 11615 -40238 11935 -40210
rect 11615 -40862 11623 -40238
rect 11927 -40862 11935 -40238
rect 11615 -40890 11935 -40862
rect 12615 -40238 12935 -40210
rect 12615 -40862 12623 -40238
rect 12927 -40862 12935 -40238
rect 12615 -40890 12935 -40862
rect 13615 -40238 13935 -40210
rect 13615 -40862 13623 -40238
rect 13927 -40862 13935 -40238
rect 13615 -40890 13935 -40862
rect 14615 -40238 14935 -40210
rect 14615 -40862 14623 -40238
rect 14927 -40862 14935 -40238
rect 14615 -40890 14935 -40862
rect 15615 -40238 15935 -40210
rect 15615 -40862 15623 -40238
rect 15927 -40862 15935 -40238
rect 15615 -40890 15935 -40862
rect 16615 -40238 16935 -40210
rect 16615 -40862 16623 -40238
rect 16927 -40862 16935 -40238
rect 16615 -40890 16935 -40862
rect 17615 -40238 17935 -40210
rect 17615 -40862 17623 -40238
rect 17927 -40862 17935 -40238
rect 17615 -40890 17935 -40862
rect 18615 -40238 18935 -40210
rect 18615 -40862 18623 -40238
rect 18927 -40862 18935 -40238
rect 18615 -40890 18935 -40862
rect 19615 -40238 19935 -40210
rect 19615 -40862 19623 -40238
rect 19927 -40862 19935 -40238
rect 19615 -40890 19935 -40862
rect 20615 -40238 20935 -40210
rect 20615 -40862 20623 -40238
rect 20927 -40862 20935 -40238
rect 20615 -40890 20935 -40862
rect 21615 -40238 21935 -40210
rect 21615 -40862 21623 -40238
rect 21927 -40862 21935 -40238
rect 21615 -40890 21935 -40862
rect 22615 -40238 22935 -40210
rect 22615 -40862 22623 -40238
rect 22927 -40862 22935 -40238
rect 22615 -40890 22935 -40862
rect 23615 -40238 23935 -40210
rect 23615 -40862 23623 -40238
rect 23927 -40862 23935 -40238
rect 23615 -40890 23935 -40862
rect 24615 -40238 24935 -40210
rect 24615 -40862 24623 -40238
rect 24927 -40862 24935 -40238
rect 24615 -40890 24935 -40862
rect 25615 -40238 25935 -40210
rect 25615 -40862 25623 -40238
rect 25927 -40862 25935 -40238
rect 25615 -40890 25935 -40862
rect 26615 -40238 26935 -40210
rect 26615 -40862 26623 -40238
rect 26927 -40862 26935 -40238
rect 26615 -40890 26935 -40862
rect 27615 -40238 27935 -40210
rect 27615 -40862 27623 -40238
rect 27927 -40862 27935 -40238
rect 27615 -40890 27935 -40862
rect 28615 -40238 28935 -40210
rect 28615 -40862 28623 -40238
rect 28927 -40862 28935 -40238
rect 28615 -40890 28935 -40862
rect 29615 -40238 29935 -40210
rect 29615 -40862 29623 -40238
rect 29927 -40862 29935 -40238
rect 29615 -40890 29935 -40862
rect 30615 -40238 30935 -40210
rect 30615 -40862 30623 -40238
rect 30927 -40862 30935 -40238
rect 30615 -40890 30935 -40862
rect 31615 -40238 31935 -40210
rect 31615 -40862 31623 -40238
rect 31927 -40862 31935 -40238
rect 31615 -40890 31935 -40862
rect 32615 -40238 32935 -40210
rect 32615 -40862 32623 -40238
rect 32927 -40862 32935 -40238
rect 32615 -40890 32935 -40862
rect 33615 -40238 33935 -40210
rect 33615 -40862 33623 -40238
rect 33927 -40862 33935 -40238
rect 33615 -40890 33935 -40862
rect 8275 -40898 34275 -40890
rect 8275 -41202 8283 -40898
rect 8587 -41202 8623 -40898
rect 8927 -41202 8963 -40898
rect 9587 -41202 9623 -40898
rect 9927 -41202 9963 -40898
rect 10587 -41202 10623 -40898
rect 10927 -41202 10963 -40898
rect 11587 -41202 11623 -40898
rect 11927 -41202 11963 -40898
rect 12587 -41202 12623 -40898
rect 12927 -41202 12963 -40898
rect 13587 -41202 13623 -40898
rect 13927 -41202 13963 -40898
rect 14587 -41202 14623 -40898
rect 14927 -41202 14963 -40898
rect 15587 -41202 15623 -40898
rect 15927 -41202 15963 -40898
rect 16587 -41202 16623 -40898
rect 16927 -41202 16963 -40898
rect 17587 -41202 17623 -40898
rect 17927 -41202 17963 -40898
rect 18587 -41202 18623 -40898
rect 18927 -41202 18963 -40898
rect 19587 -41202 19623 -40898
rect 19927 -41202 19963 -40898
rect 20587 -41202 20623 -40898
rect 20927 -41202 20963 -40898
rect 21587 -41202 21623 -40898
rect 21927 -41202 21963 -40898
rect 22587 -41202 22623 -40898
rect 22927 -41202 22963 -40898
rect 23587 -41202 23623 -40898
rect 23927 -41202 23963 -40898
rect 24587 -41202 24623 -40898
rect 24927 -41202 24963 -40898
rect 25587 -41202 25623 -40898
rect 25927 -41202 25963 -40898
rect 26587 -41202 26623 -40898
rect 26927 -41202 26963 -40898
rect 27587 -41202 27623 -40898
rect 27927 -41202 27963 -40898
rect 28587 -41202 28623 -40898
rect 28927 -41202 28963 -40898
rect 29587 -41202 29623 -40898
rect 29927 -41202 29963 -40898
rect 30587 -41202 30623 -40898
rect 30927 -41202 30963 -40898
rect 31587 -41202 31623 -40898
rect 31927 -41202 31963 -40898
rect 32587 -41202 32623 -40898
rect 32927 -41202 32963 -40898
rect 33587 -41202 33623 -40898
rect 33927 -41202 33963 -40898
rect 34267 -41202 34275 -40898
rect 8275 -41210 34275 -41202
rect 8615 -41238 8935 -41210
rect 8615 -41862 8623 -41238
rect 8927 -41862 8935 -41238
rect 8615 -41890 8935 -41862
rect 9615 -41238 9935 -41210
rect 9615 -41862 9623 -41238
rect 9927 -41862 9935 -41238
rect 9615 -41890 9935 -41862
rect 10615 -41238 10935 -41210
rect 10615 -41862 10623 -41238
rect 10927 -41862 10935 -41238
rect 10615 -41890 10935 -41862
rect 11615 -41238 11935 -41210
rect 11615 -41862 11623 -41238
rect 11927 -41862 11935 -41238
rect 11615 -41890 11935 -41862
rect 12615 -41238 12935 -41210
rect 12615 -41862 12623 -41238
rect 12927 -41862 12935 -41238
rect 12615 -41890 12935 -41862
rect 13615 -41238 13935 -41210
rect 13615 -41862 13623 -41238
rect 13927 -41862 13935 -41238
rect 13615 -41890 13935 -41862
rect 14615 -41238 14935 -41210
rect 14615 -41862 14623 -41238
rect 14927 -41862 14935 -41238
rect 14615 -41890 14935 -41862
rect 15615 -41238 15935 -41210
rect 15615 -41862 15623 -41238
rect 15927 -41862 15935 -41238
rect 15615 -41890 15935 -41862
rect 16615 -41238 16935 -41210
rect 16615 -41862 16623 -41238
rect 16927 -41862 16935 -41238
rect 16615 -41890 16935 -41862
rect 17615 -41238 17935 -41210
rect 17615 -41862 17623 -41238
rect 17927 -41862 17935 -41238
rect 17615 -41890 17935 -41862
rect 18615 -41238 18935 -41210
rect 18615 -41862 18623 -41238
rect 18927 -41862 18935 -41238
rect 18615 -41890 18935 -41862
rect 19615 -41238 19935 -41210
rect 19615 -41862 19623 -41238
rect 19927 -41862 19935 -41238
rect 19615 -41890 19935 -41862
rect 20615 -41238 20935 -41210
rect 20615 -41862 20623 -41238
rect 20927 -41862 20935 -41238
rect 20615 -41890 20935 -41862
rect 21615 -41238 21935 -41210
rect 21615 -41862 21623 -41238
rect 21927 -41862 21935 -41238
rect 21615 -41890 21935 -41862
rect 22615 -41238 22935 -41210
rect 22615 -41862 22623 -41238
rect 22927 -41862 22935 -41238
rect 22615 -41890 22935 -41862
rect 23615 -41238 23935 -41210
rect 23615 -41862 23623 -41238
rect 23927 -41862 23935 -41238
rect 23615 -41890 23935 -41862
rect 24615 -41238 24935 -41210
rect 24615 -41862 24623 -41238
rect 24927 -41862 24935 -41238
rect 24615 -41890 24935 -41862
rect 25615 -41238 25935 -41210
rect 25615 -41862 25623 -41238
rect 25927 -41862 25935 -41238
rect 25615 -41890 25935 -41862
rect 26615 -41238 26935 -41210
rect 26615 -41862 26623 -41238
rect 26927 -41862 26935 -41238
rect 26615 -41890 26935 -41862
rect 27615 -41238 27935 -41210
rect 27615 -41862 27623 -41238
rect 27927 -41862 27935 -41238
rect 27615 -41890 27935 -41862
rect 28615 -41238 28935 -41210
rect 28615 -41862 28623 -41238
rect 28927 -41862 28935 -41238
rect 28615 -41890 28935 -41862
rect 29615 -41238 29935 -41210
rect 29615 -41862 29623 -41238
rect 29927 -41862 29935 -41238
rect 29615 -41890 29935 -41862
rect 30615 -41238 30935 -41210
rect 30615 -41862 30623 -41238
rect 30927 -41862 30935 -41238
rect 30615 -41890 30935 -41862
rect 31615 -41238 31935 -41210
rect 31615 -41862 31623 -41238
rect 31927 -41862 31935 -41238
rect 31615 -41890 31935 -41862
rect 32615 -41238 32935 -41210
rect 32615 -41862 32623 -41238
rect 32927 -41862 32935 -41238
rect 32615 -41890 32935 -41862
rect 33615 -41238 33935 -41210
rect 33615 -41862 33623 -41238
rect 33927 -41862 33935 -41238
rect 33615 -41890 33935 -41862
rect 8275 -41898 34275 -41890
rect 8275 -42202 8283 -41898
rect 8587 -42202 8623 -41898
rect 8927 -42202 8963 -41898
rect 9587 -42202 9623 -41898
rect 9927 -42202 9963 -41898
rect 10587 -42202 10623 -41898
rect 10927 -42202 10963 -41898
rect 11587 -42202 11623 -41898
rect 11927 -42202 11963 -41898
rect 12587 -42202 12623 -41898
rect 12927 -42202 12963 -41898
rect 13587 -42202 13623 -41898
rect 13927 -42202 13963 -41898
rect 14587 -42202 14623 -41898
rect 14927 -42202 14963 -41898
rect 15587 -42202 15623 -41898
rect 15927 -42202 15963 -41898
rect 16587 -42202 16623 -41898
rect 16927 -42202 16963 -41898
rect 17587 -42202 17623 -41898
rect 17927 -42202 17963 -41898
rect 18587 -42202 18623 -41898
rect 18927 -42202 18963 -41898
rect 19587 -42202 19623 -41898
rect 19927 -42202 19963 -41898
rect 20587 -42202 20623 -41898
rect 20927 -42202 20963 -41898
rect 21587 -42202 21623 -41898
rect 21927 -42202 21963 -41898
rect 22587 -42202 22623 -41898
rect 22927 -42202 22963 -41898
rect 23587 -42202 23623 -41898
rect 23927 -42202 23963 -41898
rect 24587 -42202 24623 -41898
rect 24927 -42202 24963 -41898
rect 25587 -42202 25623 -41898
rect 25927 -42202 25963 -41898
rect 26587 -42202 26623 -41898
rect 26927 -42202 26963 -41898
rect 27587 -42202 27623 -41898
rect 27927 -42202 27963 -41898
rect 28587 -42202 28623 -41898
rect 28927 -42202 28963 -41898
rect 29587 -42202 29623 -41898
rect 29927 -42202 29963 -41898
rect 30587 -42202 30623 -41898
rect 30927 -42202 30963 -41898
rect 31587 -42202 31623 -41898
rect 31927 -42202 31963 -41898
rect 32587 -42202 32623 -41898
rect 32927 -42202 32963 -41898
rect 33587 -42202 33623 -41898
rect 33927 -42202 33963 -41898
rect 34267 -42202 34275 -41898
rect 8275 -42210 34275 -42202
rect 8615 -42238 8935 -42210
rect 8615 -42862 8623 -42238
rect 8927 -42862 8935 -42238
rect 8615 -42890 8935 -42862
rect 9615 -42238 9935 -42210
rect 9615 -42862 9623 -42238
rect 9927 -42862 9935 -42238
rect 9615 -42890 9935 -42862
rect 10615 -42238 10935 -42210
rect 10615 -42862 10623 -42238
rect 10927 -42862 10935 -42238
rect 10615 -42890 10935 -42862
rect 11615 -42238 11935 -42210
rect 11615 -42862 11623 -42238
rect 11927 -42862 11935 -42238
rect 11615 -42890 11935 -42862
rect 12615 -42238 12935 -42210
rect 12615 -42862 12623 -42238
rect 12927 -42862 12935 -42238
rect 12615 -42890 12935 -42862
rect 13615 -42238 13935 -42210
rect 13615 -42862 13623 -42238
rect 13927 -42862 13935 -42238
rect 13615 -42890 13935 -42862
rect 14615 -42238 14935 -42210
rect 14615 -42862 14623 -42238
rect 14927 -42862 14935 -42238
rect 14615 -42890 14935 -42862
rect 15615 -42238 15935 -42210
rect 15615 -42862 15623 -42238
rect 15927 -42862 15935 -42238
rect 15615 -42890 15935 -42862
rect 16615 -42238 16935 -42210
rect 16615 -42862 16623 -42238
rect 16927 -42862 16935 -42238
rect 16615 -42890 16935 -42862
rect 17615 -42238 17935 -42210
rect 17615 -42862 17623 -42238
rect 17927 -42862 17935 -42238
rect 17615 -42890 17935 -42862
rect 18615 -42238 18935 -42210
rect 18615 -42862 18623 -42238
rect 18927 -42862 18935 -42238
rect 18615 -42890 18935 -42862
rect 19615 -42238 19935 -42210
rect 19615 -42862 19623 -42238
rect 19927 -42862 19935 -42238
rect 19615 -42890 19935 -42862
rect 20615 -42238 20935 -42210
rect 20615 -42862 20623 -42238
rect 20927 -42862 20935 -42238
rect 20615 -42890 20935 -42862
rect 21615 -42238 21935 -42210
rect 21615 -42862 21623 -42238
rect 21927 -42862 21935 -42238
rect 21615 -42890 21935 -42862
rect 22615 -42238 22935 -42210
rect 22615 -42862 22623 -42238
rect 22927 -42862 22935 -42238
rect 22615 -42890 22935 -42862
rect 23615 -42238 23935 -42210
rect 23615 -42862 23623 -42238
rect 23927 -42862 23935 -42238
rect 23615 -42890 23935 -42862
rect 24615 -42238 24935 -42210
rect 24615 -42862 24623 -42238
rect 24927 -42862 24935 -42238
rect 24615 -42890 24935 -42862
rect 25615 -42238 25935 -42210
rect 25615 -42862 25623 -42238
rect 25927 -42862 25935 -42238
rect 25615 -42890 25935 -42862
rect 26615 -42238 26935 -42210
rect 26615 -42862 26623 -42238
rect 26927 -42862 26935 -42238
rect 26615 -42890 26935 -42862
rect 27615 -42238 27935 -42210
rect 27615 -42862 27623 -42238
rect 27927 -42862 27935 -42238
rect 27615 -42890 27935 -42862
rect 28615 -42238 28935 -42210
rect 28615 -42862 28623 -42238
rect 28927 -42862 28935 -42238
rect 28615 -42890 28935 -42862
rect 29615 -42238 29935 -42210
rect 29615 -42862 29623 -42238
rect 29927 -42862 29935 -42238
rect 29615 -42890 29935 -42862
rect 30615 -42238 30935 -42210
rect 30615 -42862 30623 -42238
rect 30927 -42862 30935 -42238
rect 30615 -42890 30935 -42862
rect 31615 -42238 31935 -42210
rect 31615 -42862 31623 -42238
rect 31927 -42862 31935 -42238
rect 31615 -42890 31935 -42862
rect 32615 -42238 32935 -42210
rect 32615 -42862 32623 -42238
rect 32927 -42862 32935 -42238
rect 32615 -42890 32935 -42862
rect 33615 -42238 33935 -42210
rect 33615 -42862 33623 -42238
rect 33927 -42862 33935 -42238
rect 33615 -42890 33935 -42862
rect 8275 -42898 34275 -42890
rect 8275 -43202 8283 -42898
rect 8587 -43202 8623 -42898
rect 8927 -43202 8963 -42898
rect 9587 -43202 9623 -42898
rect 9927 -43202 9963 -42898
rect 10587 -43202 10623 -42898
rect 10927 -43202 10963 -42898
rect 11587 -43202 11623 -42898
rect 11927 -43202 11963 -42898
rect 12587 -43202 12623 -42898
rect 12927 -43202 12963 -42898
rect 13587 -43202 13623 -42898
rect 13927 -43202 13963 -42898
rect 14587 -43202 14623 -42898
rect 14927 -43202 14963 -42898
rect 15587 -43202 15623 -42898
rect 15927 -43202 15963 -42898
rect 16587 -43202 16623 -42898
rect 16927 -43202 16963 -42898
rect 17587 -43202 17623 -42898
rect 17927 -43202 17963 -42898
rect 18587 -43202 18623 -42898
rect 18927 -43202 18963 -42898
rect 19587 -43202 19623 -42898
rect 19927 -43202 19963 -42898
rect 20587 -43202 20623 -42898
rect 20927 -43202 20963 -42898
rect 21587 -43202 21623 -42898
rect 21927 -43202 21963 -42898
rect 22587 -43202 22623 -42898
rect 22927 -43202 22963 -42898
rect 23587 -43202 23623 -42898
rect 23927 -43202 23963 -42898
rect 24587 -43202 24623 -42898
rect 24927 -43202 24963 -42898
rect 25587 -43202 25623 -42898
rect 25927 -43202 25963 -42898
rect 26587 -43202 26623 -42898
rect 26927 -43202 26963 -42898
rect 27587 -43202 27623 -42898
rect 27927 -43202 27963 -42898
rect 28587 -43202 28623 -42898
rect 28927 -43202 28963 -42898
rect 29587 -43202 29623 -42898
rect 29927 -43202 29963 -42898
rect 30587 -43202 30623 -42898
rect 30927 -43202 30963 -42898
rect 31587 -43202 31623 -42898
rect 31927 -43202 31963 -42898
rect 32587 -43202 32623 -42898
rect 32927 -43202 32963 -42898
rect 33587 -43202 33623 -42898
rect 33927 -43202 33963 -42898
rect 34267 -43202 34275 -42898
rect 8275 -43210 34275 -43202
rect 8615 -43238 8935 -43210
rect 8615 -43862 8623 -43238
rect 8927 -43862 8935 -43238
rect 8615 -43890 8935 -43862
rect 9615 -43238 9935 -43210
rect 9615 -43862 9623 -43238
rect 9927 -43862 9935 -43238
rect 9615 -43890 9935 -43862
rect 10615 -43238 10935 -43210
rect 10615 -43862 10623 -43238
rect 10927 -43862 10935 -43238
rect 10615 -43890 10935 -43862
rect 11615 -43238 11935 -43210
rect 11615 -43862 11623 -43238
rect 11927 -43862 11935 -43238
rect 11615 -43890 11935 -43862
rect 12615 -43238 12935 -43210
rect 12615 -43862 12623 -43238
rect 12927 -43862 12935 -43238
rect 12615 -43890 12935 -43862
rect 13615 -43238 13935 -43210
rect 13615 -43862 13623 -43238
rect 13927 -43862 13935 -43238
rect 13615 -43890 13935 -43862
rect 14615 -43238 14935 -43210
rect 14615 -43862 14623 -43238
rect 14927 -43862 14935 -43238
rect 14615 -43890 14935 -43862
rect 15615 -43238 15935 -43210
rect 15615 -43862 15623 -43238
rect 15927 -43862 15935 -43238
rect 15615 -43890 15935 -43862
rect 16615 -43238 16935 -43210
rect 16615 -43862 16623 -43238
rect 16927 -43862 16935 -43238
rect 16615 -43890 16935 -43862
rect 17615 -43238 17935 -43210
rect 17615 -43862 17623 -43238
rect 17927 -43862 17935 -43238
rect 17615 -43890 17935 -43862
rect 18615 -43238 18935 -43210
rect 18615 -43862 18623 -43238
rect 18927 -43862 18935 -43238
rect 18615 -43890 18935 -43862
rect 19615 -43238 19935 -43210
rect 19615 -43862 19623 -43238
rect 19927 -43862 19935 -43238
rect 19615 -43890 19935 -43862
rect 20615 -43238 20935 -43210
rect 20615 -43862 20623 -43238
rect 20927 -43862 20935 -43238
rect 20615 -43890 20935 -43862
rect 21615 -43238 21935 -43210
rect 21615 -43862 21623 -43238
rect 21927 -43862 21935 -43238
rect 21615 -43890 21935 -43862
rect 22615 -43238 22935 -43210
rect 22615 -43862 22623 -43238
rect 22927 -43862 22935 -43238
rect 22615 -43890 22935 -43862
rect 23615 -43238 23935 -43210
rect 23615 -43862 23623 -43238
rect 23927 -43862 23935 -43238
rect 23615 -43890 23935 -43862
rect 24615 -43238 24935 -43210
rect 24615 -43862 24623 -43238
rect 24927 -43862 24935 -43238
rect 24615 -43890 24935 -43862
rect 25615 -43238 25935 -43210
rect 25615 -43862 25623 -43238
rect 25927 -43862 25935 -43238
rect 25615 -43890 25935 -43862
rect 26615 -43238 26935 -43210
rect 26615 -43862 26623 -43238
rect 26927 -43862 26935 -43238
rect 26615 -43890 26935 -43862
rect 27615 -43238 27935 -43210
rect 27615 -43862 27623 -43238
rect 27927 -43862 27935 -43238
rect 27615 -43890 27935 -43862
rect 28615 -43238 28935 -43210
rect 28615 -43862 28623 -43238
rect 28927 -43862 28935 -43238
rect 28615 -43890 28935 -43862
rect 29615 -43238 29935 -43210
rect 29615 -43862 29623 -43238
rect 29927 -43862 29935 -43238
rect 29615 -43890 29935 -43862
rect 30615 -43238 30935 -43210
rect 30615 -43862 30623 -43238
rect 30927 -43862 30935 -43238
rect 30615 -43890 30935 -43862
rect 31615 -43238 31935 -43210
rect 31615 -43862 31623 -43238
rect 31927 -43862 31935 -43238
rect 31615 -43890 31935 -43862
rect 32615 -43238 32935 -43210
rect 32615 -43862 32623 -43238
rect 32927 -43862 32935 -43238
rect 32615 -43890 32935 -43862
rect 33615 -43238 33935 -43210
rect 33615 -43862 33623 -43238
rect 33927 -43862 33935 -43238
rect 33615 -43890 33935 -43862
rect 8275 -43898 34275 -43890
rect 8275 -44202 8283 -43898
rect 8587 -44202 8623 -43898
rect 8927 -44202 8963 -43898
rect 9587 -44202 9623 -43898
rect 9927 -44202 9963 -43898
rect 10587 -44202 10623 -43898
rect 10927 -44202 10963 -43898
rect 11587 -44202 11623 -43898
rect 11927 -44202 11963 -43898
rect 12587 -44202 12623 -43898
rect 12927 -44202 12963 -43898
rect 13587 -44202 13623 -43898
rect 13927 -44202 13963 -43898
rect 14587 -44202 14623 -43898
rect 14927 -44202 14963 -43898
rect 15587 -44202 15623 -43898
rect 15927 -44202 15963 -43898
rect 16587 -44202 16623 -43898
rect 16927 -44202 16963 -43898
rect 17587 -44202 17623 -43898
rect 17927 -44202 17963 -43898
rect 18587 -44202 18623 -43898
rect 18927 -44202 18963 -43898
rect 19587 -44202 19623 -43898
rect 19927 -44202 19963 -43898
rect 20587 -44202 20623 -43898
rect 20927 -44202 20963 -43898
rect 21587 -44202 21623 -43898
rect 21927 -44202 21963 -43898
rect 22587 -44202 22623 -43898
rect 22927 -44202 22963 -43898
rect 23587 -44202 23623 -43898
rect 23927 -44202 23963 -43898
rect 24587 -44202 24623 -43898
rect 24927 -44202 24963 -43898
rect 25587 -44202 25623 -43898
rect 25927 -44202 25963 -43898
rect 26587 -44202 26623 -43898
rect 26927 -44202 26963 -43898
rect 27587 -44202 27623 -43898
rect 27927 -44202 27963 -43898
rect 28587 -44202 28623 -43898
rect 28927 -44202 28963 -43898
rect 29587 -44202 29623 -43898
rect 29927 -44202 29963 -43898
rect 30587 -44202 30623 -43898
rect 30927 -44202 30963 -43898
rect 31587 -44202 31623 -43898
rect 31927 -44202 31963 -43898
rect 32587 -44202 32623 -43898
rect 32927 -44202 32963 -43898
rect 33587 -44202 33623 -43898
rect 33927 -44202 33963 -43898
rect 34267 -44202 34275 -43898
rect 8275 -44210 34275 -44202
rect -4275 -44550 5725 -44502
rect 8615 -44238 8935 -44210
rect -49485 -44890 -49165 -44862
rect 8615 -44862 8623 -44238
rect 8927 -44862 8935 -44238
rect 8615 -44890 8935 -44862
rect 9615 -44238 9935 -44210
rect 9615 -44862 9623 -44238
rect 9927 -44862 9935 -44238
rect 9615 -44890 9935 -44862
rect 10615 -44238 10935 -44210
rect 10615 -44862 10623 -44238
rect 10927 -44862 10935 -44238
rect 10615 -44890 10935 -44862
rect 11615 -44238 11935 -44210
rect 11615 -44862 11623 -44238
rect 11927 -44862 11935 -44238
rect 11615 -44890 11935 -44862
rect 12615 -44238 12935 -44210
rect 12615 -44862 12623 -44238
rect 12927 -44862 12935 -44238
rect 12615 -44890 12935 -44862
rect 13615 -44238 13935 -44210
rect 13615 -44862 13623 -44238
rect 13927 -44862 13935 -44238
rect 13615 -44890 13935 -44862
rect 14615 -44238 14935 -44210
rect 14615 -44862 14623 -44238
rect 14927 -44862 14935 -44238
rect 14615 -44890 14935 -44862
rect 15615 -44238 15935 -44210
rect 15615 -44862 15623 -44238
rect 15927 -44862 15935 -44238
rect 15615 -44890 15935 -44862
rect 16615 -44238 16935 -44210
rect 16615 -44862 16623 -44238
rect 16927 -44862 16935 -44238
rect 16615 -44890 16935 -44862
rect 17615 -44238 17935 -44210
rect 17615 -44862 17623 -44238
rect 17927 -44862 17935 -44238
rect 17615 -44890 17935 -44862
rect 18615 -44238 18935 -44210
rect 18615 -44862 18623 -44238
rect 18927 -44862 18935 -44238
rect 18615 -44890 18935 -44862
rect 19615 -44238 19935 -44210
rect 19615 -44862 19623 -44238
rect 19927 -44862 19935 -44238
rect 19615 -44890 19935 -44862
rect 20615 -44238 20935 -44210
rect 20615 -44862 20623 -44238
rect 20927 -44862 20935 -44238
rect 20615 -44890 20935 -44862
rect 21615 -44238 21935 -44210
rect 21615 -44862 21623 -44238
rect 21927 -44862 21935 -44238
rect 21615 -44890 21935 -44862
rect 22615 -44238 22935 -44210
rect 22615 -44862 22623 -44238
rect 22927 -44862 22935 -44238
rect 22615 -44890 22935 -44862
rect 23615 -44238 23935 -44210
rect 23615 -44862 23623 -44238
rect 23927 -44862 23935 -44238
rect 23615 -44890 23935 -44862
rect 24615 -44238 24935 -44210
rect 24615 -44862 24623 -44238
rect 24927 -44862 24935 -44238
rect 24615 -44890 24935 -44862
rect 25615 -44238 25935 -44210
rect 25615 -44862 25623 -44238
rect 25927 -44862 25935 -44238
rect 25615 -44890 25935 -44862
rect 26615 -44238 26935 -44210
rect 26615 -44862 26623 -44238
rect 26927 -44862 26935 -44238
rect 26615 -44890 26935 -44862
rect 27615 -44238 27935 -44210
rect 27615 -44862 27623 -44238
rect 27927 -44862 27935 -44238
rect 27615 -44890 27935 -44862
rect 28615 -44238 28935 -44210
rect 28615 -44862 28623 -44238
rect 28927 -44862 28935 -44238
rect 28615 -44890 28935 -44862
rect 29615 -44238 29935 -44210
rect 29615 -44862 29623 -44238
rect 29927 -44862 29935 -44238
rect 29615 -44890 29935 -44862
rect 30615 -44238 30935 -44210
rect 30615 -44862 30623 -44238
rect 30927 -44862 30935 -44238
rect 30615 -44890 30935 -44862
rect 31615 -44238 31935 -44210
rect 31615 -44862 31623 -44238
rect 31927 -44862 31935 -44238
rect 31615 -44890 31935 -44862
rect 32615 -44238 32935 -44210
rect 32615 -44862 32623 -44238
rect 32927 -44862 32935 -44238
rect 32615 -44890 32935 -44862
rect 33615 -44238 33935 -44210
rect 33615 -44862 33623 -44238
rect 33927 -44862 33935 -44238
rect 33615 -44890 33935 -44862
rect -74825 -44898 -48825 -44890
rect -74825 -45202 -74817 -44898
rect -74513 -45202 -74477 -44898
rect -74173 -45202 -74137 -44898
rect -73513 -45202 -73477 -44898
rect -73173 -45202 -73137 -44898
rect -72513 -45202 -72477 -44898
rect -72173 -45202 -72137 -44898
rect -71513 -45202 -71477 -44898
rect -71173 -45202 -71137 -44898
rect -70513 -45202 -70477 -44898
rect -70173 -45202 -70137 -44898
rect -69513 -45202 -69477 -44898
rect -69173 -45202 -69137 -44898
rect -68513 -45202 -68477 -44898
rect -68173 -45202 -68137 -44898
rect -67513 -45202 -67477 -44898
rect -67173 -45202 -67137 -44898
rect -66513 -45202 -66477 -44898
rect -66173 -45202 -66137 -44898
rect -65513 -45202 -65477 -44898
rect -65173 -45202 -65137 -44898
rect -64513 -45202 -64477 -44898
rect -64173 -45202 -64137 -44898
rect -63513 -45202 -63477 -44898
rect -63173 -45202 -63137 -44898
rect -62513 -45202 -62477 -44898
rect -62173 -45202 -62137 -44898
rect -61513 -45202 -61477 -44898
rect -61173 -45202 -61137 -44898
rect -60513 -45202 -60477 -44898
rect -60173 -45202 -60137 -44898
rect -59513 -45202 -59477 -44898
rect -59173 -45202 -59137 -44898
rect -58513 -45202 -58477 -44898
rect -58173 -45202 -58137 -44898
rect -57513 -45202 -57477 -44898
rect -57173 -45202 -57137 -44898
rect -56513 -45202 -56477 -44898
rect -56173 -45202 -56137 -44898
rect -55513 -45202 -55477 -44898
rect -55173 -45202 -55137 -44898
rect -54513 -45202 -54477 -44898
rect -54173 -45202 -54137 -44898
rect -53513 -45202 -53477 -44898
rect -53173 -45202 -53137 -44898
rect -52513 -45202 -52477 -44898
rect -52173 -45202 -52137 -44898
rect -51513 -45202 -51477 -44898
rect -51173 -45202 -51137 -44898
rect -50513 -45202 -50477 -44898
rect -50173 -45202 -50137 -44898
rect -49513 -45202 -49477 -44898
rect -49173 -45202 -49137 -44898
rect -48833 -45202 -48825 -44898
rect -74825 -45210 -48825 -45202
rect 8275 -44898 34275 -44890
rect 8275 -45202 8283 -44898
rect 8587 -45202 8623 -44898
rect 8927 -45202 8963 -44898
rect 9587 -45202 9623 -44898
rect 9927 -45202 9963 -44898
rect 10587 -45202 10623 -44898
rect 10927 -45202 10963 -44898
rect 11587 -45202 11623 -44898
rect 11927 -45202 11963 -44898
rect 12587 -45202 12623 -44898
rect 12927 -45202 12963 -44898
rect 13587 -45202 13623 -44898
rect 13927 -45202 13963 -44898
rect 14587 -45202 14623 -44898
rect 14927 -45202 14963 -44898
rect 15587 -45202 15623 -44898
rect 15927 -45202 15963 -44898
rect 16587 -45202 16623 -44898
rect 16927 -45202 16963 -44898
rect 17587 -45202 17623 -44898
rect 17927 -45202 17963 -44898
rect 18587 -45202 18623 -44898
rect 18927 -45202 18963 -44898
rect 19587 -45202 19623 -44898
rect 19927 -45202 19963 -44898
rect 20587 -45202 20623 -44898
rect 20927 -45202 20963 -44898
rect 21587 -45202 21623 -44898
rect 21927 -45202 21963 -44898
rect 22587 -45202 22623 -44898
rect 22927 -45202 22963 -44898
rect 23587 -45202 23623 -44898
rect 23927 -45202 23963 -44898
rect 24587 -45202 24623 -44898
rect 24927 -45202 24963 -44898
rect 25587 -45202 25623 -44898
rect 25927 -45202 25963 -44898
rect 26587 -45202 26623 -44898
rect 26927 -45202 26963 -44898
rect 27587 -45202 27623 -44898
rect 27927 -45202 27963 -44898
rect 28587 -45202 28623 -44898
rect 28927 -45202 28963 -44898
rect 29587 -45202 29623 -44898
rect 29927 -45202 29963 -44898
rect 30587 -45202 30623 -44898
rect 30927 -45202 30963 -44898
rect 31587 -45202 31623 -44898
rect 31927 -45202 31963 -44898
rect 32587 -45202 32623 -44898
rect 32927 -45202 32963 -44898
rect 33587 -45202 33623 -44898
rect 33927 -45202 33963 -44898
rect 34267 -45202 34275 -44898
rect 8275 -45210 34275 -45202
rect -74485 -45238 -74165 -45210
rect -74485 -45862 -74477 -45238
rect -74173 -45862 -74165 -45238
rect -74485 -45890 -74165 -45862
rect -73485 -45238 -73165 -45210
rect -73485 -45862 -73477 -45238
rect -73173 -45862 -73165 -45238
rect -73485 -45890 -73165 -45862
rect -72485 -45238 -72165 -45210
rect -72485 -45862 -72477 -45238
rect -72173 -45862 -72165 -45238
rect -72485 -45890 -72165 -45862
rect -71485 -45238 -71165 -45210
rect -71485 -45862 -71477 -45238
rect -71173 -45862 -71165 -45238
rect -71485 -45890 -71165 -45862
rect -70485 -45238 -70165 -45210
rect -70485 -45862 -70477 -45238
rect -70173 -45862 -70165 -45238
rect -70485 -45890 -70165 -45862
rect -69485 -45238 -69165 -45210
rect -69485 -45862 -69477 -45238
rect -69173 -45862 -69165 -45238
rect -69485 -45890 -69165 -45862
rect -68485 -45238 -68165 -45210
rect -68485 -45862 -68477 -45238
rect -68173 -45862 -68165 -45238
rect -68485 -45890 -68165 -45862
rect -67485 -45238 -67165 -45210
rect -67485 -45862 -67477 -45238
rect -67173 -45862 -67165 -45238
rect -67485 -45890 -67165 -45862
rect -66485 -45238 -66165 -45210
rect -66485 -45862 -66477 -45238
rect -66173 -45862 -66165 -45238
rect -66485 -45890 -66165 -45862
rect -65485 -45238 -65165 -45210
rect -65485 -45862 -65477 -45238
rect -65173 -45862 -65165 -45238
rect -65485 -45890 -65165 -45862
rect -64485 -45238 -64165 -45210
rect -64485 -45862 -64477 -45238
rect -64173 -45862 -64165 -45238
rect -64485 -45890 -64165 -45862
rect -63485 -45238 -63165 -45210
rect -63485 -45862 -63477 -45238
rect -63173 -45862 -63165 -45238
rect -63485 -45890 -63165 -45862
rect -62485 -45238 -62165 -45210
rect -62485 -45862 -62477 -45238
rect -62173 -45862 -62165 -45238
rect -62485 -45890 -62165 -45862
rect -61485 -45238 -61165 -45210
rect -61485 -45862 -61477 -45238
rect -61173 -45862 -61165 -45238
rect -61485 -45890 -61165 -45862
rect -60485 -45238 -60165 -45210
rect -60485 -45862 -60477 -45238
rect -60173 -45862 -60165 -45238
rect -60485 -45890 -60165 -45862
rect -59485 -45238 -59165 -45210
rect -59485 -45862 -59477 -45238
rect -59173 -45862 -59165 -45238
rect -59485 -45890 -59165 -45862
rect -58485 -45238 -58165 -45210
rect -58485 -45862 -58477 -45238
rect -58173 -45862 -58165 -45238
rect -58485 -45890 -58165 -45862
rect -57485 -45238 -57165 -45210
rect -57485 -45862 -57477 -45238
rect -57173 -45862 -57165 -45238
rect -57485 -45890 -57165 -45862
rect -56485 -45238 -56165 -45210
rect -56485 -45862 -56477 -45238
rect -56173 -45862 -56165 -45238
rect -56485 -45890 -56165 -45862
rect -55485 -45238 -55165 -45210
rect -55485 -45862 -55477 -45238
rect -55173 -45862 -55165 -45238
rect -55485 -45890 -55165 -45862
rect -54485 -45238 -54165 -45210
rect -54485 -45862 -54477 -45238
rect -54173 -45862 -54165 -45238
rect -54485 -45890 -54165 -45862
rect -53485 -45238 -53165 -45210
rect -53485 -45862 -53477 -45238
rect -53173 -45862 -53165 -45238
rect -53485 -45890 -53165 -45862
rect -52485 -45238 -52165 -45210
rect -52485 -45862 -52477 -45238
rect -52173 -45862 -52165 -45238
rect -52485 -45890 -52165 -45862
rect -51485 -45238 -51165 -45210
rect -51485 -45862 -51477 -45238
rect -51173 -45862 -51165 -45238
rect -51485 -45890 -51165 -45862
rect -50485 -45238 -50165 -45210
rect -50485 -45862 -50477 -45238
rect -50173 -45862 -50165 -45238
rect -50485 -45890 -50165 -45862
rect -49485 -45238 -49165 -45210
rect -49485 -45862 -49477 -45238
rect -49173 -45862 -49165 -45238
rect -49485 -45890 -49165 -45862
rect 8615 -45238 8935 -45210
rect 8615 -45862 8623 -45238
rect 8927 -45862 8935 -45238
rect 8615 -45890 8935 -45862
rect 9615 -45238 9935 -45210
rect 9615 -45862 9623 -45238
rect 9927 -45862 9935 -45238
rect 9615 -45890 9935 -45862
rect 10615 -45238 10935 -45210
rect 10615 -45862 10623 -45238
rect 10927 -45862 10935 -45238
rect 10615 -45890 10935 -45862
rect 11615 -45238 11935 -45210
rect 11615 -45862 11623 -45238
rect 11927 -45862 11935 -45238
rect 11615 -45890 11935 -45862
rect 12615 -45238 12935 -45210
rect 12615 -45862 12623 -45238
rect 12927 -45862 12935 -45238
rect 12615 -45890 12935 -45862
rect 13615 -45238 13935 -45210
rect 13615 -45862 13623 -45238
rect 13927 -45862 13935 -45238
rect 13615 -45890 13935 -45862
rect 14615 -45238 14935 -45210
rect 14615 -45862 14623 -45238
rect 14927 -45862 14935 -45238
rect 14615 -45890 14935 -45862
rect 15615 -45238 15935 -45210
rect 15615 -45862 15623 -45238
rect 15927 -45862 15935 -45238
rect 15615 -45890 15935 -45862
rect 16615 -45238 16935 -45210
rect 16615 -45862 16623 -45238
rect 16927 -45862 16935 -45238
rect 16615 -45890 16935 -45862
rect 17615 -45238 17935 -45210
rect 17615 -45862 17623 -45238
rect 17927 -45862 17935 -45238
rect 17615 -45890 17935 -45862
rect 18615 -45238 18935 -45210
rect 18615 -45862 18623 -45238
rect 18927 -45862 18935 -45238
rect 18615 -45890 18935 -45862
rect 19615 -45238 19935 -45210
rect 19615 -45862 19623 -45238
rect 19927 -45862 19935 -45238
rect 19615 -45890 19935 -45862
rect 20615 -45238 20935 -45210
rect 20615 -45862 20623 -45238
rect 20927 -45862 20935 -45238
rect 20615 -45890 20935 -45862
rect 21615 -45238 21935 -45210
rect 21615 -45862 21623 -45238
rect 21927 -45862 21935 -45238
rect 21615 -45890 21935 -45862
rect 22615 -45238 22935 -45210
rect 22615 -45862 22623 -45238
rect 22927 -45862 22935 -45238
rect 22615 -45890 22935 -45862
rect 23615 -45238 23935 -45210
rect 23615 -45862 23623 -45238
rect 23927 -45862 23935 -45238
rect 23615 -45890 23935 -45862
rect 24615 -45238 24935 -45210
rect 24615 -45862 24623 -45238
rect 24927 -45862 24935 -45238
rect 24615 -45890 24935 -45862
rect 25615 -45238 25935 -45210
rect 25615 -45862 25623 -45238
rect 25927 -45862 25935 -45238
rect 25615 -45890 25935 -45862
rect 26615 -45238 26935 -45210
rect 26615 -45862 26623 -45238
rect 26927 -45862 26935 -45238
rect 26615 -45890 26935 -45862
rect 27615 -45238 27935 -45210
rect 27615 -45862 27623 -45238
rect 27927 -45862 27935 -45238
rect 27615 -45890 27935 -45862
rect 28615 -45238 28935 -45210
rect 28615 -45862 28623 -45238
rect 28927 -45862 28935 -45238
rect 28615 -45890 28935 -45862
rect 29615 -45238 29935 -45210
rect 29615 -45862 29623 -45238
rect 29927 -45862 29935 -45238
rect 29615 -45890 29935 -45862
rect 30615 -45238 30935 -45210
rect 30615 -45862 30623 -45238
rect 30927 -45862 30935 -45238
rect 30615 -45890 30935 -45862
rect 31615 -45238 31935 -45210
rect 31615 -45862 31623 -45238
rect 31927 -45862 31935 -45238
rect 31615 -45890 31935 -45862
rect 32615 -45238 32935 -45210
rect 32615 -45862 32623 -45238
rect 32927 -45862 32935 -45238
rect 32615 -45890 32935 -45862
rect 33615 -45238 33935 -45210
rect 33615 -45862 33623 -45238
rect 33927 -45862 33935 -45238
rect 33615 -45890 33935 -45862
rect -74825 -45898 -48825 -45890
rect -74825 -46202 -74817 -45898
rect -74513 -46202 -74477 -45898
rect -74173 -46202 -74137 -45898
rect -73513 -46202 -73477 -45898
rect -73173 -46202 -73137 -45898
rect -72513 -46202 -72477 -45898
rect -72173 -46202 -72137 -45898
rect -71513 -46202 -71477 -45898
rect -71173 -46202 -71137 -45898
rect -70513 -46202 -70477 -45898
rect -70173 -46202 -70137 -45898
rect -69513 -46202 -69477 -45898
rect -69173 -46202 -69137 -45898
rect -68513 -46202 -68477 -45898
rect -68173 -46202 -68137 -45898
rect -67513 -46202 -67477 -45898
rect -67173 -46202 -67137 -45898
rect -66513 -46202 -66477 -45898
rect -66173 -46202 -66137 -45898
rect -65513 -46202 -65477 -45898
rect -65173 -46202 -65137 -45898
rect -64513 -46202 -64477 -45898
rect -64173 -46202 -64137 -45898
rect -63513 -46202 -63477 -45898
rect -63173 -46202 -63137 -45898
rect -62513 -46202 -62477 -45898
rect -62173 -46202 -62137 -45898
rect -61513 -46202 -61477 -45898
rect -61173 -46202 -61137 -45898
rect -60513 -46202 -60477 -45898
rect -60173 -46202 -60137 -45898
rect -59513 -46202 -59477 -45898
rect -59173 -46202 -59137 -45898
rect -58513 -46202 -58477 -45898
rect -58173 -46202 -58137 -45898
rect -57513 -46202 -57477 -45898
rect -57173 -46202 -57137 -45898
rect -56513 -46202 -56477 -45898
rect -56173 -46202 -56137 -45898
rect -55513 -46202 -55477 -45898
rect -55173 -46202 -55137 -45898
rect -54513 -46202 -54477 -45898
rect -54173 -46202 -54137 -45898
rect -53513 -46202 -53477 -45898
rect -53173 -46202 -53137 -45898
rect -52513 -46202 -52477 -45898
rect -52173 -46202 -52137 -45898
rect -51513 -46202 -51477 -45898
rect -51173 -46202 -51137 -45898
rect -50513 -46202 -50477 -45898
rect -50173 -46202 -50137 -45898
rect -49513 -46202 -49477 -45898
rect -49173 -46202 -49137 -45898
rect -48833 -46202 -48825 -45898
rect -74825 -46210 -48825 -46202
rect 8275 -45898 34275 -45890
rect 8275 -46202 8283 -45898
rect 8587 -46202 8623 -45898
rect 8927 -46202 8963 -45898
rect 9587 -46202 9623 -45898
rect 9927 -46202 9963 -45898
rect 10587 -46202 10623 -45898
rect 10927 -46202 10963 -45898
rect 11587 -46202 11623 -45898
rect 11927 -46202 11963 -45898
rect 12587 -46202 12623 -45898
rect 12927 -46202 12963 -45898
rect 13587 -46202 13623 -45898
rect 13927 -46202 13963 -45898
rect 14587 -46202 14623 -45898
rect 14927 -46202 14963 -45898
rect 15587 -46202 15623 -45898
rect 15927 -46202 15963 -45898
rect 16587 -46202 16623 -45898
rect 16927 -46202 16963 -45898
rect 17587 -46202 17623 -45898
rect 17927 -46202 17963 -45898
rect 18587 -46202 18623 -45898
rect 18927 -46202 18963 -45898
rect 19587 -46202 19623 -45898
rect 19927 -46202 19963 -45898
rect 20587 -46202 20623 -45898
rect 20927 -46202 20963 -45898
rect 21587 -46202 21623 -45898
rect 21927 -46202 21963 -45898
rect 22587 -46202 22623 -45898
rect 22927 -46202 22963 -45898
rect 23587 -46202 23623 -45898
rect 23927 -46202 23963 -45898
rect 24587 -46202 24623 -45898
rect 24927 -46202 24963 -45898
rect 25587 -46202 25623 -45898
rect 25927 -46202 25963 -45898
rect 26587 -46202 26623 -45898
rect 26927 -46202 26963 -45898
rect 27587 -46202 27623 -45898
rect 27927 -46202 27963 -45898
rect 28587 -46202 28623 -45898
rect 28927 -46202 28963 -45898
rect 29587 -46202 29623 -45898
rect 29927 -46202 29963 -45898
rect 30587 -46202 30623 -45898
rect 30927 -46202 30963 -45898
rect 31587 -46202 31623 -45898
rect 31927 -46202 31963 -45898
rect 32587 -46202 32623 -45898
rect 32927 -46202 32963 -45898
rect 33587 -46202 33623 -45898
rect 33927 -46202 33963 -45898
rect 34267 -46202 34275 -45898
rect 8275 -46210 34275 -46202
rect -74485 -46238 -74165 -46210
rect -74485 -46542 -74477 -46238
rect -74173 -46542 -74165 -46238
rect -74485 -46550 -74165 -46542
rect -73485 -46238 -73165 -46210
rect -73485 -46542 -73477 -46238
rect -73173 -46542 -73165 -46238
rect -73485 -46550 -73165 -46542
rect -72485 -46238 -72165 -46210
rect -72485 -46542 -72477 -46238
rect -72173 -46542 -72165 -46238
rect -72485 -46550 -72165 -46542
rect -71485 -46238 -71165 -46210
rect -71485 -46542 -71477 -46238
rect -71173 -46542 -71165 -46238
rect -71485 -46550 -71165 -46542
rect -70485 -46238 -70165 -46210
rect -70485 -46542 -70477 -46238
rect -70173 -46542 -70165 -46238
rect -70485 -46550 -70165 -46542
rect -69485 -46238 -69165 -46210
rect -69485 -46542 -69477 -46238
rect -69173 -46542 -69165 -46238
rect -69485 -46550 -69165 -46542
rect -68485 -46238 -68165 -46210
rect -68485 -46542 -68477 -46238
rect -68173 -46542 -68165 -46238
rect -68485 -46550 -68165 -46542
rect -67485 -46238 -67165 -46210
rect -67485 -46542 -67477 -46238
rect -67173 -46542 -67165 -46238
rect -67485 -46550 -67165 -46542
rect -66485 -46238 -66165 -46210
rect -66485 -46542 -66477 -46238
rect -66173 -46542 -66165 -46238
rect -66485 -46550 -66165 -46542
rect -65485 -46238 -65165 -46210
rect -65485 -46542 -65477 -46238
rect -65173 -46542 -65165 -46238
rect -65485 -46550 -65165 -46542
rect -64485 -46238 -64165 -46210
rect -64485 -46542 -64477 -46238
rect -64173 -46542 -64165 -46238
rect -64485 -46550 -64165 -46542
rect -63485 -46238 -63165 -46210
rect -63485 -46542 -63477 -46238
rect -63173 -46542 -63165 -46238
rect -63485 -46550 -63165 -46542
rect -62485 -46238 -62165 -46210
rect -62485 -46542 -62477 -46238
rect -62173 -46542 -62165 -46238
rect -62485 -46550 -62165 -46542
rect -61485 -46238 -61165 -46210
rect -61485 -46542 -61477 -46238
rect -61173 -46542 -61165 -46238
rect -61485 -46550 -61165 -46542
rect -60485 -46238 -60165 -46210
rect -60485 -46542 -60477 -46238
rect -60173 -46542 -60165 -46238
rect -60485 -46550 -60165 -46542
rect -59485 -46238 -59165 -46210
rect -59485 -46542 -59477 -46238
rect -59173 -46542 -59165 -46238
rect -59485 -46550 -59165 -46542
rect -58485 -46238 -58165 -46210
rect -58485 -46542 -58477 -46238
rect -58173 -46542 -58165 -46238
rect -58485 -46550 -58165 -46542
rect -57485 -46238 -57165 -46210
rect -57485 -46542 -57477 -46238
rect -57173 -46542 -57165 -46238
rect -57485 -46550 -57165 -46542
rect -56485 -46238 -56165 -46210
rect -56485 -46542 -56477 -46238
rect -56173 -46542 -56165 -46238
rect -56485 -46550 -56165 -46542
rect -55485 -46238 -55165 -46210
rect -55485 -46542 -55477 -46238
rect -55173 -46542 -55165 -46238
rect -55485 -46550 -55165 -46542
rect -54485 -46238 -54165 -46210
rect -54485 -46542 -54477 -46238
rect -54173 -46542 -54165 -46238
rect -54485 -46550 -54165 -46542
rect -53485 -46238 -53165 -46210
rect -53485 -46542 -53477 -46238
rect -53173 -46542 -53165 -46238
rect -53485 -46550 -53165 -46542
rect -52485 -46238 -52165 -46210
rect -52485 -46542 -52477 -46238
rect -52173 -46542 -52165 -46238
rect -52485 -46550 -52165 -46542
rect -51485 -46238 -51165 -46210
rect -51485 -46542 -51477 -46238
rect -51173 -46542 -51165 -46238
rect -51485 -46550 -51165 -46542
rect -50485 -46238 -50165 -46210
rect -50485 -46542 -50477 -46238
rect -50173 -46542 -50165 -46238
rect -50485 -46550 -50165 -46542
rect -49485 -46238 -49165 -46210
rect -49485 -46542 -49477 -46238
rect -49173 -46542 -49165 -46238
rect -49485 -46550 -49165 -46542
rect 8615 -46238 8935 -46210
rect 8615 -46542 8623 -46238
rect 8927 -46542 8935 -46238
rect 8615 -46550 8935 -46542
rect 9615 -46238 9935 -46210
rect 9615 -46542 9623 -46238
rect 9927 -46542 9935 -46238
rect 9615 -46550 9935 -46542
rect 10615 -46238 10935 -46210
rect 10615 -46542 10623 -46238
rect 10927 -46542 10935 -46238
rect 10615 -46550 10935 -46542
rect 11615 -46238 11935 -46210
rect 11615 -46542 11623 -46238
rect 11927 -46542 11935 -46238
rect 11615 -46550 11935 -46542
rect 12615 -46238 12935 -46210
rect 12615 -46542 12623 -46238
rect 12927 -46542 12935 -46238
rect 12615 -46550 12935 -46542
rect 13615 -46238 13935 -46210
rect 13615 -46542 13623 -46238
rect 13927 -46542 13935 -46238
rect 13615 -46550 13935 -46542
rect 14615 -46238 14935 -46210
rect 14615 -46542 14623 -46238
rect 14927 -46542 14935 -46238
rect 14615 -46550 14935 -46542
rect 15615 -46238 15935 -46210
rect 15615 -46542 15623 -46238
rect 15927 -46542 15935 -46238
rect 15615 -46550 15935 -46542
rect 16615 -46238 16935 -46210
rect 16615 -46542 16623 -46238
rect 16927 -46542 16935 -46238
rect 16615 -46550 16935 -46542
rect 17615 -46238 17935 -46210
rect 17615 -46542 17623 -46238
rect 17927 -46542 17935 -46238
rect 17615 -46550 17935 -46542
rect 18615 -46238 18935 -46210
rect 18615 -46542 18623 -46238
rect 18927 -46542 18935 -46238
rect 18615 -46550 18935 -46542
rect 19615 -46238 19935 -46210
rect 19615 -46542 19623 -46238
rect 19927 -46542 19935 -46238
rect 19615 -46550 19935 -46542
rect 20615 -46238 20935 -46210
rect 20615 -46542 20623 -46238
rect 20927 -46542 20935 -46238
rect 20615 -46550 20935 -46542
rect 21615 -46238 21935 -46210
rect 21615 -46542 21623 -46238
rect 21927 -46542 21935 -46238
rect 21615 -46550 21935 -46542
rect 22615 -46238 22935 -46210
rect 22615 -46542 22623 -46238
rect 22927 -46542 22935 -46238
rect 22615 -46550 22935 -46542
rect 23615 -46238 23935 -46210
rect 23615 -46542 23623 -46238
rect 23927 -46542 23935 -46238
rect 23615 -46550 23935 -46542
rect 24615 -46238 24935 -46210
rect 24615 -46542 24623 -46238
rect 24927 -46542 24935 -46238
rect 24615 -46550 24935 -46542
rect 25615 -46238 25935 -46210
rect 25615 -46542 25623 -46238
rect 25927 -46542 25935 -46238
rect 25615 -46550 25935 -46542
rect 26615 -46238 26935 -46210
rect 26615 -46542 26623 -46238
rect 26927 -46542 26935 -46238
rect 26615 -46550 26935 -46542
rect 27615 -46238 27935 -46210
rect 27615 -46542 27623 -46238
rect 27927 -46542 27935 -46238
rect 27615 -46550 27935 -46542
rect 28615 -46238 28935 -46210
rect 28615 -46542 28623 -46238
rect 28927 -46542 28935 -46238
rect 28615 -46550 28935 -46542
rect 29615 -46238 29935 -46210
rect 29615 -46542 29623 -46238
rect 29927 -46542 29935 -46238
rect 29615 -46550 29935 -46542
rect 30615 -46238 30935 -46210
rect 30615 -46542 30623 -46238
rect 30927 -46542 30935 -46238
rect 30615 -46550 30935 -46542
rect 31615 -46238 31935 -46210
rect 31615 -46542 31623 -46238
rect 31927 -46542 31935 -46238
rect 31615 -46550 31935 -46542
rect 32615 -46238 32935 -46210
rect 32615 -46542 32623 -46238
rect 32927 -46542 32935 -46238
rect 32615 -46550 32935 -46542
rect 33615 -46238 33935 -46210
rect 33615 -46542 33623 -46238
rect 33927 -46542 33935 -46238
rect 33615 -46550 33935 -46542
<< via4 >>
rect -74443 38272 -74207 38508
rect -73443 38272 -73207 38508
rect -72443 38272 -72207 38508
rect -71443 38272 -71207 38508
rect -70443 38272 -70207 38508
rect -69443 38272 -69207 38508
rect -68443 38272 -68207 38508
rect -67443 38272 -67207 38508
rect -66443 38272 -66207 38508
rect -65443 38272 -65207 38508
rect -64443 38272 -64207 38508
rect -63443 38272 -63207 38508
rect -62443 38272 -62207 38508
rect -61443 38272 -61207 38508
rect -60443 38272 -60207 38508
rect -59443 38272 -59207 38508
rect 10036 38272 10272 38508
rect 11036 38272 11272 38508
rect 12036 38272 12272 38508
rect 13036 38272 13272 38508
rect 14036 38272 14272 38508
rect 15036 38272 15272 38508
rect 16036 38272 16272 38508
rect 17036 38272 17272 38508
rect 18036 38272 18272 38508
rect 19036 38272 19272 38508
rect 20036 38272 20272 38508
rect 21036 38272 21272 38508
rect 22036 38272 22272 38508
rect 23036 38272 23272 38508
rect 24036 38272 24272 38508
rect 25036 38272 25272 38508
rect 26036 38272 26272 38508
rect 27036 38272 27272 38508
rect 28036 38272 28272 38508
rect 29036 38272 29272 38508
rect 30036 38272 30272 38508
rect 31036 38272 31272 38508
rect 32036 38272 32272 38508
rect 33036 38272 33272 38508
rect 34036 38272 34272 38508
rect -74783 37932 -74547 38168
rect -74443 37932 -74207 38168
rect -74103 37932 -73867 38168
rect -73783 37932 -73547 38168
rect -73443 37932 -73207 38168
rect -73103 37932 -72867 38168
rect -72783 37932 -72547 38168
rect -72443 37932 -72207 38168
rect -72103 37932 -71867 38168
rect -71783 37932 -71547 38168
rect -71443 37932 -71207 38168
rect -71103 37932 -70867 38168
rect -70783 37932 -70547 38168
rect -70443 37932 -70207 38168
rect -70103 37932 -69867 38168
rect -69783 37932 -69547 38168
rect -69443 37932 -69207 38168
rect -69103 37932 -68867 38168
rect -68783 37932 -68547 38168
rect -68443 37932 -68207 38168
rect -68103 37932 -67867 38168
rect -67783 37932 -67547 38168
rect -67443 37932 -67207 38168
rect -67103 37932 -66867 38168
rect -66783 37932 -66547 38168
rect -66443 37932 -66207 38168
rect -66103 37932 -65867 38168
rect -65783 37932 -65547 38168
rect -65443 37932 -65207 38168
rect -65103 37932 -64867 38168
rect -64783 37932 -64547 38168
rect -64443 37932 -64207 38168
rect -64103 37932 -63867 38168
rect -63783 37932 -63547 38168
rect -63443 37932 -63207 38168
rect -63103 37932 -62867 38168
rect -62783 37932 -62547 38168
rect -62443 37932 -62207 38168
rect -62103 37932 -61867 38168
rect -61783 37932 -61547 38168
rect -61443 37932 -61207 38168
rect -61103 37932 -60867 38168
rect -60783 37932 -60547 38168
rect -60443 37932 -60207 38168
rect -60103 37932 -59867 38168
rect -59783 37932 -59547 38168
rect -59443 37932 -59207 38168
rect -59103 37932 -58867 38168
rect 9696 37932 9932 38168
rect 10036 37932 10272 38168
rect 10376 37932 10612 38168
rect 10696 37932 10932 38168
rect 11036 37932 11272 38168
rect 11376 37932 11612 38168
rect 11696 37932 11932 38168
rect 12036 37932 12272 38168
rect 12376 37932 12612 38168
rect 12696 37932 12932 38168
rect 13036 37932 13272 38168
rect 13376 37932 13612 38168
rect 13696 37932 13932 38168
rect 14036 37932 14272 38168
rect 14376 37932 14612 38168
rect 14696 37932 14932 38168
rect 15036 37932 15272 38168
rect 15376 37932 15612 38168
rect 15696 37932 15932 38168
rect 16036 37932 16272 38168
rect 16376 37932 16612 38168
rect 16696 37932 16932 38168
rect 17036 37932 17272 38168
rect 17376 37932 17612 38168
rect 17696 37932 17932 38168
rect 18036 37932 18272 38168
rect 18376 37932 18612 38168
rect 18696 37932 18932 38168
rect 19036 37932 19272 38168
rect 19376 37932 19612 38168
rect 19696 37932 19932 38168
rect 20036 37932 20272 38168
rect 20376 37932 20612 38168
rect 20696 37932 20932 38168
rect 21036 37932 21272 38168
rect 21376 37932 21612 38168
rect 21696 37932 21932 38168
rect 22036 37932 22272 38168
rect 22376 37932 22612 38168
rect 22696 37932 22932 38168
rect 23036 37932 23272 38168
rect 23376 37932 23612 38168
rect 23696 37932 23932 38168
rect 24036 37932 24272 38168
rect 24376 37932 24612 38168
rect 24696 37932 24932 38168
rect 25036 37932 25272 38168
rect 25376 37932 25612 38168
rect 25696 37932 25932 38168
rect 26036 37932 26272 38168
rect 26376 37932 26612 38168
rect 26696 37932 26932 38168
rect 27036 37932 27272 38168
rect 27376 37932 27612 38168
rect 27696 37932 27932 38168
rect 28036 37932 28272 38168
rect 28376 37932 28612 38168
rect 28696 37932 28932 38168
rect 29036 37932 29272 38168
rect 29376 37932 29612 38168
rect 29696 37932 29932 38168
rect 30036 37932 30272 38168
rect 30376 37932 30612 38168
rect 30696 37932 30932 38168
rect 31036 37932 31272 38168
rect 31376 37932 31612 38168
rect 31696 37932 31932 38168
rect 32036 37932 32272 38168
rect 32376 37932 32612 38168
rect 32696 37932 32932 38168
rect 33036 37932 33272 38168
rect 33376 37932 33612 38168
rect 33696 37932 33932 38168
rect 34036 37932 34272 38168
rect 34376 37932 34612 38168
rect -74443 37592 -74207 37828
rect -74443 37272 -74207 37508
rect -73443 37592 -73207 37828
rect -73443 37272 -73207 37508
rect -72443 37592 -72207 37828
rect -72443 37272 -72207 37508
rect -71443 37592 -71207 37828
rect -71443 37272 -71207 37508
rect -70443 37592 -70207 37828
rect -70443 37272 -70207 37508
rect -69443 37592 -69207 37828
rect -69443 37272 -69207 37508
rect -68443 37592 -68207 37828
rect -68443 37272 -68207 37508
rect -67443 37592 -67207 37828
rect -67443 37272 -67207 37508
rect -66443 37592 -66207 37828
rect -66443 37272 -66207 37508
rect -65443 37592 -65207 37828
rect -65443 37272 -65207 37508
rect -64443 37592 -64207 37828
rect -64443 37272 -64207 37508
rect -63443 37592 -63207 37828
rect -63443 37272 -63207 37508
rect -62443 37592 -62207 37828
rect -62443 37272 -62207 37508
rect -61443 37592 -61207 37828
rect -61443 37272 -61207 37508
rect -60443 37592 -60207 37828
rect -60443 37272 -60207 37508
rect -59443 37592 -59207 37828
rect -59443 37272 -59207 37508
rect 10036 37592 10272 37828
rect 10036 37272 10272 37508
rect 11036 37592 11272 37828
rect 11036 37272 11272 37508
rect 12036 37592 12272 37828
rect 12036 37272 12272 37508
rect 13036 37592 13272 37828
rect 13036 37272 13272 37508
rect 14036 37592 14272 37828
rect 14036 37272 14272 37508
rect 15036 37592 15272 37828
rect 15036 37272 15272 37508
rect 16036 37592 16272 37828
rect 16036 37272 16272 37508
rect 17036 37592 17272 37828
rect 17036 37272 17272 37508
rect 18036 37592 18272 37828
rect 18036 37272 18272 37508
rect 19036 37592 19272 37828
rect 19036 37272 19272 37508
rect 20036 37592 20272 37828
rect 20036 37272 20272 37508
rect 21036 37592 21272 37828
rect 21036 37272 21272 37508
rect 22036 37592 22272 37828
rect 22036 37272 22272 37508
rect 23036 37592 23272 37828
rect 23036 37272 23272 37508
rect 24036 37592 24272 37828
rect 24036 37272 24272 37508
rect 25036 37592 25272 37828
rect 25036 37272 25272 37508
rect 26036 37592 26272 37828
rect 26036 37272 26272 37508
rect 27036 37592 27272 37828
rect 27036 37272 27272 37508
rect 28036 37592 28272 37828
rect 28036 37272 28272 37508
rect 29036 37592 29272 37828
rect 29036 37272 29272 37508
rect 30036 37592 30272 37828
rect 30036 37272 30272 37508
rect 31036 37592 31272 37828
rect 31036 37272 31272 37508
rect 32036 37592 32272 37828
rect 32036 37272 32272 37508
rect 33036 37592 33272 37828
rect 33036 37272 33272 37508
rect 34036 37592 34272 37828
rect 34036 37272 34272 37508
rect -74783 36932 -74547 37168
rect -74443 36932 -74207 37168
rect -74103 36932 -73867 37168
rect -73783 36932 -73547 37168
rect -73443 36932 -73207 37168
rect -73103 36932 -72867 37168
rect -72783 36932 -72547 37168
rect -72443 36932 -72207 37168
rect -72103 36932 -71867 37168
rect -71783 36932 -71547 37168
rect -71443 36932 -71207 37168
rect -71103 36932 -70867 37168
rect -70783 36932 -70547 37168
rect -70443 36932 -70207 37168
rect -70103 36932 -69867 37168
rect -69783 36932 -69547 37168
rect -69443 36932 -69207 37168
rect -69103 36932 -68867 37168
rect -68783 36932 -68547 37168
rect -68443 36932 -68207 37168
rect -68103 36932 -67867 37168
rect -67783 36932 -67547 37168
rect -67443 36932 -67207 37168
rect -67103 36932 -66867 37168
rect -66783 36932 -66547 37168
rect -66443 36932 -66207 37168
rect -66103 36932 -65867 37168
rect -65783 36932 -65547 37168
rect -65443 36932 -65207 37168
rect -65103 36932 -64867 37168
rect -64783 36932 -64547 37168
rect -64443 36932 -64207 37168
rect -64103 36932 -63867 37168
rect -63783 36932 -63547 37168
rect -63443 36932 -63207 37168
rect -63103 36932 -62867 37168
rect -62783 36932 -62547 37168
rect -62443 36932 -62207 37168
rect -62103 36932 -61867 37168
rect -61783 36932 -61547 37168
rect -61443 36932 -61207 37168
rect -61103 36932 -60867 37168
rect -60783 36932 -60547 37168
rect -60443 36932 -60207 37168
rect -60103 36932 -59867 37168
rect -59783 36932 -59547 37168
rect -59443 36932 -59207 37168
rect -59103 36932 -58867 37168
rect 9696 36932 9932 37168
rect 10036 36932 10272 37168
rect 10376 36932 10612 37168
rect 10696 36932 10932 37168
rect 11036 36932 11272 37168
rect 11376 36932 11612 37168
rect 11696 36932 11932 37168
rect 12036 36932 12272 37168
rect 12376 36932 12612 37168
rect 12696 36932 12932 37168
rect 13036 36932 13272 37168
rect 13376 36932 13612 37168
rect 13696 36932 13932 37168
rect 14036 36932 14272 37168
rect 14376 36932 14612 37168
rect 14696 36932 14932 37168
rect 15036 36932 15272 37168
rect 15376 36932 15612 37168
rect 15696 36932 15932 37168
rect 16036 36932 16272 37168
rect 16376 36932 16612 37168
rect 16696 36932 16932 37168
rect 17036 36932 17272 37168
rect 17376 36932 17612 37168
rect 17696 36932 17932 37168
rect 18036 36932 18272 37168
rect 18376 36932 18612 37168
rect 18696 36932 18932 37168
rect 19036 36932 19272 37168
rect 19376 36932 19612 37168
rect 19696 36932 19932 37168
rect 20036 36932 20272 37168
rect 20376 36932 20612 37168
rect 20696 36932 20932 37168
rect 21036 36932 21272 37168
rect 21376 36932 21612 37168
rect 21696 36932 21932 37168
rect 22036 36932 22272 37168
rect 22376 36932 22612 37168
rect 22696 36932 22932 37168
rect 23036 36932 23272 37168
rect 23376 36932 23612 37168
rect 23696 36932 23932 37168
rect 24036 36932 24272 37168
rect 24376 36932 24612 37168
rect 24696 36932 24932 37168
rect 25036 36932 25272 37168
rect 25376 36932 25612 37168
rect 25696 36932 25932 37168
rect 26036 36932 26272 37168
rect 26376 36932 26612 37168
rect 26696 36932 26932 37168
rect 27036 36932 27272 37168
rect 27376 36932 27612 37168
rect 27696 36932 27932 37168
rect 28036 36932 28272 37168
rect 28376 36932 28612 37168
rect 28696 36932 28932 37168
rect 29036 36932 29272 37168
rect 29376 36932 29612 37168
rect 29696 36932 29932 37168
rect 30036 36932 30272 37168
rect 30376 36932 30612 37168
rect 30696 36932 30932 37168
rect 31036 36932 31272 37168
rect 31376 36932 31612 37168
rect 31696 36932 31932 37168
rect 32036 36932 32272 37168
rect 32376 36932 32612 37168
rect 32696 36932 32932 37168
rect 33036 36932 33272 37168
rect 33376 36932 33612 37168
rect 33696 36932 33932 37168
rect 34036 36932 34272 37168
rect 34376 36932 34612 37168
rect -74443 36592 -74207 36828
rect -74443 36272 -74207 36508
rect -73443 36592 -73207 36828
rect -73443 36272 -73207 36508
rect -72443 36592 -72207 36828
rect -72443 36272 -72207 36508
rect -71443 36592 -71207 36828
rect -71443 36272 -71207 36508
rect -70443 36592 -70207 36828
rect -70443 36272 -70207 36508
rect -69443 36592 -69207 36828
rect -69443 36272 -69207 36508
rect -68443 36592 -68207 36828
rect -68443 36272 -68207 36508
rect -67443 36592 -67207 36828
rect -67443 36272 -67207 36508
rect -66443 36592 -66207 36828
rect -66443 36272 -66207 36508
rect -65443 36592 -65207 36828
rect -65443 36272 -65207 36508
rect -64443 36592 -64207 36828
rect -64443 36272 -64207 36508
rect -63443 36592 -63207 36828
rect -63443 36272 -63207 36508
rect -62443 36592 -62207 36828
rect -62443 36272 -62207 36508
rect -61443 36592 -61207 36828
rect -61443 36272 -61207 36508
rect -60443 36592 -60207 36828
rect -60443 36272 -60207 36508
rect -59443 36592 -59207 36828
rect -59443 36272 -59207 36508
rect 10036 36592 10272 36828
rect 10036 36272 10272 36508
rect 11036 36592 11272 36828
rect 11036 36272 11272 36508
rect 12036 36592 12272 36828
rect 12036 36272 12272 36508
rect 13036 36592 13272 36828
rect 13036 36272 13272 36508
rect 14036 36592 14272 36828
rect 14036 36272 14272 36508
rect 15036 36592 15272 36828
rect 15036 36272 15272 36508
rect 16036 36592 16272 36828
rect 16036 36272 16272 36508
rect 17036 36592 17272 36828
rect 17036 36272 17272 36508
rect 18036 36592 18272 36828
rect 18036 36272 18272 36508
rect 19036 36592 19272 36828
rect 19036 36272 19272 36508
rect 20036 36592 20272 36828
rect 20036 36272 20272 36508
rect 21036 36592 21272 36828
rect 21036 36272 21272 36508
rect 22036 36592 22272 36828
rect 22036 36272 22272 36508
rect 23036 36592 23272 36828
rect 23036 36272 23272 36508
rect 24036 36592 24272 36828
rect 24036 36272 24272 36508
rect 25036 36592 25272 36828
rect 25036 36272 25272 36508
rect 26036 36592 26272 36828
rect 26036 36272 26272 36508
rect 27036 36592 27272 36828
rect 27036 36272 27272 36508
rect 28036 36592 28272 36828
rect 28036 36272 28272 36508
rect 29036 36592 29272 36828
rect 29036 36272 29272 36508
rect 30036 36592 30272 36828
rect 30036 36272 30272 36508
rect 31036 36592 31272 36828
rect 31036 36272 31272 36508
rect 32036 36592 32272 36828
rect 32036 36272 32272 36508
rect 33036 36592 33272 36828
rect 33036 36272 33272 36508
rect 34036 36592 34272 36828
rect 34036 36272 34272 36508
rect -74783 35932 -74547 36168
rect -74443 35932 -74207 36168
rect -74103 35932 -73867 36168
rect -73783 35932 -73547 36168
rect -73443 35932 -73207 36168
rect -73103 35932 -72867 36168
rect -72783 35932 -72547 36168
rect -72443 35932 -72207 36168
rect -72103 35932 -71867 36168
rect -71783 35932 -71547 36168
rect -71443 35932 -71207 36168
rect -71103 35932 -70867 36168
rect -70783 35932 -70547 36168
rect -70443 35932 -70207 36168
rect -70103 35932 -69867 36168
rect -69783 35932 -69547 36168
rect -69443 35932 -69207 36168
rect -69103 35932 -68867 36168
rect -68783 35932 -68547 36168
rect -68443 35932 -68207 36168
rect -68103 35932 -67867 36168
rect -67783 35932 -67547 36168
rect -67443 35932 -67207 36168
rect -67103 35932 -66867 36168
rect -66783 35932 -66547 36168
rect -66443 35932 -66207 36168
rect -66103 35932 -65867 36168
rect -65783 35932 -65547 36168
rect -65443 35932 -65207 36168
rect -65103 35932 -64867 36168
rect -64783 35932 -64547 36168
rect -64443 35932 -64207 36168
rect -64103 35932 -63867 36168
rect -63783 35932 -63547 36168
rect -63443 35932 -63207 36168
rect -63103 35932 -62867 36168
rect -62783 35932 -62547 36168
rect -62443 35932 -62207 36168
rect -62103 35932 -61867 36168
rect -61783 35932 -61547 36168
rect -61443 35932 -61207 36168
rect -61103 35932 -60867 36168
rect -60783 35932 -60547 36168
rect -60443 35932 -60207 36168
rect -60103 35932 -59867 36168
rect -59783 35932 -59547 36168
rect -59443 35932 -59207 36168
rect -59103 35932 -58867 36168
rect 9696 35932 9932 36168
rect 10036 35932 10272 36168
rect 10376 35932 10612 36168
rect 10696 35932 10932 36168
rect 11036 35932 11272 36168
rect 11376 35932 11612 36168
rect 11696 35932 11932 36168
rect 12036 35932 12272 36168
rect 12376 35932 12612 36168
rect 12696 35932 12932 36168
rect 13036 35932 13272 36168
rect 13376 35932 13612 36168
rect 13696 35932 13932 36168
rect 14036 35932 14272 36168
rect 14376 35932 14612 36168
rect 14696 35932 14932 36168
rect 15036 35932 15272 36168
rect 15376 35932 15612 36168
rect 15696 35932 15932 36168
rect 16036 35932 16272 36168
rect 16376 35932 16612 36168
rect 16696 35932 16932 36168
rect 17036 35932 17272 36168
rect 17376 35932 17612 36168
rect 17696 35932 17932 36168
rect 18036 35932 18272 36168
rect 18376 35932 18612 36168
rect 18696 35932 18932 36168
rect 19036 35932 19272 36168
rect 19376 35932 19612 36168
rect 19696 35932 19932 36168
rect 20036 35932 20272 36168
rect 20376 35932 20612 36168
rect 20696 35932 20932 36168
rect 21036 35932 21272 36168
rect 21376 35932 21612 36168
rect 21696 35932 21932 36168
rect 22036 35932 22272 36168
rect 22376 35932 22612 36168
rect 22696 35932 22932 36168
rect 23036 35932 23272 36168
rect 23376 35932 23612 36168
rect 23696 35932 23932 36168
rect 24036 35932 24272 36168
rect 24376 35932 24612 36168
rect 24696 35932 24932 36168
rect 25036 35932 25272 36168
rect 25376 35932 25612 36168
rect 25696 35932 25932 36168
rect 26036 35932 26272 36168
rect 26376 35932 26612 36168
rect 26696 35932 26932 36168
rect 27036 35932 27272 36168
rect 27376 35932 27612 36168
rect 27696 35932 27932 36168
rect 28036 35932 28272 36168
rect 28376 35932 28612 36168
rect 28696 35932 28932 36168
rect 29036 35932 29272 36168
rect 29376 35932 29612 36168
rect 29696 35932 29932 36168
rect 30036 35932 30272 36168
rect 30376 35932 30612 36168
rect 30696 35932 30932 36168
rect 31036 35932 31272 36168
rect 31376 35932 31612 36168
rect 31696 35932 31932 36168
rect 32036 35932 32272 36168
rect 32376 35932 32612 36168
rect 32696 35932 32932 36168
rect 33036 35932 33272 36168
rect 33376 35932 33612 36168
rect 33696 35932 33932 36168
rect 34036 35932 34272 36168
rect 34376 35932 34612 36168
rect -74443 35592 -74207 35828
rect -74443 35272 -74207 35508
rect -73443 35592 -73207 35828
rect -73443 35272 -73207 35508
rect -72443 35592 -72207 35828
rect -72443 35272 -72207 35508
rect -71443 35592 -71207 35828
rect -71443 35272 -71207 35508
rect -70443 35592 -70207 35828
rect -70443 35272 -70207 35508
rect -69443 35592 -69207 35828
rect -69443 35272 -69207 35508
rect -68443 35592 -68207 35828
rect -68443 35272 -68207 35508
rect -67443 35592 -67207 35828
rect -67443 35272 -67207 35508
rect -66443 35592 -66207 35828
rect -66443 35272 -66207 35508
rect -65443 35592 -65207 35828
rect -65443 35272 -65207 35508
rect -64443 35592 -64207 35828
rect -64443 35272 -64207 35508
rect -63443 35592 -63207 35828
rect -63443 35272 -63207 35508
rect -62443 35592 -62207 35828
rect -62443 35272 -62207 35508
rect -61443 35592 -61207 35828
rect -61443 35272 -61207 35508
rect -60443 35592 -60207 35828
rect -60443 35272 -60207 35508
rect -59443 35592 -59207 35828
rect -59443 35272 -59207 35508
rect 10036 35592 10272 35828
rect 10036 35272 10272 35508
rect 11036 35592 11272 35828
rect 11036 35272 11272 35508
rect 12036 35592 12272 35828
rect 12036 35272 12272 35508
rect 13036 35592 13272 35828
rect 13036 35272 13272 35508
rect 14036 35592 14272 35828
rect 14036 35272 14272 35508
rect 15036 35592 15272 35828
rect 15036 35272 15272 35508
rect 16036 35592 16272 35828
rect 16036 35272 16272 35508
rect 17036 35592 17272 35828
rect 17036 35272 17272 35508
rect 18036 35592 18272 35828
rect 18036 35272 18272 35508
rect 19036 35592 19272 35828
rect 19036 35272 19272 35508
rect 20036 35592 20272 35828
rect 20036 35272 20272 35508
rect 21036 35592 21272 35828
rect 21036 35272 21272 35508
rect 22036 35592 22272 35828
rect 22036 35272 22272 35508
rect 23036 35592 23272 35828
rect 23036 35272 23272 35508
rect 24036 35592 24272 35828
rect 24036 35272 24272 35508
rect 25036 35592 25272 35828
rect 25036 35272 25272 35508
rect 26036 35592 26272 35828
rect 26036 35272 26272 35508
rect 27036 35592 27272 35828
rect 27036 35272 27272 35508
rect 28036 35592 28272 35828
rect 28036 35272 28272 35508
rect 29036 35592 29272 35828
rect 29036 35272 29272 35508
rect 30036 35592 30272 35828
rect 30036 35272 30272 35508
rect 31036 35592 31272 35828
rect 31036 35272 31272 35508
rect 32036 35592 32272 35828
rect 32036 35272 32272 35508
rect 33036 35592 33272 35828
rect 33036 35272 33272 35508
rect 34036 35592 34272 35828
rect 34036 35272 34272 35508
rect -74783 34932 -74547 35168
rect -74443 34932 -74207 35168
rect -74103 34932 -73867 35168
rect -73783 34932 -73547 35168
rect -73443 34932 -73207 35168
rect -73103 34932 -72867 35168
rect -72783 34932 -72547 35168
rect -72443 34932 -72207 35168
rect -72103 34932 -71867 35168
rect -71783 34932 -71547 35168
rect -71443 34932 -71207 35168
rect -71103 34932 -70867 35168
rect -70783 34932 -70547 35168
rect -70443 34932 -70207 35168
rect -70103 34932 -69867 35168
rect -69783 34932 -69547 35168
rect -69443 34932 -69207 35168
rect -69103 34932 -68867 35168
rect -68783 34932 -68547 35168
rect -68443 34932 -68207 35168
rect -68103 34932 -67867 35168
rect -67783 34932 -67547 35168
rect -67443 34932 -67207 35168
rect -67103 34932 -66867 35168
rect -66783 34932 -66547 35168
rect -66443 34932 -66207 35168
rect -66103 34932 -65867 35168
rect -65783 34932 -65547 35168
rect -65443 34932 -65207 35168
rect -65103 34932 -64867 35168
rect -64783 34932 -64547 35168
rect -64443 34932 -64207 35168
rect -64103 34932 -63867 35168
rect -63783 34932 -63547 35168
rect -63443 34932 -63207 35168
rect -63103 34932 -62867 35168
rect -62783 34932 -62547 35168
rect -62443 34932 -62207 35168
rect -62103 34932 -61867 35168
rect -61783 34932 -61547 35168
rect -61443 34932 -61207 35168
rect -61103 34932 -60867 35168
rect -60783 34932 -60547 35168
rect -60443 34932 -60207 35168
rect -60103 34932 -59867 35168
rect -59783 34932 -59547 35168
rect -59443 34932 -59207 35168
rect -59103 34932 -58867 35168
rect 9696 34932 9932 35168
rect 10036 34932 10272 35168
rect 10376 34932 10612 35168
rect 10696 34932 10932 35168
rect 11036 34932 11272 35168
rect 11376 34932 11612 35168
rect 11696 34932 11932 35168
rect 12036 34932 12272 35168
rect 12376 34932 12612 35168
rect 12696 34932 12932 35168
rect 13036 34932 13272 35168
rect 13376 34932 13612 35168
rect 13696 34932 13932 35168
rect 14036 34932 14272 35168
rect 14376 34932 14612 35168
rect 14696 34932 14932 35168
rect 15036 34932 15272 35168
rect 15376 34932 15612 35168
rect 15696 34932 15932 35168
rect 16036 34932 16272 35168
rect 16376 34932 16612 35168
rect 16696 34932 16932 35168
rect 17036 34932 17272 35168
rect 17376 34932 17612 35168
rect 17696 34932 17932 35168
rect 18036 34932 18272 35168
rect 18376 34932 18612 35168
rect 18696 34932 18932 35168
rect 19036 34932 19272 35168
rect 19376 34932 19612 35168
rect 19696 34932 19932 35168
rect 20036 34932 20272 35168
rect 20376 34932 20612 35168
rect 20696 34932 20932 35168
rect 21036 34932 21272 35168
rect 21376 34932 21612 35168
rect 21696 34932 21932 35168
rect 22036 34932 22272 35168
rect 22376 34932 22612 35168
rect 22696 34932 22932 35168
rect 23036 34932 23272 35168
rect 23376 34932 23612 35168
rect 23696 34932 23932 35168
rect 24036 34932 24272 35168
rect 24376 34932 24612 35168
rect 24696 34932 24932 35168
rect 25036 34932 25272 35168
rect 25376 34932 25612 35168
rect 25696 34932 25932 35168
rect 26036 34932 26272 35168
rect 26376 34932 26612 35168
rect 26696 34932 26932 35168
rect 27036 34932 27272 35168
rect 27376 34932 27612 35168
rect 27696 34932 27932 35168
rect 28036 34932 28272 35168
rect 28376 34932 28612 35168
rect 28696 34932 28932 35168
rect 29036 34932 29272 35168
rect 29376 34932 29612 35168
rect 29696 34932 29932 35168
rect 30036 34932 30272 35168
rect 30376 34932 30612 35168
rect 30696 34932 30932 35168
rect 31036 34932 31272 35168
rect 31376 34932 31612 35168
rect 31696 34932 31932 35168
rect 32036 34932 32272 35168
rect 32376 34932 32612 35168
rect 32696 34932 32932 35168
rect 33036 34932 33272 35168
rect 33376 34932 33612 35168
rect 33696 34932 33932 35168
rect 34036 34932 34272 35168
rect 34376 34932 34612 35168
rect -74443 34592 -74207 34828
rect -74443 34272 -74207 34508
rect -73443 34592 -73207 34828
rect -73443 34272 -73207 34508
rect -72443 34592 -72207 34828
rect -72443 34272 -72207 34508
rect -71443 34592 -71207 34828
rect -71443 34272 -71207 34508
rect -70443 34592 -70207 34828
rect -70443 34272 -70207 34508
rect -69443 34592 -69207 34828
rect -69443 34272 -69207 34508
rect -68443 34592 -68207 34828
rect -68443 34272 -68207 34508
rect -67443 34592 -67207 34828
rect -67443 34272 -67207 34508
rect -66443 34592 -66207 34828
rect -66443 34272 -66207 34508
rect -65443 34592 -65207 34828
rect -65443 34272 -65207 34508
rect -64443 34592 -64207 34828
rect -64443 34272 -64207 34508
rect -63443 34592 -63207 34828
rect -63443 34272 -63207 34508
rect -62443 34592 -62207 34828
rect -62443 34272 -62207 34508
rect -61443 34592 -61207 34828
rect -61443 34272 -61207 34508
rect -60443 34592 -60207 34828
rect -60443 34272 -60207 34508
rect -59443 34592 -59207 34828
rect -59443 34272 -59207 34508
rect 10036 34592 10272 34828
rect 10036 34272 10272 34508
rect 11036 34592 11272 34828
rect 11036 34272 11272 34508
rect 12036 34592 12272 34828
rect 12036 34272 12272 34508
rect 13036 34592 13272 34828
rect 13036 34272 13272 34508
rect 14036 34592 14272 34828
rect 14036 34272 14272 34508
rect 15036 34592 15272 34828
rect 15036 34272 15272 34508
rect 16036 34592 16272 34828
rect 16036 34272 16272 34508
rect 17036 34592 17272 34828
rect 17036 34272 17272 34508
rect 18036 34592 18272 34828
rect 18036 34272 18272 34508
rect 19036 34592 19272 34828
rect 19036 34272 19272 34508
rect 20036 34592 20272 34828
rect 20036 34272 20272 34508
rect 21036 34592 21272 34828
rect 21036 34272 21272 34508
rect 22036 34592 22272 34828
rect 22036 34272 22272 34508
rect 23036 34592 23272 34828
rect 23036 34272 23272 34508
rect 24036 34592 24272 34828
rect 24036 34272 24272 34508
rect 25036 34592 25272 34828
rect 25036 34272 25272 34508
rect 26036 34592 26272 34828
rect 26036 34272 26272 34508
rect 27036 34592 27272 34828
rect 27036 34272 27272 34508
rect 28036 34592 28272 34828
rect 28036 34272 28272 34508
rect 29036 34592 29272 34828
rect 29036 34272 29272 34508
rect 30036 34592 30272 34828
rect 30036 34272 30272 34508
rect 31036 34592 31272 34828
rect 31036 34272 31272 34508
rect 32036 34592 32272 34828
rect 32036 34272 32272 34508
rect 33036 34592 33272 34828
rect 33036 34272 33272 34508
rect 34036 34592 34272 34828
rect 34036 34272 34272 34508
rect -74783 33932 -74547 34168
rect -74443 33932 -74207 34168
rect -74103 33932 -73867 34168
rect -73783 33932 -73547 34168
rect -73443 33932 -73207 34168
rect -73103 33932 -72867 34168
rect -72783 33932 -72547 34168
rect -72443 33932 -72207 34168
rect -72103 33932 -71867 34168
rect -71783 33932 -71547 34168
rect -71443 33932 -71207 34168
rect -71103 33932 -70867 34168
rect -70783 33932 -70547 34168
rect -70443 33932 -70207 34168
rect -70103 33932 -69867 34168
rect -69783 33932 -69547 34168
rect -69443 33932 -69207 34168
rect -69103 33932 -68867 34168
rect -68783 33932 -68547 34168
rect -68443 33932 -68207 34168
rect -68103 33932 -67867 34168
rect -67783 33932 -67547 34168
rect -67443 33932 -67207 34168
rect -67103 33932 -66867 34168
rect -66783 33932 -66547 34168
rect -66443 33932 -66207 34168
rect -66103 33932 -65867 34168
rect -65783 33932 -65547 34168
rect -65443 33932 -65207 34168
rect -65103 33932 -64867 34168
rect -64783 33932 -64547 34168
rect -64443 33932 -64207 34168
rect -64103 33932 -63867 34168
rect -63783 33932 -63547 34168
rect -63443 33932 -63207 34168
rect -63103 33932 -62867 34168
rect -62783 33932 -62547 34168
rect -62443 33932 -62207 34168
rect -62103 33932 -61867 34168
rect -61783 33932 -61547 34168
rect -61443 33932 -61207 34168
rect -61103 33932 -60867 34168
rect -60783 33932 -60547 34168
rect -60443 33932 -60207 34168
rect -60103 33932 -59867 34168
rect -59783 33932 -59547 34168
rect -59443 33932 -59207 34168
rect -59103 33932 -58867 34168
rect 9696 33932 9932 34168
rect 10036 33932 10272 34168
rect 10376 33932 10612 34168
rect 10696 33932 10932 34168
rect 11036 33932 11272 34168
rect 11376 33932 11612 34168
rect 11696 33932 11932 34168
rect 12036 33932 12272 34168
rect 12376 33932 12612 34168
rect 12696 33932 12932 34168
rect 13036 33932 13272 34168
rect 13376 33932 13612 34168
rect 13696 33932 13932 34168
rect 14036 33932 14272 34168
rect 14376 33932 14612 34168
rect 14696 33932 14932 34168
rect 15036 33932 15272 34168
rect 15376 33932 15612 34168
rect 15696 33932 15932 34168
rect 16036 33932 16272 34168
rect 16376 33932 16612 34168
rect 16696 33932 16932 34168
rect 17036 33932 17272 34168
rect 17376 33932 17612 34168
rect 17696 33932 17932 34168
rect 18036 33932 18272 34168
rect 18376 33932 18612 34168
rect 18696 33932 18932 34168
rect 19036 33932 19272 34168
rect 19376 33932 19612 34168
rect 19696 33932 19932 34168
rect 20036 33932 20272 34168
rect 20376 33932 20612 34168
rect 20696 33932 20932 34168
rect 21036 33932 21272 34168
rect 21376 33932 21612 34168
rect 21696 33932 21932 34168
rect 22036 33932 22272 34168
rect 22376 33932 22612 34168
rect 22696 33932 22932 34168
rect 23036 33932 23272 34168
rect 23376 33932 23612 34168
rect 23696 33932 23932 34168
rect 24036 33932 24272 34168
rect 24376 33932 24612 34168
rect 24696 33932 24932 34168
rect 25036 33932 25272 34168
rect 25376 33932 25612 34168
rect 25696 33932 25932 34168
rect 26036 33932 26272 34168
rect 26376 33932 26612 34168
rect 26696 33932 26932 34168
rect 27036 33932 27272 34168
rect 27376 33932 27612 34168
rect 27696 33932 27932 34168
rect 28036 33932 28272 34168
rect 28376 33932 28612 34168
rect 28696 33932 28932 34168
rect 29036 33932 29272 34168
rect 29376 33932 29612 34168
rect 29696 33932 29932 34168
rect 30036 33932 30272 34168
rect 30376 33932 30612 34168
rect 30696 33932 30932 34168
rect 31036 33932 31272 34168
rect 31376 33932 31612 34168
rect 31696 33932 31932 34168
rect 32036 33932 32272 34168
rect 32376 33932 32612 34168
rect 32696 33932 32932 34168
rect 33036 33932 33272 34168
rect 33376 33932 33612 34168
rect 33696 33932 33932 34168
rect 34036 33932 34272 34168
rect 34376 33932 34612 34168
rect -74443 33592 -74207 33828
rect -74443 33272 -74207 33508
rect -73443 33592 -73207 33828
rect -73443 33272 -73207 33508
rect -72443 33592 -72207 33828
rect -72443 33272 -72207 33508
rect -71443 33592 -71207 33828
rect -71443 33272 -71207 33508
rect -70443 33592 -70207 33828
rect -70443 33272 -70207 33508
rect -69443 33592 -69207 33828
rect -69443 33272 -69207 33508
rect -68443 33592 -68207 33828
rect -68443 33272 -68207 33508
rect -67443 33592 -67207 33828
rect -67443 33272 -67207 33508
rect -66443 33592 -66207 33828
rect -66443 33272 -66207 33508
rect -65443 33592 -65207 33828
rect -65443 33272 -65207 33508
rect -64443 33592 -64207 33828
rect -64443 33272 -64207 33508
rect -63443 33592 -63207 33828
rect -63443 33272 -63207 33508
rect -62443 33592 -62207 33828
rect -62443 33272 -62207 33508
rect -61443 33592 -61207 33828
rect -61443 33272 -61207 33508
rect -60443 33592 -60207 33828
rect -60443 33272 -60207 33508
rect -59443 33592 -59207 33828
rect -59443 33272 -59207 33508
rect 10036 33592 10272 33828
rect 10036 33272 10272 33508
rect 11036 33592 11272 33828
rect 11036 33272 11272 33508
rect 12036 33592 12272 33828
rect 12036 33272 12272 33508
rect 13036 33592 13272 33828
rect 13036 33272 13272 33508
rect 14036 33592 14272 33828
rect 14036 33272 14272 33508
rect 15036 33592 15272 33828
rect 15036 33272 15272 33508
rect 16036 33592 16272 33828
rect 16036 33272 16272 33508
rect 17036 33592 17272 33828
rect 17036 33272 17272 33508
rect 18036 33592 18272 33828
rect 18036 33272 18272 33508
rect 19036 33592 19272 33828
rect 19036 33272 19272 33508
rect 20036 33592 20272 33828
rect 20036 33272 20272 33508
rect 21036 33592 21272 33828
rect 21036 33272 21272 33508
rect 22036 33592 22272 33828
rect 22036 33272 22272 33508
rect 23036 33592 23272 33828
rect 23036 33272 23272 33508
rect 24036 33592 24272 33828
rect 24036 33272 24272 33508
rect 25036 33592 25272 33828
rect 25036 33272 25272 33508
rect 26036 33592 26272 33828
rect 26036 33272 26272 33508
rect 27036 33592 27272 33828
rect 27036 33272 27272 33508
rect 28036 33592 28272 33828
rect 28036 33272 28272 33508
rect 29036 33592 29272 33828
rect 29036 33272 29272 33508
rect 30036 33592 30272 33828
rect 30036 33272 30272 33508
rect 31036 33592 31272 33828
rect 31036 33272 31272 33508
rect 32036 33592 32272 33828
rect 32036 33272 32272 33508
rect 33036 33592 33272 33828
rect 33036 33272 33272 33508
rect 34036 33592 34272 33828
rect 34036 33272 34272 33508
rect -74783 32932 -74547 33168
rect -74443 32932 -74207 33168
rect -74103 32932 -73867 33168
rect -73783 32932 -73547 33168
rect -73443 32932 -73207 33168
rect -73103 32932 -72867 33168
rect -72783 32932 -72547 33168
rect -72443 32932 -72207 33168
rect -72103 32932 -71867 33168
rect -71783 32932 -71547 33168
rect -71443 32932 -71207 33168
rect -71103 32932 -70867 33168
rect -70783 32932 -70547 33168
rect -70443 32932 -70207 33168
rect -70103 32932 -69867 33168
rect -69783 32932 -69547 33168
rect -69443 32932 -69207 33168
rect -69103 32932 -68867 33168
rect -68783 32932 -68547 33168
rect -68443 32932 -68207 33168
rect -68103 32932 -67867 33168
rect -67783 32932 -67547 33168
rect -67443 32932 -67207 33168
rect -67103 32932 -66867 33168
rect -66783 32932 -66547 33168
rect -66443 32932 -66207 33168
rect -66103 32932 -65867 33168
rect -65783 32932 -65547 33168
rect -65443 32932 -65207 33168
rect -65103 32932 -64867 33168
rect -64783 32932 -64547 33168
rect -64443 32932 -64207 33168
rect -64103 32932 -63867 33168
rect -63783 32932 -63547 33168
rect -63443 32932 -63207 33168
rect -63103 32932 -62867 33168
rect -62783 32932 -62547 33168
rect -62443 32932 -62207 33168
rect -62103 32932 -61867 33168
rect -61783 32932 -61547 33168
rect -61443 32932 -61207 33168
rect -61103 32932 -60867 33168
rect -60783 32932 -60547 33168
rect -60443 32932 -60207 33168
rect -60103 32932 -59867 33168
rect -59783 32932 -59547 33168
rect -59443 32932 -59207 33168
rect -59103 32932 -58867 33168
rect 9696 32932 9932 33168
rect 10036 32932 10272 33168
rect 10376 32932 10612 33168
rect 10696 32932 10932 33168
rect 11036 32932 11272 33168
rect 11376 32932 11612 33168
rect 11696 32932 11932 33168
rect 12036 32932 12272 33168
rect 12376 32932 12612 33168
rect 12696 32932 12932 33168
rect 13036 32932 13272 33168
rect 13376 32932 13612 33168
rect 13696 32932 13932 33168
rect 14036 32932 14272 33168
rect 14376 32932 14612 33168
rect 14696 32932 14932 33168
rect 15036 32932 15272 33168
rect 15376 32932 15612 33168
rect 15696 32932 15932 33168
rect 16036 32932 16272 33168
rect 16376 32932 16612 33168
rect 16696 32932 16932 33168
rect 17036 32932 17272 33168
rect 17376 32932 17612 33168
rect 17696 32932 17932 33168
rect 18036 32932 18272 33168
rect 18376 32932 18612 33168
rect 18696 32932 18932 33168
rect 19036 32932 19272 33168
rect 19376 32932 19612 33168
rect 19696 32932 19932 33168
rect 20036 32932 20272 33168
rect 20376 32932 20612 33168
rect 20696 32932 20932 33168
rect 21036 32932 21272 33168
rect 21376 32932 21612 33168
rect 21696 32932 21932 33168
rect 22036 32932 22272 33168
rect 22376 32932 22612 33168
rect 22696 32932 22932 33168
rect 23036 32932 23272 33168
rect 23376 32932 23612 33168
rect 23696 32932 23932 33168
rect 24036 32932 24272 33168
rect 24376 32932 24612 33168
rect 24696 32932 24932 33168
rect 25036 32932 25272 33168
rect 25376 32932 25612 33168
rect 25696 32932 25932 33168
rect 26036 32932 26272 33168
rect 26376 32932 26612 33168
rect 26696 32932 26932 33168
rect 27036 32932 27272 33168
rect 27376 32932 27612 33168
rect 27696 32932 27932 33168
rect 28036 32932 28272 33168
rect 28376 32932 28612 33168
rect 28696 32932 28932 33168
rect 29036 32932 29272 33168
rect 29376 32932 29612 33168
rect 29696 32932 29932 33168
rect 30036 32932 30272 33168
rect 30376 32932 30612 33168
rect 30696 32932 30932 33168
rect 31036 32932 31272 33168
rect 31376 32932 31612 33168
rect 31696 32932 31932 33168
rect 32036 32932 32272 33168
rect 32376 32932 32612 33168
rect 32696 32932 32932 33168
rect 33036 32932 33272 33168
rect 33376 32932 33612 33168
rect 33696 32932 33932 33168
rect 34036 32932 34272 33168
rect 34376 32932 34612 33168
rect -74443 32592 -74207 32828
rect -74443 32272 -74207 32508
rect -73443 32592 -73207 32828
rect -73443 32272 -73207 32508
rect -72443 32592 -72207 32828
rect -72443 32272 -72207 32508
rect -71443 32592 -71207 32828
rect -71443 32272 -71207 32508
rect -70443 32592 -70207 32828
rect -70443 32272 -70207 32508
rect -69443 32592 -69207 32828
rect -69443 32272 -69207 32508
rect -68443 32592 -68207 32828
rect -68443 32272 -68207 32508
rect -67443 32592 -67207 32828
rect -67443 32272 -67207 32508
rect -66443 32592 -66207 32828
rect -66443 32272 -66207 32508
rect -65443 32592 -65207 32828
rect -65443 32272 -65207 32508
rect -64443 32592 -64207 32828
rect -64443 32272 -64207 32508
rect -63443 32592 -63207 32828
rect -63443 32272 -63207 32508
rect -62443 32592 -62207 32828
rect -62443 32272 -62207 32508
rect -61443 32592 -61207 32828
rect -61443 32272 -61207 32508
rect -60443 32592 -60207 32828
rect -60443 32272 -60207 32508
rect -59443 32592 -59207 32828
rect -59443 32272 -59207 32508
rect 10036 32592 10272 32828
rect 10036 32272 10272 32508
rect 11036 32592 11272 32828
rect 11036 32272 11272 32508
rect 12036 32592 12272 32828
rect 12036 32272 12272 32508
rect 13036 32592 13272 32828
rect 13036 32272 13272 32508
rect 14036 32592 14272 32828
rect 14036 32272 14272 32508
rect 15036 32592 15272 32828
rect 15036 32272 15272 32508
rect 16036 32592 16272 32828
rect 16036 32272 16272 32508
rect 17036 32592 17272 32828
rect 17036 32272 17272 32508
rect 18036 32592 18272 32828
rect 18036 32272 18272 32508
rect 19036 32592 19272 32828
rect 19036 32272 19272 32508
rect 20036 32592 20272 32828
rect 20036 32272 20272 32508
rect 21036 32592 21272 32828
rect 21036 32272 21272 32508
rect 22036 32592 22272 32828
rect 22036 32272 22272 32508
rect 23036 32592 23272 32828
rect 23036 32272 23272 32508
rect 24036 32592 24272 32828
rect 24036 32272 24272 32508
rect 25036 32592 25272 32828
rect 25036 32272 25272 32508
rect 26036 32592 26272 32828
rect 26036 32272 26272 32508
rect 27036 32592 27272 32828
rect 27036 32272 27272 32508
rect 28036 32592 28272 32828
rect 28036 32272 28272 32508
rect 29036 32592 29272 32828
rect 29036 32272 29272 32508
rect 30036 32592 30272 32828
rect 30036 32272 30272 32508
rect 31036 32592 31272 32828
rect 31036 32272 31272 32508
rect 32036 32592 32272 32828
rect 32036 32272 32272 32508
rect 33036 32592 33272 32828
rect 33036 32272 33272 32508
rect 34036 32592 34272 32828
rect 34036 32272 34272 32508
rect -74783 31932 -74547 32168
rect -74443 31932 -74207 32168
rect -74103 31932 -73867 32168
rect -73783 31932 -73547 32168
rect -73443 31932 -73207 32168
rect -73103 31932 -72867 32168
rect -72783 31932 -72547 32168
rect -72443 31932 -72207 32168
rect -72103 31932 -71867 32168
rect -71783 31932 -71547 32168
rect -71443 31932 -71207 32168
rect -71103 31932 -70867 32168
rect -70783 31932 -70547 32168
rect -70443 31932 -70207 32168
rect -70103 31932 -69867 32168
rect -69783 31932 -69547 32168
rect -69443 31932 -69207 32168
rect -69103 31932 -68867 32168
rect -68783 31932 -68547 32168
rect -68443 31932 -68207 32168
rect -68103 31932 -67867 32168
rect -67783 31932 -67547 32168
rect -67443 31932 -67207 32168
rect -67103 31932 -66867 32168
rect -66783 31932 -66547 32168
rect -66443 31932 -66207 32168
rect -66103 31932 -65867 32168
rect -65783 31932 -65547 32168
rect -65443 31932 -65207 32168
rect -65103 31932 -64867 32168
rect -64783 31932 -64547 32168
rect -64443 31932 -64207 32168
rect -64103 31932 -63867 32168
rect -63783 31932 -63547 32168
rect -63443 31932 -63207 32168
rect -63103 31932 -62867 32168
rect -62783 31932 -62547 32168
rect -62443 31932 -62207 32168
rect -62103 31932 -61867 32168
rect -61783 31932 -61547 32168
rect -61443 31932 -61207 32168
rect -61103 31932 -60867 32168
rect -60783 31932 -60547 32168
rect -60443 31932 -60207 32168
rect -60103 31932 -59867 32168
rect -59783 31932 -59547 32168
rect -59443 31932 -59207 32168
rect -59103 31932 -58867 32168
rect 9696 31932 9932 32168
rect 10036 31932 10272 32168
rect 10376 31932 10612 32168
rect 10696 31932 10932 32168
rect 11036 31932 11272 32168
rect 11376 31932 11612 32168
rect 11696 31932 11932 32168
rect 12036 31932 12272 32168
rect 12376 31932 12612 32168
rect 12696 31932 12932 32168
rect 13036 31932 13272 32168
rect 13376 31932 13612 32168
rect 13696 31932 13932 32168
rect 14036 31932 14272 32168
rect 14376 31932 14612 32168
rect 14696 31932 14932 32168
rect 15036 31932 15272 32168
rect 15376 31932 15612 32168
rect 15696 31932 15932 32168
rect 16036 31932 16272 32168
rect 16376 31932 16612 32168
rect 16696 31932 16932 32168
rect 17036 31932 17272 32168
rect 17376 31932 17612 32168
rect 17696 31932 17932 32168
rect 18036 31932 18272 32168
rect 18376 31932 18612 32168
rect 18696 31932 18932 32168
rect 19036 31932 19272 32168
rect 19376 31932 19612 32168
rect 19696 31932 19932 32168
rect 20036 31932 20272 32168
rect 20376 31932 20612 32168
rect 20696 31932 20932 32168
rect 21036 31932 21272 32168
rect 21376 31932 21612 32168
rect 21696 31932 21932 32168
rect 22036 31932 22272 32168
rect 22376 31932 22612 32168
rect 22696 31932 22932 32168
rect 23036 31932 23272 32168
rect 23376 31932 23612 32168
rect 23696 31932 23932 32168
rect 24036 31932 24272 32168
rect 24376 31932 24612 32168
rect 24696 31932 24932 32168
rect 25036 31932 25272 32168
rect 25376 31932 25612 32168
rect 25696 31932 25932 32168
rect 26036 31932 26272 32168
rect 26376 31932 26612 32168
rect 26696 31932 26932 32168
rect 27036 31932 27272 32168
rect 27376 31932 27612 32168
rect 27696 31932 27932 32168
rect 28036 31932 28272 32168
rect 28376 31932 28612 32168
rect 28696 31932 28932 32168
rect 29036 31932 29272 32168
rect 29376 31932 29612 32168
rect 29696 31932 29932 32168
rect 30036 31932 30272 32168
rect 30376 31932 30612 32168
rect 30696 31932 30932 32168
rect 31036 31932 31272 32168
rect 31376 31932 31612 32168
rect 31696 31932 31932 32168
rect 32036 31932 32272 32168
rect 32376 31932 32612 32168
rect 32696 31932 32932 32168
rect 33036 31932 33272 32168
rect 33376 31932 33612 32168
rect 33696 31932 33932 32168
rect 34036 31932 34272 32168
rect 34376 31932 34612 32168
rect -74443 31592 -74207 31828
rect -74443 31272 -74207 31508
rect -73443 31592 -73207 31828
rect -73443 31272 -73207 31508
rect -72443 31592 -72207 31828
rect -72443 31272 -72207 31508
rect -71443 31592 -71207 31828
rect -71443 31272 -71207 31508
rect -70443 31592 -70207 31828
rect -70443 31272 -70207 31508
rect -69443 31592 -69207 31828
rect -69443 31272 -69207 31508
rect -68443 31592 -68207 31828
rect -68443 31272 -68207 31508
rect -67443 31592 -67207 31828
rect -67443 31272 -67207 31508
rect -66443 31592 -66207 31828
rect -66443 31272 -66207 31508
rect -65443 31592 -65207 31828
rect -65443 31272 -65207 31508
rect -64443 31592 -64207 31828
rect -64443 31272 -64207 31508
rect -63443 31592 -63207 31828
rect -63443 31272 -63207 31508
rect -62443 31592 -62207 31828
rect -62443 31272 -62207 31508
rect -61443 31592 -61207 31828
rect -61443 31272 -61207 31508
rect -60443 31592 -60207 31828
rect -60443 31272 -60207 31508
rect -59443 31592 -59207 31828
rect -59443 31272 -59207 31508
rect 10036 31592 10272 31828
rect 10036 31272 10272 31508
rect 11036 31592 11272 31828
rect 11036 31272 11272 31508
rect 12036 31592 12272 31828
rect 12036 31272 12272 31508
rect 13036 31592 13272 31828
rect 13036 31272 13272 31508
rect 14036 31592 14272 31828
rect 14036 31272 14272 31508
rect 15036 31592 15272 31828
rect 15036 31272 15272 31508
rect 16036 31592 16272 31828
rect 16036 31272 16272 31508
rect 17036 31592 17272 31828
rect 17036 31272 17272 31508
rect 18036 31592 18272 31828
rect 18036 31272 18272 31508
rect 19036 31592 19272 31828
rect 19036 31272 19272 31508
rect 20036 31592 20272 31828
rect 20036 31272 20272 31508
rect 21036 31592 21272 31828
rect 21036 31272 21272 31508
rect 22036 31592 22272 31828
rect 22036 31272 22272 31508
rect 23036 31592 23272 31828
rect 23036 31272 23272 31508
rect 24036 31592 24272 31828
rect 24036 31272 24272 31508
rect 25036 31592 25272 31828
rect 25036 31272 25272 31508
rect 26036 31592 26272 31828
rect 26036 31272 26272 31508
rect 27036 31592 27272 31828
rect 27036 31272 27272 31508
rect 28036 31592 28272 31828
rect 28036 31272 28272 31508
rect 29036 31592 29272 31828
rect 29036 31272 29272 31508
rect 30036 31592 30272 31828
rect 30036 31272 30272 31508
rect 31036 31592 31272 31828
rect 31036 31272 31272 31508
rect 32036 31592 32272 31828
rect 32036 31272 32272 31508
rect 33036 31592 33272 31828
rect 33036 31272 33272 31508
rect 34036 31592 34272 31828
rect 34036 31272 34272 31508
rect -74783 30932 -74547 31168
rect -74443 30932 -74207 31168
rect -74103 30932 -73867 31168
rect -73783 30932 -73547 31168
rect -73443 30932 -73207 31168
rect -73103 30932 -72867 31168
rect -72783 30932 -72547 31168
rect -72443 30932 -72207 31168
rect -72103 30932 -71867 31168
rect -71783 30932 -71547 31168
rect -71443 30932 -71207 31168
rect -71103 30932 -70867 31168
rect -70783 30932 -70547 31168
rect -70443 30932 -70207 31168
rect -70103 30932 -69867 31168
rect -69783 30932 -69547 31168
rect -69443 30932 -69207 31168
rect -69103 30932 -68867 31168
rect -68783 30932 -68547 31168
rect -68443 30932 -68207 31168
rect -68103 30932 -67867 31168
rect -67783 30932 -67547 31168
rect -67443 30932 -67207 31168
rect -67103 30932 -66867 31168
rect -66783 30932 -66547 31168
rect -66443 30932 -66207 31168
rect -66103 30932 -65867 31168
rect -65783 30932 -65547 31168
rect -65443 30932 -65207 31168
rect -65103 30932 -64867 31168
rect -64783 30932 -64547 31168
rect -64443 30932 -64207 31168
rect -64103 30932 -63867 31168
rect -63783 30932 -63547 31168
rect -63443 30932 -63207 31168
rect -63103 30932 -62867 31168
rect -62783 30932 -62547 31168
rect -62443 30932 -62207 31168
rect -62103 30932 -61867 31168
rect -61783 30932 -61547 31168
rect -61443 30932 -61207 31168
rect -61103 30932 -60867 31168
rect -60783 30932 -60547 31168
rect -60443 30932 -60207 31168
rect -60103 30932 -59867 31168
rect -59783 30932 -59547 31168
rect -59443 30932 -59207 31168
rect -59103 30932 -58867 31168
rect 9696 30932 9932 31168
rect 10036 30932 10272 31168
rect 10376 30932 10612 31168
rect 10696 30932 10932 31168
rect 11036 30932 11272 31168
rect 11376 30932 11612 31168
rect 11696 30932 11932 31168
rect 12036 30932 12272 31168
rect 12376 30932 12612 31168
rect 12696 30932 12932 31168
rect 13036 30932 13272 31168
rect 13376 30932 13612 31168
rect 13696 30932 13932 31168
rect 14036 30932 14272 31168
rect 14376 30932 14612 31168
rect 14696 30932 14932 31168
rect 15036 30932 15272 31168
rect 15376 30932 15612 31168
rect 15696 30932 15932 31168
rect 16036 30932 16272 31168
rect 16376 30932 16612 31168
rect 16696 30932 16932 31168
rect 17036 30932 17272 31168
rect 17376 30932 17612 31168
rect 17696 30932 17932 31168
rect 18036 30932 18272 31168
rect 18376 30932 18612 31168
rect 18696 30932 18932 31168
rect 19036 30932 19272 31168
rect 19376 30932 19612 31168
rect 19696 30932 19932 31168
rect 20036 30932 20272 31168
rect 20376 30932 20612 31168
rect 20696 30932 20932 31168
rect 21036 30932 21272 31168
rect 21376 30932 21612 31168
rect 21696 30932 21932 31168
rect 22036 30932 22272 31168
rect 22376 30932 22612 31168
rect 22696 30932 22932 31168
rect 23036 30932 23272 31168
rect 23376 30932 23612 31168
rect 23696 30932 23932 31168
rect 24036 30932 24272 31168
rect 24376 30932 24612 31168
rect 24696 30932 24932 31168
rect 25036 30932 25272 31168
rect 25376 30932 25612 31168
rect 25696 30932 25932 31168
rect 26036 30932 26272 31168
rect 26376 30932 26612 31168
rect 26696 30932 26932 31168
rect 27036 30932 27272 31168
rect 27376 30932 27612 31168
rect 27696 30932 27932 31168
rect 28036 30932 28272 31168
rect 28376 30932 28612 31168
rect 28696 30932 28932 31168
rect 29036 30932 29272 31168
rect 29376 30932 29612 31168
rect 29696 30932 29932 31168
rect 30036 30932 30272 31168
rect 30376 30932 30612 31168
rect 30696 30932 30932 31168
rect 31036 30932 31272 31168
rect 31376 30932 31612 31168
rect 31696 30932 31932 31168
rect 32036 30932 32272 31168
rect 32376 30932 32612 31168
rect 32696 30932 32932 31168
rect 33036 30932 33272 31168
rect 33376 30932 33612 31168
rect 33696 30932 33932 31168
rect 34036 30932 34272 31168
rect 34376 30932 34612 31168
rect -74443 30592 -74207 30828
rect -74443 30272 -74207 30508
rect -73443 30592 -73207 30828
rect -73443 30272 -73207 30508
rect -72443 30592 -72207 30828
rect -72443 30272 -72207 30508
rect -71443 30592 -71207 30828
rect -71443 30272 -71207 30508
rect -70443 30592 -70207 30828
rect -70443 30272 -70207 30508
rect -69443 30592 -69207 30828
rect -69443 30272 -69207 30508
rect -68443 30592 -68207 30828
rect -68443 30272 -68207 30508
rect -67443 30592 -67207 30828
rect -67443 30272 -67207 30508
rect -66443 30592 -66207 30828
rect -66443 30272 -66207 30508
rect -65443 30592 -65207 30828
rect -65443 30272 -65207 30508
rect -64443 30592 -64207 30828
rect -64443 30272 -64207 30508
rect -63443 30592 -63207 30828
rect -63443 30272 -63207 30508
rect -62443 30592 -62207 30828
rect -62443 30272 -62207 30508
rect -61443 30592 -61207 30828
rect -61443 30272 -61207 30508
rect -60443 30592 -60207 30828
rect -60443 30272 -60207 30508
rect -59443 30592 -59207 30828
rect -59443 30272 -59207 30508
rect 10036 30592 10272 30828
rect 10036 30272 10272 30508
rect 11036 30592 11272 30828
rect 11036 30272 11272 30508
rect 12036 30592 12272 30828
rect 12036 30272 12272 30508
rect 13036 30592 13272 30828
rect 13036 30272 13272 30508
rect 14036 30592 14272 30828
rect 14036 30272 14272 30508
rect 15036 30592 15272 30828
rect 15036 30272 15272 30508
rect 16036 30592 16272 30828
rect 16036 30272 16272 30508
rect 17036 30592 17272 30828
rect 17036 30272 17272 30508
rect 18036 30592 18272 30828
rect 18036 30272 18272 30508
rect 19036 30592 19272 30828
rect 19036 30272 19272 30508
rect 20036 30592 20272 30828
rect 20036 30272 20272 30508
rect 21036 30592 21272 30828
rect 21036 30272 21272 30508
rect 22036 30592 22272 30828
rect 22036 30272 22272 30508
rect 23036 30592 23272 30828
rect 23036 30272 23272 30508
rect 24036 30592 24272 30828
rect 24036 30272 24272 30508
rect 25036 30592 25272 30828
rect 25036 30272 25272 30508
rect 26036 30592 26272 30828
rect 26036 30272 26272 30508
rect 27036 30592 27272 30828
rect 27036 30272 27272 30508
rect 28036 30592 28272 30828
rect 28036 30272 28272 30508
rect 29036 30592 29272 30828
rect 29036 30272 29272 30508
rect 30036 30592 30272 30828
rect 30036 30272 30272 30508
rect 31036 30592 31272 30828
rect 31036 30272 31272 30508
rect 32036 30592 32272 30828
rect 32036 30272 32272 30508
rect 33036 30592 33272 30828
rect 33036 30272 33272 30508
rect 34036 30592 34272 30828
rect 34036 30272 34272 30508
rect -74783 29932 -74547 30168
rect -74443 29932 -74207 30168
rect -74103 29932 -73867 30168
rect -73783 29932 -73547 30168
rect -73443 29932 -73207 30168
rect -73103 29932 -72867 30168
rect -72783 29932 -72547 30168
rect -72443 29932 -72207 30168
rect -72103 29932 -71867 30168
rect -71783 29932 -71547 30168
rect -71443 29932 -71207 30168
rect -71103 29932 -70867 30168
rect -70783 29932 -70547 30168
rect -70443 29932 -70207 30168
rect -70103 29932 -69867 30168
rect -69783 29932 -69547 30168
rect -69443 29932 -69207 30168
rect -69103 29932 -68867 30168
rect -68783 29932 -68547 30168
rect -68443 29932 -68207 30168
rect -68103 29932 -67867 30168
rect -67783 29932 -67547 30168
rect -67443 29932 -67207 30168
rect -67103 29932 -66867 30168
rect -66783 29932 -66547 30168
rect -66443 29932 -66207 30168
rect -66103 29932 -65867 30168
rect -65783 29932 -65547 30168
rect -65443 29932 -65207 30168
rect -65103 29932 -64867 30168
rect -64783 29932 -64547 30168
rect -64443 29932 -64207 30168
rect -64103 29932 -63867 30168
rect -63783 29932 -63547 30168
rect -63443 29932 -63207 30168
rect -63103 29932 -62867 30168
rect -62783 29932 -62547 30168
rect -62443 29932 -62207 30168
rect -62103 29932 -61867 30168
rect -61783 29932 -61547 30168
rect -61443 29932 -61207 30168
rect -61103 29932 -60867 30168
rect -60783 29932 -60547 30168
rect -60443 29932 -60207 30168
rect -60103 29932 -59867 30168
rect -59783 29932 -59547 30168
rect -59443 29932 -59207 30168
rect -59103 29932 -58867 30168
rect 9696 29932 9932 30168
rect 10036 29932 10272 30168
rect 10376 29932 10612 30168
rect 10696 29932 10932 30168
rect 11036 29932 11272 30168
rect 11376 29932 11612 30168
rect 11696 29932 11932 30168
rect 12036 29932 12272 30168
rect 12376 29932 12612 30168
rect 12696 29932 12932 30168
rect 13036 29932 13272 30168
rect 13376 29932 13612 30168
rect 13696 29932 13932 30168
rect 14036 29932 14272 30168
rect 14376 29932 14612 30168
rect 14696 29932 14932 30168
rect 15036 29932 15272 30168
rect 15376 29932 15612 30168
rect 15696 29932 15932 30168
rect 16036 29932 16272 30168
rect 16376 29932 16612 30168
rect 16696 29932 16932 30168
rect 17036 29932 17272 30168
rect 17376 29932 17612 30168
rect 17696 29932 17932 30168
rect 18036 29932 18272 30168
rect 18376 29932 18612 30168
rect 18696 29932 18932 30168
rect 19036 29932 19272 30168
rect 19376 29932 19612 30168
rect 19696 29932 19932 30168
rect 20036 29932 20272 30168
rect 20376 29932 20612 30168
rect 20696 29932 20932 30168
rect 21036 29932 21272 30168
rect 21376 29932 21612 30168
rect 21696 29932 21932 30168
rect 22036 29932 22272 30168
rect 22376 29932 22612 30168
rect 22696 29932 22932 30168
rect 23036 29932 23272 30168
rect 23376 29932 23612 30168
rect 23696 29932 23932 30168
rect 24036 29932 24272 30168
rect 24376 29932 24612 30168
rect 24696 29932 24932 30168
rect 25036 29932 25272 30168
rect 25376 29932 25612 30168
rect 25696 29932 25932 30168
rect 26036 29932 26272 30168
rect 26376 29932 26612 30168
rect 26696 29932 26932 30168
rect 27036 29932 27272 30168
rect 27376 29932 27612 30168
rect 27696 29932 27932 30168
rect 28036 29932 28272 30168
rect 28376 29932 28612 30168
rect 28696 29932 28932 30168
rect 29036 29932 29272 30168
rect 29376 29932 29612 30168
rect 29696 29932 29932 30168
rect 30036 29932 30272 30168
rect 30376 29932 30612 30168
rect 30696 29932 30932 30168
rect 31036 29932 31272 30168
rect 31376 29932 31612 30168
rect 31696 29932 31932 30168
rect 32036 29932 32272 30168
rect 32376 29932 32612 30168
rect 32696 29932 32932 30168
rect 33036 29932 33272 30168
rect 33376 29932 33612 30168
rect 33696 29932 33932 30168
rect 34036 29932 34272 30168
rect 34376 29932 34612 30168
rect -74443 29592 -74207 29828
rect -74443 29272 -74207 29508
rect -73443 29592 -73207 29828
rect -73443 29272 -73207 29508
rect -72443 29592 -72207 29828
rect -72443 29272 -72207 29508
rect -71443 29592 -71207 29828
rect -71443 29272 -71207 29508
rect -70443 29592 -70207 29828
rect -70443 29272 -70207 29508
rect -69443 29592 -69207 29828
rect -69443 29272 -69207 29508
rect -68443 29592 -68207 29828
rect -68443 29272 -68207 29508
rect -67443 29592 -67207 29828
rect -67443 29272 -67207 29508
rect -66443 29592 -66207 29828
rect -66443 29272 -66207 29508
rect -65443 29592 -65207 29828
rect -65443 29272 -65207 29508
rect -64443 29592 -64207 29828
rect -64443 29272 -64207 29508
rect -63443 29592 -63207 29828
rect -63443 29272 -63207 29508
rect -62443 29592 -62207 29828
rect -62443 29272 -62207 29508
rect -61443 29592 -61207 29828
rect -61443 29272 -61207 29508
rect -60443 29592 -60207 29828
rect -60443 29272 -60207 29508
rect -59443 29592 -59207 29828
rect -59443 29272 -59207 29508
rect 10036 29592 10272 29828
rect 10036 29272 10272 29508
rect 11036 29592 11272 29828
rect 11036 29272 11272 29508
rect 12036 29592 12272 29828
rect 12036 29272 12272 29508
rect 13036 29592 13272 29828
rect 13036 29272 13272 29508
rect 14036 29592 14272 29828
rect 14036 29272 14272 29508
rect 15036 29592 15272 29828
rect 15036 29272 15272 29508
rect 16036 29592 16272 29828
rect 16036 29272 16272 29508
rect 17036 29592 17272 29828
rect 17036 29272 17272 29508
rect 18036 29592 18272 29828
rect 18036 29272 18272 29508
rect 19036 29592 19272 29828
rect 19036 29272 19272 29508
rect 20036 29592 20272 29828
rect 20036 29272 20272 29508
rect 21036 29592 21272 29828
rect 21036 29272 21272 29508
rect 22036 29592 22272 29828
rect 22036 29272 22272 29508
rect 23036 29592 23272 29828
rect 23036 29272 23272 29508
rect 24036 29592 24272 29828
rect 24036 29272 24272 29508
rect 25036 29592 25272 29828
rect 25036 29272 25272 29508
rect 26036 29592 26272 29828
rect 26036 29272 26272 29508
rect 27036 29592 27272 29828
rect 27036 29272 27272 29508
rect 28036 29592 28272 29828
rect 28036 29272 28272 29508
rect 29036 29592 29272 29828
rect 29036 29272 29272 29508
rect 30036 29592 30272 29828
rect 30036 29272 30272 29508
rect 31036 29592 31272 29828
rect 31036 29272 31272 29508
rect 32036 29592 32272 29828
rect 32036 29272 32272 29508
rect 33036 29592 33272 29828
rect 33036 29272 33272 29508
rect 34036 29592 34272 29828
rect 34036 29272 34272 29508
rect -74783 28932 -74547 29168
rect -74443 28932 -74207 29168
rect -74103 28932 -73867 29168
rect -73783 28932 -73547 29168
rect -73443 28932 -73207 29168
rect -73103 28932 -72867 29168
rect -72783 28932 -72547 29168
rect -72443 28932 -72207 29168
rect -72103 28932 -71867 29168
rect -71783 28932 -71547 29168
rect -71443 28932 -71207 29168
rect -71103 28932 -70867 29168
rect -70783 28932 -70547 29168
rect -70443 28932 -70207 29168
rect -70103 28932 -69867 29168
rect -69783 28932 -69547 29168
rect -69443 28932 -69207 29168
rect -69103 28932 -68867 29168
rect -68783 28932 -68547 29168
rect -68443 28932 -68207 29168
rect -68103 28932 -67867 29168
rect -67783 28932 -67547 29168
rect -67443 28932 -67207 29168
rect -67103 28932 -66867 29168
rect -66783 28932 -66547 29168
rect -66443 28932 -66207 29168
rect -66103 28932 -65867 29168
rect -65783 28932 -65547 29168
rect -65443 28932 -65207 29168
rect -65103 28932 -64867 29168
rect -64783 28932 -64547 29168
rect -64443 28932 -64207 29168
rect -64103 28932 -63867 29168
rect -63783 28932 -63547 29168
rect -63443 28932 -63207 29168
rect -63103 28932 -62867 29168
rect -62783 28932 -62547 29168
rect -62443 28932 -62207 29168
rect -62103 28932 -61867 29168
rect -61783 28932 -61547 29168
rect -61443 28932 -61207 29168
rect -61103 28932 -60867 29168
rect -60783 28932 -60547 29168
rect -60443 28932 -60207 29168
rect -60103 28932 -59867 29168
rect -59783 28932 -59547 29168
rect -59443 28932 -59207 29168
rect -59103 28932 -58867 29168
rect 9696 28932 9932 29168
rect 10036 28932 10272 29168
rect 10376 28932 10612 29168
rect 10696 28932 10932 29168
rect 11036 28932 11272 29168
rect 11376 28932 11612 29168
rect 11696 28932 11932 29168
rect 12036 28932 12272 29168
rect 12376 28932 12612 29168
rect 12696 28932 12932 29168
rect 13036 28932 13272 29168
rect 13376 28932 13612 29168
rect 13696 28932 13932 29168
rect 14036 28932 14272 29168
rect 14376 28932 14612 29168
rect 14696 28932 14932 29168
rect 15036 28932 15272 29168
rect 15376 28932 15612 29168
rect 15696 28932 15932 29168
rect 16036 28932 16272 29168
rect 16376 28932 16612 29168
rect 16696 28932 16932 29168
rect 17036 28932 17272 29168
rect 17376 28932 17612 29168
rect 17696 28932 17932 29168
rect 18036 28932 18272 29168
rect 18376 28932 18612 29168
rect 18696 28932 18932 29168
rect 19036 28932 19272 29168
rect 19376 28932 19612 29168
rect 19696 28932 19932 29168
rect 20036 28932 20272 29168
rect 20376 28932 20612 29168
rect 20696 28932 20932 29168
rect 21036 28932 21272 29168
rect 21376 28932 21612 29168
rect 21696 28932 21932 29168
rect 22036 28932 22272 29168
rect 22376 28932 22612 29168
rect 22696 28932 22932 29168
rect 23036 28932 23272 29168
rect 23376 28932 23612 29168
rect 23696 28932 23932 29168
rect 24036 28932 24272 29168
rect 24376 28932 24612 29168
rect 24696 28932 24932 29168
rect 25036 28932 25272 29168
rect 25376 28932 25612 29168
rect 25696 28932 25932 29168
rect 26036 28932 26272 29168
rect 26376 28932 26612 29168
rect 26696 28932 26932 29168
rect 27036 28932 27272 29168
rect 27376 28932 27612 29168
rect 27696 28932 27932 29168
rect 28036 28932 28272 29168
rect 28376 28932 28612 29168
rect 28696 28932 28932 29168
rect 29036 28932 29272 29168
rect 29376 28932 29612 29168
rect 29696 28932 29932 29168
rect 30036 28932 30272 29168
rect 30376 28932 30612 29168
rect 30696 28932 30932 29168
rect 31036 28932 31272 29168
rect 31376 28932 31612 29168
rect 31696 28932 31932 29168
rect 32036 28932 32272 29168
rect 32376 28932 32612 29168
rect 32696 28932 32932 29168
rect 33036 28932 33272 29168
rect 33376 28932 33612 29168
rect 33696 28932 33932 29168
rect 34036 28932 34272 29168
rect 34376 28932 34612 29168
rect -74443 28592 -74207 28828
rect -73443 28592 -73207 28828
rect -72443 28592 -72207 28828
rect -71443 28592 -71207 28828
rect -70443 28592 -70207 28828
rect -69443 28592 -69207 28828
rect -68443 28592 -68207 28828
rect -67443 28592 -67207 28828
rect -66443 28592 -66207 28828
rect -65443 28592 -65207 28828
rect -64443 28592 -64207 28828
rect -63443 28592 -63207 28828
rect -62443 28592 -62207 28828
rect -61443 28592 -61207 28828
rect -60443 28592 -60207 28828
rect -59443 28592 -59207 28828
rect 10036 28592 10272 28828
rect 11036 28592 11272 28828
rect 12036 28592 12272 28828
rect 13036 28592 13272 28828
rect 14036 28592 14272 28828
rect 15036 28592 15272 28828
rect 16036 28592 16272 28828
rect 17036 28592 17272 28828
rect 18036 28592 18272 28828
rect 19036 28592 19272 28828
rect 20036 28592 20272 28828
rect 21036 28592 21272 28828
rect 22036 28592 22272 28828
rect 23036 28592 23272 28828
rect 24036 28592 24272 28828
rect 25036 28592 25272 28828
rect 26036 28592 26272 28828
rect 27036 28592 27272 28828
rect 28036 28592 28272 28828
rect 29036 28592 29272 28828
rect 30036 28592 30272 28828
rect 31036 28592 31272 28828
rect 32036 28592 32272 28828
rect 33036 28592 33272 28828
rect 34036 28592 34272 28828
rect -72708 16082 -60952 25918
rect 20392 16082 32148 25918
rect -42308 8012 -40792 13688
rect -24233 8012 -16317 13688
rect -42308 -2198 -40792 2198
rect 242 8012 1758 13688
rect 242 -2198 1758 2198
rect -42308 -13688 -40792 -8012
rect -29423 -13693 -28227 -8017
rect -12323 -13702 -11127 -8026
rect 242 -13688 1758 -8012
rect -72708 -25918 -60952 -16082
rect 20392 -25918 32148 -16082
rect -74443 -28828 -74207 -28592
rect -73443 -28828 -73207 -28592
rect -72443 -28828 -72207 -28592
rect -71443 -28828 -71207 -28592
rect -70443 -28828 -70207 -28592
rect -69443 -28828 -69207 -28592
rect -68443 -28828 -68207 -28592
rect -67443 -28828 -67207 -28592
rect -66443 -28828 -66207 -28592
rect -65443 -28828 -65207 -28592
rect -64443 -28828 -64207 -28592
rect -63443 -28828 -63207 -28592
rect -62443 -28828 -62207 -28592
rect -61443 -28828 -61207 -28592
rect -60443 -28828 -60207 -28592
rect -59443 -28828 -59207 -28592
rect -58443 -28828 -58207 -28592
rect -57443 -28828 -57207 -28592
rect -56443 -28828 -56207 -28592
rect -55443 -28828 -55207 -28592
rect -54443 -28828 -54207 -28592
rect -53443 -28828 -53207 -28592
rect -52443 -28828 -52207 -28592
rect -51443 -28828 -51207 -28592
rect -50443 -28828 -50207 -28592
rect -49443 -28828 -49207 -28592
rect 8657 -28828 8893 -28592
rect 9657 -28828 9893 -28592
rect 10657 -28828 10893 -28592
rect 11657 -28828 11893 -28592
rect 12657 -28828 12893 -28592
rect 13657 -28828 13893 -28592
rect 14657 -28828 14893 -28592
rect 15657 -28828 15893 -28592
rect 16657 -28828 16893 -28592
rect 17657 -28828 17893 -28592
rect 18657 -28828 18893 -28592
rect 19657 -28828 19893 -28592
rect 20657 -28828 20893 -28592
rect 21657 -28828 21893 -28592
rect 22657 -28828 22893 -28592
rect 23657 -28828 23893 -28592
rect 24657 -28828 24893 -28592
rect 25657 -28828 25893 -28592
rect 26657 -28828 26893 -28592
rect 27657 -28828 27893 -28592
rect 28657 -28828 28893 -28592
rect 29657 -28828 29893 -28592
rect 30657 -28828 30893 -28592
rect 31657 -28828 31893 -28592
rect 32657 -28828 32893 -28592
rect 33657 -28828 33893 -28592
rect -74783 -29168 -74547 -28932
rect -74443 -29168 -74207 -28932
rect -74103 -29168 -73867 -28932
rect -73783 -29168 -73547 -28932
rect -73443 -29168 -73207 -28932
rect -73103 -29168 -72867 -28932
rect -72783 -29168 -72547 -28932
rect -72443 -29168 -72207 -28932
rect -72103 -29168 -71867 -28932
rect -71783 -29168 -71547 -28932
rect -71443 -29168 -71207 -28932
rect -71103 -29168 -70867 -28932
rect -70783 -29168 -70547 -28932
rect -70443 -29168 -70207 -28932
rect -70103 -29168 -69867 -28932
rect -69783 -29168 -69547 -28932
rect -69443 -29168 -69207 -28932
rect -69103 -29168 -68867 -28932
rect -68783 -29168 -68547 -28932
rect -68443 -29168 -68207 -28932
rect -68103 -29168 -67867 -28932
rect -67783 -29168 -67547 -28932
rect -67443 -29168 -67207 -28932
rect -67103 -29168 -66867 -28932
rect -66783 -29168 -66547 -28932
rect -66443 -29168 -66207 -28932
rect -66103 -29168 -65867 -28932
rect -65783 -29168 -65547 -28932
rect -65443 -29168 -65207 -28932
rect -65103 -29168 -64867 -28932
rect -64783 -29168 -64547 -28932
rect -64443 -29168 -64207 -28932
rect -64103 -29168 -63867 -28932
rect -63783 -29168 -63547 -28932
rect -63443 -29168 -63207 -28932
rect -63103 -29168 -62867 -28932
rect -62783 -29168 -62547 -28932
rect -62443 -29168 -62207 -28932
rect -62103 -29168 -61867 -28932
rect -61783 -29168 -61547 -28932
rect -61443 -29168 -61207 -28932
rect -61103 -29168 -60867 -28932
rect -60783 -29168 -60547 -28932
rect -60443 -29168 -60207 -28932
rect -60103 -29168 -59867 -28932
rect -59783 -29168 -59547 -28932
rect -59443 -29168 -59207 -28932
rect -59103 -29168 -58867 -28932
rect -58783 -29168 -58547 -28932
rect -58443 -29168 -58207 -28932
rect -58103 -29168 -57867 -28932
rect -57783 -29168 -57547 -28932
rect -57443 -29168 -57207 -28932
rect -57103 -29168 -56867 -28932
rect -56783 -29168 -56547 -28932
rect -56443 -29168 -56207 -28932
rect -56103 -29168 -55867 -28932
rect -55783 -29168 -55547 -28932
rect -55443 -29168 -55207 -28932
rect -55103 -29168 -54867 -28932
rect -54783 -29168 -54547 -28932
rect -54443 -29168 -54207 -28932
rect -54103 -29168 -53867 -28932
rect -53783 -29168 -53547 -28932
rect -53443 -29168 -53207 -28932
rect -53103 -29168 -52867 -28932
rect -52783 -29168 -52547 -28932
rect -52443 -29168 -52207 -28932
rect -52103 -29168 -51867 -28932
rect -51783 -29168 -51547 -28932
rect -51443 -29168 -51207 -28932
rect -51103 -29168 -50867 -28932
rect -50783 -29168 -50547 -28932
rect -50443 -29168 -50207 -28932
rect -50103 -29168 -49867 -28932
rect -49783 -29168 -49547 -28932
rect -49443 -29168 -49207 -28932
rect -49103 -29168 -48867 -28932
rect 8317 -29168 8553 -28932
rect 8657 -29168 8893 -28932
rect 8997 -29168 9233 -28932
rect 9317 -29168 9553 -28932
rect 9657 -29168 9893 -28932
rect 9997 -29168 10233 -28932
rect 10317 -29168 10553 -28932
rect 10657 -29168 10893 -28932
rect 10997 -29168 11233 -28932
rect 11317 -29168 11553 -28932
rect 11657 -29168 11893 -28932
rect 11997 -29168 12233 -28932
rect 12317 -29168 12553 -28932
rect 12657 -29168 12893 -28932
rect 12997 -29168 13233 -28932
rect 13317 -29168 13553 -28932
rect 13657 -29168 13893 -28932
rect 13997 -29168 14233 -28932
rect 14317 -29168 14553 -28932
rect 14657 -29168 14893 -28932
rect 14997 -29168 15233 -28932
rect 15317 -29168 15553 -28932
rect 15657 -29168 15893 -28932
rect 15997 -29168 16233 -28932
rect 16317 -29168 16553 -28932
rect 16657 -29168 16893 -28932
rect 16997 -29168 17233 -28932
rect 17317 -29168 17553 -28932
rect 17657 -29168 17893 -28932
rect 17997 -29168 18233 -28932
rect 18317 -29168 18553 -28932
rect 18657 -29168 18893 -28932
rect 18997 -29168 19233 -28932
rect 19317 -29168 19553 -28932
rect 19657 -29168 19893 -28932
rect 19997 -29168 20233 -28932
rect 20317 -29168 20553 -28932
rect 20657 -29168 20893 -28932
rect 20997 -29168 21233 -28932
rect 21317 -29168 21553 -28932
rect 21657 -29168 21893 -28932
rect 21997 -29168 22233 -28932
rect 22317 -29168 22553 -28932
rect 22657 -29168 22893 -28932
rect 22997 -29168 23233 -28932
rect 23317 -29168 23553 -28932
rect 23657 -29168 23893 -28932
rect 23997 -29168 24233 -28932
rect 24317 -29168 24553 -28932
rect 24657 -29168 24893 -28932
rect 24997 -29168 25233 -28932
rect 25317 -29168 25553 -28932
rect 25657 -29168 25893 -28932
rect 25997 -29168 26233 -28932
rect 26317 -29168 26553 -28932
rect 26657 -29168 26893 -28932
rect 26997 -29168 27233 -28932
rect 27317 -29168 27553 -28932
rect 27657 -29168 27893 -28932
rect 27997 -29168 28233 -28932
rect 28317 -29168 28553 -28932
rect 28657 -29168 28893 -28932
rect 28997 -29168 29233 -28932
rect 29317 -29168 29553 -28932
rect 29657 -29168 29893 -28932
rect 29997 -29168 30233 -28932
rect 30317 -29168 30553 -28932
rect 30657 -29168 30893 -28932
rect 30997 -29168 31233 -28932
rect 31317 -29168 31553 -28932
rect 31657 -29168 31893 -28932
rect 31997 -29168 32233 -28932
rect 32317 -29168 32553 -28932
rect 32657 -29168 32893 -28932
rect 32997 -29168 33233 -28932
rect 33317 -29168 33553 -28932
rect 33657 -29168 33893 -28932
rect 33997 -29168 34233 -28932
rect -74443 -29508 -74207 -29272
rect -74443 -29828 -74207 -29592
rect -73443 -29508 -73207 -29272
rect -73443 -29828 -73207 -29592
rect -72443 -29508 -72207 -29272
rect -72443 -29828 -72207 -29592
rect -71443 -29508 -71207 -29272
rect -71443 -29828 -71207 -29592
rect -70443 -29508 -70207 -29272
rect -70443 -29828 -70207 -29592
rect -69443 -29508 -69207 -29272
rect -69443 -29828 -69207 -29592
rect -68443 -29508 -68207 -29272
rect -68443 -29828 -68207 -29592
rect -67443 -29508 -67207 -29272
rect -67443 -29828 -67207 -29592
rect -66443 -29508 -66207 -29272
rect -66443 -29828 -66207 -29592
rect -65443 -29508 -65207 -29272
rect -65443 -29828 -65207 -29592
rect -64443 -29508 -64207 -29272
rect -64443 -29828 -64207 -29592
rect -63443 -29508 -63207 -29272
rect -63443 -29828 -63207 -29592
rect -62443 -29508 -62207 -29272
rect -62443 -29828 -62207 -29592
rect -61443 -29508 -61207 -29272
rect -61443 -29828 -61207 -29592
rect -60443 -29508 -60207 -29272
rect -60443 -29828 -60207 -29592
rect -59443 -29508 -59207 -29272
rect -59443 -29828 -59207 -29592
rect -58443 -29508 -58207 -29272
rect -58443 -29828 -58207 -29592
rect -57443 -29508 -57207 -29272
rect -57443 -29828 -57207 -29592
rect -56443 -29508 -56207 -29272
rect -56443 -29828 -56207 -29592
rect -55443 -29508 -55207 -29272
rect -55443 -29828 -55207 -29592
rect -54443 -29508 -54207 -29272
rect -54443 -29828 -54207 -29592
rect -53443 -29508 -53207 -29272
rect -53443 -29828 -53207 -29592
rect -52443 -29508 -52207 -29272
rect -52443 -29828 -52207 -29592
rect -51443 -29508 -51207 -29272
rect -51443 -29828 -51207 -29592
rect -50443 -29508 -50207 -29272
rect -50443 -29828 -50207 -29592
rect -49443 -29508 -49207 -29272
rect -49443 -29828 -49207 -29592
rect 8657 -29508 8893 -29272
rect 8657 -29828 8893 -29592
rect 9657 -29508 9893 -29272
rect 9657 -29828 9893 -29592
rect 10657 -29508 10893 -29272
rect 10657 -29828 10893 -29592
rect 11657 -29508 11893 -29272
rect 11657 -29828 11893 -29592
rect 12657 -29508 12893 -29272
rect 12657 -29828 12893 -29592
rect 13657 -29508 13893 -29272
rect 13657 -29828 13893 -29592
rect 14657 -29508 14893 -29272
rect 14657 -29828 14893 -29592
rect 15657 -29508 15893 -29272
rect 15657 -29828 15893 -29592
rect 16657 -29508 16893 -29272
rect 16657 -29828 16893 -29592
rect 17657 -29508 17893 -29272
rect 17657 -29828 17893 -29592
rect 18657 -29508 18893 -29272
rect 18657 -29828 18893 -29592
rect 19657 -29508 19893 -29272
rect 19657 -29828 19893 -29592
rect 20657 -29508 20893 -29272
rect 20657 -29828 20893 -29592
rect 21657 -29508 21893 -29272
rect 21657 -29828 21893 -29592
rect 22657 -29508 22893 -29272
rect 22657 -29828 22893 -29592
rect 23657 -29508 23893 -29272
rect 23657 -29828 23893 -29592
rect 24657 -29508 24893 -29272
rect 24657 -29828 24893 -29592
rect 25657 -29508 25893 -29272
rect 25657 -29828 25893 -29592
rect 26657 -29508 26893 -29272
rect 26657 -29828 26893 -29592
rect 27657 -29508 27893 -29272
rect 27657 -29828 27893 -29592
rect 28657 -29508 28893 -29272
rect 28657 -29828 28893 -29592
rect 29657 -29508 29893 -29272
rect 29657 -29828 29893 -29592
rect 30657 -29508 30893 -29272
rect 30657 -29828 30893 -29592
rect 31657 -29508 31893 -29272
rect 31657 -29828 31893 -29592
rect 32657 -29508 32893 -29272
rect 32657 -29828 32893 -29592
rect 33657 -29508 33893 -29272
rect 33657 -29828 33893 -29592
rect -74783 -30168 -74547 -29932
rect -74443 -30168 -74207 -29932
rect -74103 -30168 -73867 -29932
rect -73783 -30168 -73547 -29932
rect -73443 -30168 -73207 -29932
rect -73103 -30168 -72867 -29932
rect -72783 -30168 -72547 -29932
rect -72443 -30168 -72207 -29932
rect -72103 -30168 -71867 -29932
rect -71783 -30168 -71547 -29932
rect -71443 -30168 -71207 -29932
rect -71103 -30168 -70867 -29932
rect -70783 -30168 -70547 -29932
rect -70443 -30168 -70207 -29932
rect -70103 -30168 -69867 -29932
rect -69783 -30168 -69547 -29932
rect -69443 -30168 -69207 -29932
rect -69103 -30168 -68867 -29932
rect -68783 -30168 -68547 -29932
rect -68443 -30168 -68207 -29932
rect -68103 -30168 -67867 -29932
rect -67783 -30168 -67547 -29932
rect -67443 -30168 -67207 -29932
rect -67103 -30168 -66867 -29932
rect -66783 -30168 -66547 -29932
rect -66443 -30168 -66207 -29932
rect -66103 -30168 -65867 -29932
rect -65783 -30168 -65547 -29932
rect -65443 -30168 -65207 -29932
rect -65103 -30168 -64867 -29932
rect -64783 -30168 -64547 -29932
rect -64443 -30168 -64207 -29932
rect -64103 -30168 -63867 -29932
rect -63783 -30168 -63547 -29932
rect -63443 -30168 -63207 -29932
rect -63103 -30168 -62867 -29932
rect -62783 -30168 -62547 -29932
rect -62443 -30168 -62207 -29932
rect -62103 -30168 -61867 -29932
rect -61783 -30168 -61547 -29932
rect -61443 -30168 -61207 -29932
rect -61103 -30168 -60867 -29932
rect -60783 -30168 -60547 -29932
rect -60443 -30168 -60207 -29932
rect -60103 -30168 -59867 -29932
rect -59783 -30168 -59547 -29932
rect -59443 -30168 -59207 -29932
rect -59103 -30168 -58867 -29932
rect -58783 -30168 -58547 -29932
rect -58443 -30168 -58207 -29932
rect -58103 -30168 -57867 -29932
rect -57783 -30168 -57547 -29932
rect -57443 -30168 -57207 -29932
rect -57103 -30168 -56867 -29932
rect -56783 -30168 -56547 -29932
rect -56443 -30168 -56207 -29932
rect -56103 -30168 -55867 -29932
rect -55783 -30168 -55547 -29932
rect -55443 -30168 -55207 -29932
rect -55103 -30168 -54867 -29932
rect -54783 -30168 -54547 -29932
rect -54443 -30168 -54207 -29932
rect -54103 -30168 -53867 -29932
rect -53783 -30168 -53547 -29932
rect -53443 -30168 -53207 -29932
rect -53103 -30168 -52867 -29932
rect -52783 -30168 -52547 -29932
rect -52443 -30168 -52207 -29932
rect -52103 -30168 -51867 -29932
rect -51783 -30168 -51547 -29932
rect -51443 -30168 -51207 -29932
rect -51103 -30168 -50867 -29932
rect -50783 -30168 -50547 -29932
rect -50443 -30168 -50207 -29932
rect -50103 -30168 -49867 -29932
rect -49783 -30168 -49547 -29932
rect -49443 -30168 -49207 -29932
rect -49103 -30168 -48867 -29932
rect 8317 -30168 8553 -29932
rect 8657 -30168 8893 -29932
rect 8997 -30168 9233 -29932
rect 9317 -30168 9553 -29932
rect 9657 -30168 9893 -29932
rect 9997 -30168 10233 -29932
rect 10317 -30168 10553 -29932
rect 10657 -30168 10893 -29932
rect 10997 -30168 11233 -29932
rect 11317 -30168 11553 -29932
rect 11657 -30168 11893 -29932
rect 11997 -30168 12233 -29932
rect 12317 -30168 12553 -29932
rect 12657 -30168 12893 -29932
rect 12997 -30168 13233 -29932
rect 13317 -30168 13553 -29932
rect 13657 -30168 13893 -29932
rect 13997 -30168 14233 -29932
rect 14317 -30168 14553 -29932
rect 14657 -30168 14893 -29932
rect 14997 -30168 15233 -29932
rect 15317 -30168 15553 -29932
rect 15657 -30168 15893 -29932
rect 15997 -30168 16233 -29932
rect 16317 -30168 16553 -29932
rect 16657 -30168 16893 -29932
rect 16997 -30168 17233 -29932
rect 17317 -30168 17553 -29932
rect 17657 -30168 17893 -29932
rect 17997 -30168 18233 -29932
rect 18317 -30168 18553 -29932
rect 18657 -30168 18893 -29932
rect 18997 -30168 19233 -29932
rect 19317 -30168 19553 -29932
rect 19657 -30168 19893 -29932
rect 19997 -30168 20233 -29932
rect 20317 -30168 20553 -29932
rect 20657 -30168 20893 -29932
rect 20997 -30168 21233 -29932
rect 21317 -30168 21553 -29932
rect 21657 -30168 21893 -29932
rect 21997 -30168 22233 -29932
rect 22317 -30168 22553 -29932
rect 22657 -30168 22893 -29932
rect 22997 -30168 23233 -29932
rect 23317 -30168 23553 -29932
rect 23657 -30168 23893 -29932
rect 23997 -30168 24233 -29932
rect 24317 -30168 24553 -29932
rect 24657 -30168 24893 -29932
rect 24997 -30168 25233 -29932
rect 25317 -30168 25553 -29932
rect 25657 -30168 25893 -29932
rect 25997 -30168 26233 -29932
rect 26317 -30168 26553 -29932
rect 26657 -30168 26893 -29932
rect 26997 -30168 27233 -29932
rect 27317 -30168 27553 -29932
rect 27657 -30168 27893 -29932
rect 27997 -30168 28233 -29932
rect 28317 -30168 28553 -29932
rect 28657 -30168 28893 -29932
rect 28997 -30168 29233 -29932
rect 29317 -30168 29553 -29932
rect 29657 -30168 29893 -29932
rect 29997 -30168 30233 -29932
rect 30317 -30168 30553 -29932
rect 30657 -30168 30893 -29932
rect 30997 -30168 31233 -29932
rect 31317 -30168 31553 -29932
rect 31657 -30168 31893 -29932
rect 31997 -30168 32233 -29932
rect 32317 -30168 32553 -29932
rect 32657 -30168 32893 -29932
rect 32997 -30168 33233 -29932
rect 33317 -30168 33553 -29932
rect 33657 -30168 33893 -29932
rect 33997 -30168 34233 -29932
rect -74443 -30508 -74207 -30272
rect -74443 -30828 -74207 -30592
rect -73443 -30508 -73207 -30272
rect -73443 -30828 -73207 -30592
rect -72443 -30508 -72207 -30272
rect -72443 -30828 -72207 -30592
rect -71443 -30508 -71207 -30272
rect -71443 -30828 -71207 -30592
rect -70443 -30508 -70207 -30272
rect -70443 -30828 -70207 -30592
rect -69443 -30508 -69207 -30272
rect -69443 -30828 -69207 -30592
rect -68443 -30508 -68207 -30272
rect -68443 -30828 -68207 -30592
rect -67443 -30508 -67207 -30272
rect -67443 -30828 -67207 -30592
rect -66443 -30508 -66207 -30272
rect -66443 -30828 -66207 -30592
rect -65443 -30508 -65207 -30272
rect -65443 -30828 -65207 -30592
rect -64443 -30508 -64207 -30272
rect -64443 -30828 -64207 -30592
rect -63443 -30508 -63207 -30272
rect -63443 -30828 -63207 -30592
rect -62443 -30508 -62207 -30272
rect -62443 -30828 -62207 -30592
rect -61443 -30508 -61207 -30272
rect -61443 -30828 -61207 -30592
rect -60443 -30508 -60207 -30272
rect -60443 -30828 -60207 -30592
rect -59443 -30508 -59207 -30272
rect -59443 -30828 -59207 -30592
rect -58443 -30508 -58207 -30272
rect -58443 -30828 -58207 -30592
rect -57443 -30508 -57207 -30272
rect -57443 -30828 -57207 -30592
rect -56443 -30508 -56207 -30272
rect -56443 -30828 -56207 -30592
rect -55443 -30508 -55207 -30272
rect -55443 -30828 -55207 -30592
rect -54443 -30508 -54207 -30272
rect -54443 -30828 -54207 -30592
rect -53443 -30508 -53207 -30272
rect -53443 -30828 -53207 -30592
rect -52443 -30508 -52207 -30272
rect -52443 -30828 -52207 -30592
rect -51443 -30508 -51207 -30272
rect -51443 -30828 -51207 -30592
rect -50443 -30508 -50207 -30272
rect -50443 -30828 -50207 -30592
rect -49443 -30508 -49207 -30272
rect -49443 -30828 -49207 -30592
rect 8657 -30508 8893 -30272
rect 8657 -30828 8893 -30592
rect 9657 -30508 9893 -30272
rect 9657 -30828 9893 -30592
rect 10657 -30508 10893 -30272
rect 10657 -30828 10893 -30592
rect 11657 -30508 11893 -30272
rect 11657 -30828 11893 -30592
rect 12657 -30508 12893 -30272
rect 12657 -30828 12893 -30592
rect 13657 -30508 13893 -30272
rect 13657 -30828 13893 -30592
rect 14657 -30508 14893 -30272
rect 14657 -30828 14893 -30592
rect 15657 -30508 15893 -30272
rect 15657 -30828 15893 -30592
rect 16657 -30508 16893 -30272
rect 16657 -30828 16893 -30592
rect 17657 -30508 17893 -30272
rect 17657 -30828 17893 -30592
rect 18657 -30508 18893 -30272
rect 18657 -30828 18893 -30592
rect 19657 -30508 19893 -30272
rect 19657 -30828 19893 -30592
rect 20657 -30508 20893 -30272
rect 20657 -30828 20893 -30592
rect 21657 -30508 21893 -30272
rect 21657 -30828 21893 -30592
rect 22657 -30508 22893 -30272
rect 22657 -30828 22893 -30592
rect 23657 -30508 23893 -30272
rect 23657 -30828 23893 -30592
rect 24657 -30508 24893 -30272
rect 24657 -30828 24893 -30592
rect 25657 -30508 25893 -30272
rect 25657 -30828 25893 -30592
rect 26657 -30508 26893 -30272
rect 26657 -30828 26893 -30592
rect 27657 -30508 27893 -30272
rect 27657 -30828 27893 -30592
rect 28657 -30508 28893 -30272
rect 28657 -30828 28893 -30592
rect 29657 -30508 29893 -30272
rect 29657 -30828 29893 -30592
rect 30657 -30508 30893 -30272
rect 30657 -30828 30893 -30592
rect 31657 -30508 31893 -30272
rect 31657 -30828 31893 -30592
rect 32657 -30508 32893 -30272
rect 32657 -30828 32893 -30592
rect 33657 -30508 33893 -30272
rect 33657 -30828 33893 -30592
rect -74783 -31168 -74547 -30932
rect -74443 -31168 -74207 -30932
rect -74103 -31168 -73867 -30932
rect -73783 -31168 -73547 -30932
rect -73443 -31168 -73207 -30932
rect -73103 -31168 -72867 -30932
rect -72783 -31168 -72547 -30932
rect -72443 -31168 -72207 -30932
rect -72103 -31168 -71867 -30932
rect -71783 -31168 -71547 -30932
rect -71443 -31168 -71207 -30932
rect -71103 -31168 -70867 -30932
rect -70783 -31168 -70547 -30932
rect -70443 -31168 -70207 -30932
rect -70103 -31168 -69867 -30932
rect -69783 -31168 -69547 -30932
rect -69443 -31168 -69207 -30932
rect -69103 -31168 -68867 -30932
rect -68783 -31168 -68547 -30932
rect -68443 -31168 -68207 -30932
rect -68103 -31168 -67867 -30932
rect -67783 -31168 -67547 -30932
rect -67443 -31168 -67207 -30932
rect -67103 -31168 -66867 -30932
rect -66783 -31168 -66547 -30932
rect -66443 -31168 -66207 -30932
rect -66103 -31168 -65867 -30932
rect -65783 -31168 -65547 -30932
rect -65443 -31168 -65207 -30932
rect -65103 -31168 -64867 -30932
rect -64783 -31168 -64547 -30932
rect -64443 -31168 -64207 -30932
rect -64103 -31168 -63867 -30932
rect -63783 -31168 -63547 -30932
rect -63443 -31168 -63207 -30932
rect -63103 -31168 -62867 -30932
rect -62783 -31168 -62547 -30932
rect -62443 -31168 -62207 -30932
rect -62103 -31168 -61867 -30932
rect -61783 -31168 -61547 -30932
rect -61443 -31168 -61207 -30932
rect -61103 -31168 -60867 -30932
rect -60783 -31168 -60547 -30932
rect -60443 -31168 -60207 -30932
rect -60103 -31168 -59867 -30932
rect -59783 -31168 -59547 -30932
rect -59443 -31168 -59207 -30932
rect -59103 -31168 -58867 -30932
rect -58783 -31168 -58547 -30932
rect -58443 -31168 -58207 -30932
rect -58103 -31168 -57867 -30932
rect -57783 -31168 -57547 -30932
rect -57443 -31168 -57207 -30932
rect -57103 -31168 -56867 -30932
rect -56783 -31168 -56547 -30932
rect -56443 -31168 -56207 -30932
rect -56103 -31168 -55867 -30932
rect -55783 -31168 -55547 -30932
rect -55443 -31168 -55207 -30932
rect -55103 -31168 -54867 -30932
rect -54783 -31168 -54547 -30932
rect -54443 -31168 -54207 -30932
rect -54103 -31168 -53867 -30932
rect -53783 -31168 -53547 -30932
rect -53443 -31168 -53207 -30932
rect -53103 -31168 -52867 -30932
rect -52783 -31168 -52547 -30932
rect -52443 -31168 -52207 -30932
rect -52103 -31168 -51867 -30932
rect -51783 -31168 -51547 -30932
rect -51443 -31168 -51207 -30932
rect -51103 -31168 -50867 -30932
rect -50783 -31168 -50547 -30932
rect -50443 -31168 -50207 -30932
rect -50103 -31168 -49867 -30932
rect -49783 -31168 -49547 -30932
rect -49443 -31168 -49207 -30932
rect -49103 -31168 -48867 -30932
rect 8317 -31168 8553 -30932
rect 8657 -31168 8893 -30932
rect 8997 -31168 9233 -30932
rect 9317 -31168 9553 -30932
rect 9657 -31168 9893 -30932
rect 9997 -31168 10233 -30932
rect 10317 -31168 10553 -30932
rect 10657 -31168 10893 -30932
rect 10997 -31168 11233 -30932
rect 11317 -31168 11553 -30932
rect 11657 -31168 11893 -30932
rect 11997 -31168 12233 -30932
rect 12317 -31168 12553 -30932
rect 12657 -31168 12893 -30932
rect 12997 -31168 13233 -30932
rect 13317 -31168 13553 -30932
rect 13657 -31168 13893 -30932
rect 13997 -31168 14233 -30932
rect 14317 -31168 14553 -30932
rect 14657 -31168 14893 -30932
rect 14997 -31168 15233 -30932
rect 15317 -31168 15553 -30932
rect 15657 -31168 15893 -30932
rect 15997 -31168 16233 -30932
rect 16317 -31168 16553 -30932
rect 16657 -31168 16893 -30932
rect 16997 -31168 17233 -30932
rect 17317 -31168 17553 -30932
rect 17657 -31168 17893 -30932
rect 17997 -31168 18233 -30932
rect 18317 -31168 18553 -30932
rect 18657 -31168 18893 -30932
rect 18997 -31168 19233 -30932
rect 19317 -31168 19553 -30932
rect 19657 -31168 19893 -30932
rect 19997 -31168 20233 -30932
rect 20317 -31168 20553 -30932
rect 20657 -31168 20893 -30932
rect 20997 -31168 21233 -30932
rect 21317 -31168 21553 -30932
rect 21657 -31168 21893 -30932
rect 21997 -31168 22233 -30932
rect 22317 -31168 22553 -30932
rect 22657 -31168 22893 -30932
rect 22997 -31168 23233 -30932
rect 23317 -31168 23553 -30932
rect 23657 -31168 23893 -30932
rect 23997 -31168 24233 -30932
rect 24317 -31168 24553 -30932
rect 24657 -31168 24893 -30932
rect 24997 -31168 25233 -30932
rect 25317 -31168 25553 -30932
rect 25657 -31168 25893 -30932
rect 25997 -31168 26233 -30932
rect 26317 -31168 26553 -30932
rect 26657 -31168 26893 -30932
rect 26997 -31168 27233 -30932
rect 27317 -31168 27553 -30932
rect 27657 -31168 27893 -30932
rect 27997 -31168 28233 -30932
rect 28317 -31168 28553 -30932
rect 28657 -31168 28893 -30932
rect 28997 -31168 29233 -30932
rect 29317 -31168 29553 -30932
rect 29657 -31168 29893 -30932
rect 29997 -31168 30233 -30932
rect 30317 -31168 30553 -30932
rect 30657 -31168 30893 -30932
rect 30997 -31168 31233 -30932
rect 31317 -31168 31553 -30932
rect 31657 -31168 31893 -30932
rect 31997 -31168 32233 -30932
rect 32317 -31168 32553 -30932
rect 32657 -31168 32893 -30932
rect 32997 -31168 33233 -30932
rect 33317 -31168 33553 -30932
rect 33657 -31168 33893 -30932
rect 33997 -31168 34233 -30932
rect -74443 -31508 -74207 -31272
rect -74443 -31828 -74207 -31592
rect -73443 -31508 -73207 -31272
rect -73443 -31828 -73207 -31592
rect -72443 -31508 -72207 -31272
rect -72443 -31828 -72207 -31592
rect -71443 -31508 -71207 -31272
rect -71443 -31828 -71207 -31592
rect -70443 -31508 -70207 -31272
rect -70443 -31828 -70207 -31592
rect -69443 -31508 -69207 -31272
rect -69443 -31828 -69207 -31592
rect -68443 -31508 -68207 -31272
rect -68443 -31828 -68207 -31592
rect -67443 -31508 -67207 -31272
rect -67443 -31828 -67207 -31592
rect -66443 -31508 -66207 -31272
rect -66443 -31828 -66207 -31592
rect -65443 -31508 -65207 -31272
rect -65443 -31828 -65207 -31592
rect -64443 -31508 -64207 -31272
rect -64443 -31828 -64207 -31592
rect -63443 -31508 -63207 -31272
rect -63443 -31828 -63207 -31592
rect -62443 -31508 -62207 -31272
rect -62443 -31828 -62207 -31592
rect -61443 -31508 -61207 -31272
rect -61443 -31828 -61207 -31592
rect -60443 -31508 -60207 -31272
rect -60443 -31828 -60207 -31592
rect -59443 -31508 -59207 -31272
rect -59443 -31828 -59207 -31592
rect -58443 -31508 -58207 -31272
rect -58443 -31828 -58207 -31592
rect -57443 -31508 -57207 -31272
rect -57443 -31828 -57207 -31592
rect -56443 -31508 -56207 -31272
rect -56443 -31828 -56207 -31592
rect -55443 -31508 -55207 -31272
rect -55443 -31828 -55207 -31592
rect -54443 -31508 -54207 -31272
rect -54443 -31828 -54207 -31592
rect -53443 -31508 -53207 -31272
rect -53443 -31828 -53207 -31592
rect -52443 -31508 -52207 -31272
rect -52443 -31828 -52207 -31592
rect -51443 -31508 -51207 -31272
rect -51443 -31828 -51207 -31592
rect -50443 -31508 -50207 -31272
rect -50443 -31828 -50207 -31592
rect -49443 -31508 -49207 -31272
rect -49443 -31828 -49207 -31592
rect 8657 -31508 8893 -31272
rect 8657 -31828 8893 -31592
rect 9657 -31508 9893 -31272
rect 9657 -31828 9893 -31592
rect 10657 -31508 10893 -31272
rect 10657 -31828 10893 -31592
rect 11657 -31508 11893 -31272
rect 11657 -31828 11893 -31592
rect 12657 -31508 12893 -31272
rect 12657 -31828 12893 -31592
rect 13657 -31508 13893 -31272
rect 13657 -31828 13893 -31592
rect 14657 -31508 14893 -31272
rect 14657 -31828 14893 -31592
rect 15657 -31508 15893 -31272
rect 15657 -31828 15893 -31592
rect 16657 -31508 16893 -31272
rect 16657 -31828 16893 -31592
rect 17657 -31508 17893 -31272
rect 17657 -31828 17893 -31592
rect 18657 -31508 18893 -31272
rect 18657 -31828 18893 -31592
rect 19657 -31508 19893 -31272
rect 19657 -31828 19893 -31592
rect 20657 -31508 20893 -31272
rect 20657 -31828 20893 -31592
rect 21657 -31508 21893 -31272
rect 21657 -31828 21893 -31592
rect 22657 -31508 22893 -31272
rect 22657 -31828 22893 -31592
rect 23657 -31508 23893 -31272
rect 23657 -31828 23893 -31592
rect 24657 -31508 24893 -31272
rect 24657 -31828 24893 -31592
rect 25657 -31508 25893 -31272
rect 25657 -31828 25893 -31592
rect 26657 -31508 26893 -31272
rect 26657 -31828 26893 -31592
rect 27657 -31508 27893 -31272
rect 27657 -31828 27893 -31592
rect 28657 -31508 28893 -31272
rect 28657 -31828 28893 -31592
rect 29657 -31508 29893 -31272
rect 29657 -31828 29893 -31592
rect 30657 -31508 30893 -31272
rect 30657 -31828 30893 -31592
rect 31657 -31508 31893 -31272
rect 31657 -31828 31893 -31592
rect 32657 -31508 32893 -31272
rect 32657 -31828 32893 -31592
rect 33657 -31508 33893 -31272
rect 33657 -31828 33893 -31592
rect -74783 -32168 -74547 -31932
rect -74443 -32168 -74207 -31932
rect -74103 -32168 -73867 -31932
rect -73783 -32168 -73547 -31932
rect -73443 -32168 -73207 -31932
rect -73103 -32168 -72867 -31932
rect -72783 -32168 -72547 -31932
rect -72443 -32168 -72207 -31932
rect -72103 -32168 -71867 -31932
rect -71783 -32168 -71547 -31932
rect -71443 -32168 -71207 -31932
rect -71103 -32168 -70867 -31932
rect -70783 -32168 -70547 -31932
rect -70443 -32168 -70207 -31932
rect -70103 -32168 -69867 -31932
rect -69783 -32168 -69547 -31932
rect -69443 -32168 -69207 -31932
rect -69103 -32168 -68867 -31932
rect -68783 -32168 -68547 -31932
rect -68443 -32168 -68207 -31932
rect -68103 -32168 -67867 -31932
rect -67783 -32168 -67547 -31932
rect -67443 -32168 -67207 -31932
rect -67103 -32168 -66867 -31932
rect -66783 -32168 -66547 -31932
rect -66443 -32168 -66207 -31932
rect -66103 -32168 -65867 -31932
rect -65783 -32168 -65547 -31932
rect -65443 -32168 -65207 -31932
rect -65103 -32168 -64867 -31932
rect -64783 -32168 -64547 -31932
rect -64443 -32168 -64207 -31932
rect -64103 -32168 -63867 -31932
rect -63783 -32168 -63547 -31932
rect -63443 -32168 -63207 -31932
rect -63103 -32168 -62867 -31932
rect -62783 -32168 -62547 -31932
rect -62443 -32168 -62207 -31932
rect -62103 -32168 -61867 -31932
rect -61783 -32168 -61547 -31932
rect -61443 -32168 -61207 -31932
rect -61103 -32168 -60867 -31932
rect -60783 -32168 -60547 -31932
rect -60443 -32168 -60207 -31932
rect -60103 -32168 -59867 -31932
rect -59783 -32168 -59547 -31932
rect -59443 -32168 -59207 -31932
rect -59103 -32168 -58867 -31932
rect -58783 -32168 -58547 -31932
rect -58443 -32168 -58207 -31932
rect -58103 -32168 -57867 -31932
rect -57783 -32168 -57547 -31932
rect -57443 -32168 -57207 -31932
rect -57103 -32168 -56867 -31932
rect -56783 -32168 -56547 -31932
rect -56443 -32168 -56207 -31932
rect -56103 -32168 -55867 -31932
rect -55783 -32168 -55547 -31932
rect -55443 -32168 -55207 -31932
rect -55103 -32168 -54867 -31932
rect -54783 -32168 -54547 -31932
rect -54443 -32168 -54207 -31932
rect -54103 -32168 -53867 -31932
rect -53783 -32168 -53547 -31932
rect -53443 -32168 -53207 -31932
rect -53103 -32168 -52867 -31932
rect -52783 -32168 -52547 -31932
rect -52443 -32168 -52207 -31932
rect -52103 -32168 -51867 -31932
rect -51783 -32168 -51547 -31932
rect -51443 -32168 -51207 -31932
rect -51103 -32168 -50867 -31932
rect -50783 -32168 -50547 -31932
rect -50443 -32168 -50207 -31932
rect -50103 -32168 -49867 -31932
rect -49783 -32168 -49547 -31932
rect -49443 -32168 -49207 -31932
rect -49103 -32168 -48867 -31932
rect 8317 -32168 8553 -31932
rect 8657 -32168 8893 -31932
rect 8997 -32168 9233 -31932
rect 9317 -32168 9553 -31932
rect 9657 -32168 9893 -31932
rect 9997 -32168 10233 -31932
rect 10317 -32168 10553 -31932
rect 10657 -32168 10893 -31932
rect 10997 -32168 11233 -31932
rect 11317 -32168 11553 -31932
rect 11657 -32168 11893 -31932
rect 11997 -32168 12233 -31932
rect 12317 -32168 12553 -31932
rect 12657 -32168 12893 -31932
rect 12997 -32168 13233 -31932
rect 13317 -32168 13553 -31932
rect 13657 -32168 13893 -31932
rect 13997 -32168 14233 -31932
rect 14317 -32168 14553 -31932
rect 14657 -32168 14893 -31932
rect 14997 -32168 15233 -31932
rect 15317 -32168 15553 -31932
rect 15657 -32168 15893 -31932
rect 15997 -32168 16233 -31932
rect 16317 -32168 16553 -31932
rect 16657 -32168 16893 -31932
rect 16997 -32168 17233 -31932
rect 17317 -32168 17553 -31932
rect 17657 -32168 17893 -31932
rect 17997 -32168 18233 -31932
rect 18317 -32168 18553 -31932
rect 18657 -32168 18893 -31932
rect 18997 -32168 19233 -31932
rect 19317 -32168 19553 -31932
rect 19657 -32168 19893 -31932
rect 19997 -32168 20233 -31932
rect 20317 -32168 20553 -31932
rect 20657 -32168 20893 -31932
rect 20997 -32168 21233 -31932
rect 21317 -32168 21553 -31932
rect 21657 -32168 21893 -31932
rect 21997 -32168 22233 -31932
rect 22317 -32168 22553 -31932
rect 22657 -32168 22893 -31932
rect 22997 -32168 23233 -31932
rect 23317 -32168 23553 -31932
rect 23657 -32168 23893 -31932
rect 23997 -32168 24233 -31932
rect 24317 -32168 24553 -31932
rect 24657 -32168 24893 -31932
rect 24997 -32168 25233 -31932
rect 25317 -32168 25553 -31932
rect 25657 -32168 25893 -31932
rect 25997 -32168 26233 -31932
rect 26317 -32168 26553 -31932
rect 26657 -32168 26893 -31932
rect 26997 -32168 27233 -31932
rect 27317 -32168 27553 -31932
rect 27657 -32168 27893 -31932
rect 27997 -32168 28233 -31932
rect 28317 -32168 28553 -31932
rect 28657 -32168 28893 -31932
rect 28997 -32168 29233 -31932
rect 29317 -32168 29553 -31932
rect 29657 -32168 29893 -31932
rect 29997 -32168 30233 -31932
rect 30317 -32168 30553 -31932
rect 30657 -32168 30893 -31932
rect 30997 -32168 31233 -31932
rect 31317 -32168 31553 -31932
rect 31657 -32168 31893 -31932
rect 31997 -32168 32233 -31932
rect 32317 -32168 32553 -31932
rect 32657 -32168 32893 -31932
rect 32997 -32168 33233 -31932
rect 33317 -32168 33553 -31932
rect 33657 -32168 33893 -31932
rect 33997 -32168 34233 -31932
rect -74443 -32508 -74207 -32272
rect -74443 -32828 -74207 -32592
rect -73443 -32508 -73207 -32272
rect -73443 -32828 -73207 -32592
rect -72443 -32508 -72207 -32272
rect -72443 -32828 -72207 -32592
rect -71443 -32508 -71207 -32272
rect -71443 -32828 -71207 -32592
rect -70443 -32508 -70207 -32272
rect -70443 -32828 -70207 -32592
rect -69443 -32508 -69207 -32272
rect -69443 -32828 -69207 -32592
rect -68443 -32508 -68207 -32272
rect -68443 -32828 -68207 -32592
rect -67443 -32508 -67207 -32272
rect -67443 -32828 -67207 -32592
rect -66443 -32508 -66207 -32272
rect -66443 -32828 -66207 -32592
rect -65443 -32508 -65207 -32272
rect -65443 -32828 -65207 -32592
rect -64443 -32508 -64207 -32272
rect -64443 -32828 -64207 -32592
rect -63443 -32508 -63207 -32272
rect -63443 -32828 -63207 -32592
rect -62443 -32508 -62207 -32272
rect -62443 -32828 -62207 -32592
rect -61443 -32508 -61207 -32272
rect -61443 -32828 -61207 -32592
rect -60443 -32508 -60207 -32272
rect -60443 -32828 -60207 -32592
rect -59443 -32508 -59207 -32272
rect -59443 -32828 -59207 -32592
rect -58443 -32508 -58207 -32272
rect -58443 -32828 -58207 -32592
rect -57443 -32508 -57207 -32272
rect -57443 -32828 -57207 -32592
rect -56443 -32508 -56207 -32272
rect -56443 -32828 -56207 -32592
rect -55443 -32508 -55207 -32272
rect -55443 -32828 -55207 -32592
rect -54443 -32508 -54207 -32272
rect -54443 -32828 -54207 -32592
rect -53443 -32508 -53207 -32272
rect -53443 -32828 -53207 -32592
rect -52443 -32508 -52207 -32272
rect -52443 -32828 -52207 -32592
rect -51443 -32508 -51207 -32272
rect -51443 -32828 -51207 -32592
rect -50443 -32508 -50207 -32272
rect -50443 -32828 -50207 -32592
rect -49443 -32508 -49207 -32272
rect -49443 -32828 -49207 -32592
rect -74783 -33168 -74547 -32932
rect -74443 -33168 -74207 -32932
rect -74103 -33168 -73867 -32932
rect -73783 -33168 -73547 -32932
rect -73443 -33168 -73207 -32932
rect -73103 -33168 -72867 -32932
rect -72783 -33168 -72547 -32932
rect -72443 -33168 -72207 -32932
rect -72103 -33168 -71867 -32932
rect -71783 -33168 -71547 -32932
rect -71443 -33168 -71207 -32932
rect -71103 -33168 -70867 -32932
rect -70783 -33168 -70547 -32932
rect -70443 -33168 -70207 -32932
rect -70103 -33168 -69867 -32932
rect -69783 -33168 -69547 -32932
rect -69443 -33168 -69207 -32932
rect -69103 -33168 -68867 -32932
rect -68783 -33168 -68547 -32932
rect -68443 -33168 -68207 -32932
rect -68103 -33168 -67867 -32932
rect -67783 -33168 -67547 -32932
rect -67443 -33168 -67207 -32932
rect -67103 -33168 -66867 -32932
rect -66783 -33168 -66547 -32932
rect -66443 -33168 -66207 -32932
rect -66103 -33168 -65867 -32932
rect -65783 -33168 -65547 -32932
rect -65443 -33168 -65207 -32932
rect -65103 -33168 -64867 -32932
rect -64783 -33168 -64547 -32932
rect -64443 -33168 -64207 -32932
rect -64103 -33168 -63867 -32932
rect -63783 -33168 -63547 -32932
rect -63443 -33168 -63207 -32932
rect -63103 -33168 -62867 -32932
rect -62783 -33168 -62547 -32932
rect -62443 -33168 -62207 -32932
rect -62103 -33168 -61867 -32932
rect -61783 -33168 -61547 -32932
rect -61443 -33168 -61207 -32932
rect -61103 -33168 -60867 -32932
rect -60783 -33168 -60547 -32932
rect -60443 -33168 -60207 -32932
rect -60103 -33168 -59867 -32932
rect -59783 -33168 -59547 -32932
rect -59443 -33168 -59207 -32932
rect -59103 -33168 -58867 -32932
rect -58783 -33168 -58547 -32932
rect -58443 -33168 -58207 -32932
rect -58103 -33168 -57867 -32932
rect -57783 -33168 -57547 -32932
rect -57443 -33168 -57207 -32932
rect -57103 -33168 -56867 -32932
rect -56783 -33168 -56547 -32932
rect -56443 -33168 -56207 -32932
rect -56103 -33168 -55867 -32932
rect -55783 -33168 -55547 -32932
rect -55443 -33168 -55207 -32932
rect -55103 -33168 -54867 -32932
rect -54783 -33168 -54547 -32932
rect -54443 -33168 -54207 -32932
rect -54103 -33168 -53867 -32932
rect -53783 -33168 -53547 -32932
rect -53443 -33168 -53207 -32932
rect -53103 -33168 -52867 -32932
rect -52783 -33168 -52547 -32932
rect -52443 -33168 -52207 -32932
rect -52103 -33168 -51867 -32932
rect -51783 -33168 -51547 -32932
rect -51443 -33168 -51207 -32932
rect -51103 -33168 -50867 -32932
rect -50783 -33168 -50547 -32932
rect -50443 -33168 -50207 -32932
rect -50103 -33168 -49867 -32932
rect -49783 -33168 -49547 -32932
rect -49443 -33168 -49207 -32932
rect -49103 -33168 -48867 -32932
rect -74443 -33508 -74207 -33272
rect -74443 -33828 -74207 -33592
rect -73443 -33508 -73207 -33272
rect -73443 -33828 -73207 -33592
rect -72443 -33508 -72207 -33272
rect -72443 -33828 -72207 -33592
rect -71443 -33508 -71207 -33272
rect -71443 -33828 -71207 -33592
rect -70443 -33508 -70207 -33272
rect -70443 -33828 -70207 -33592
rect -69443 -33508 -69207 -33272
rect -69443 -33828 -69207 -33592
rect -68443 -33508 -68207 -33272
rect -68443 -33828 -68207 -33592
rect -67443 -33508 -67207 -33272
rect -67443 -33828 -67207 -33592
rect -66443 -33508 -66207 -33272
rect -66443 -33828 -66207 -33592
rect -65443 -33508 -65207 -33272
rect -65443 -33828 -65207 -33592
rect -64443 -33508 -64207 -33272
rect -64443 -33828 -64207 -33592
rect -63443 -33508 -63207 -33272
rect -63443 -33828 -63207 -33592
rect -62443 -33508 -62207 -33272
rect -62443 -33828 -62207 -33592
rect -61443 -33508 -61207 -33272
rect -61443 -33828 -61207 -33592
rect -60443 -33508 -60207 -33272
rect -60443 -33828 -60207 -33592
rect -59443 -33508 -59207 -33272
rect -59443 -33828 -59207 -33592
rect -58443 -33508 -58207 -33272
rect -58443 -33828 -58207 -33592
rect -57443 -33508 -57207 -33272
rect -57443 -33828 -57207 -33592
rect -56443 -33508 -56207 -33272
rect -56443 -33828 -56207 -33592
rect -55443 -33508 -55207 -33272
rect -55443 -33828 -55207 -33592
rect -54443 -33508 -54207 -33272
rect -54443 -33828 -54207 -33592
rect -53443 -33508 -53207 -33272
rect -53443 -33828 -53207 -33592
rect -52443 -33508 -52207 -33272
rect -52443 -33828 -52207 -33592
rect -51443 -33508 -51207 -33272
rect -51443 -33828 -51207 -33592
rect -50443 -33508 -50207 -33272
rect -50443 -33828 -50207 -33592
rect -49443 -33508 -49207 -33272
rect -49443 -33828 -49207 -33592
rect -74783 -34168 -74547 -33932
rect -74443 -34168 -74207 -33932
rect -74103 -34168 -73867 -33932
rect -73783 -34168 -73547 -33932
rect -73443 -34168 -73207 -33932
rect -73103 -34168 -72867 -33932
rect -72783 -34168 -72547 -33932
rect -72443 -34168 -72207 -33932
rect -72103 -34168 -71867 -33932
rect -71783 -34168 -71547 -33932
rect -71443 -34168 -71207 -33932
rect -71103 -34168 -70867 -33932
rect -70783 -34168 -70547 -33932
rect -70443 -34168 -70207 -33932
rect -70103 -34168 -69867 -33932
rect -69783 -34168 -69547 -33932
rect -69443 -34168 -69207 -33932
rect -69103 -34168 -68867 -33932
rect -68783 -34168 -68547 -33932
rect -68443 -34168 -68207 -33932
rect -68103 -34168 -67867 -33932
rect -67783 -34168 -67547 -33932
rect -67443 -34168 -67207 -33932
rect -67103 -34168 -66867 -33932
rect -66783 -34168 -66547 -33932
rect -66443 -34168 -66207 -33932
rect -66103 -34168 -65867 -33932
rect -65783 -34168 -65547 -33932
rect -65443 -34168 -65207 -33932
rect -65103 -34168 -64867 -33932
rect -64783 -34168 -64547 -33932
rect -64443 -34168 -64207 -33932
rect -64103 -34168 -63867 -33932
rect -63783 -34168 -63547 -33932
rect -63443 -34168 -63207 -33932
rect -63103 -34168 -62867 -33932
rect -62783 -34168 -62547 -33932
rect -62443 -34168 -62207 -33932
rect -62103 -34168 -61867 -33932
rect -61783 -34168 -61547 -33932
rect -61443 -34168 -61207 -33932
rect -61103 -34168 -60867 -33932
rect -60783 -34168 -60547 -33932
rect -60443 -34168 -60207 -33932
rect -60103 -34168 -59867 -33932
rect -59783 -34168 -59547 -33932
rect -59443 -34168 -59207 -33932
rect -59103 -34168 -58867 -33932
rect -58783 -34168 -58547 -33932
rect -58443 -34168 -58207 -33932
rect -58103 -34168 -57867 -33932
rect -57783 -34168 -57547 -33932
rect -57443 -34168 -57207 -33932
rect -57103 -34168 -56867 -33932
rect -56783 -34168 -56547 -33932
rect -56443 -34168 -56207 -33932
rect -56103 -34168 -55867 -33932
rect -55783 -34168 -55547 -33932
rect -55443 -34168 -55207 -33932
rect -55103 -34168 -54867 -33932
rect -54783 -34168 -54547 -33932
rect -54443 -34168 -54207 -33932
rect -54103 -34168 -53867 -33932
rect -53783 -34168 -53547 -33932
rect -53443 -34168 -53207 -33932
rect -53103 -34168 -52867 -33932
rect -52783 -34168 -52547 -33932
rect -52443 -34168 -52207 -33932
rect -52103 -34168 -51867 -33932
rect -51783 -34168 -51547 -33932
rect -51443 -34168 -51207 -33932
rect -51103 -34168 -50867 -33932
rect -50783 -34168 -50547 -33932
rect -50443 -34168 -50207 -33932
rect -50103 -34168 -49867 -33932
rect -49783 -34168 -49547 -33932
rect -49443 -34168 -49207 -33932
rect -49103 -34168 -48867 -33932
rect -74443 -34508 -74207 -34272
rect -74443 -34828 -74207 -34592
rect -73443 -34508 -73207 -34272
rect -73443 -34828 -73207 -34592
rect -72443 -34508 -72207 -34272
rect -72443 -34828 -72207 -34592
rect -71443 -34508 -71207 -34272
rect -71443 -34828 -71207 -34592
rect -70443 -34508 -70207 -34272
rect -70443 -34828 -70207 -34592
rect -69443 -34508 -69207 -34272
rect -69443 -34828 -69207 -34592
rect -68443 -34508 -68207 -34272
rect -68443 -34828 -68207 -34592
rect -67443 -34508 -67207 -34272
rect -67443 -34828 -67207 -34592
rect -66443 -34508 -66207 -34272
rect -66443 -34828 -66207 -34592
rect -65443 -34508 -65207 -34272
rect -65443 -34828 -65207 -34592
rect -64443 -34508 -64207 -34272
rect -64443 -34828 -64207 -34592
rect -63443 -34508 -63207 -34272
rect -63443 -34828 -63207 -34592
rect -62443 -34508 -62207 -34272
rect -62443 -34828 -62207 -34592
rect -61443 -34508 -61207 -34272
rect -61443 -34828 -61207 -34592
rect -60443 -34508 -60207 -34272
rect -60443 -34828 -60207 -34592
rect -59443 -34508 -59207 -34272
rect -59443 -34828 -59207 -34592
rect -58443 -34508 -58207 -34272
rect -58443 -34828 -58207 -34592
rect -57443 -34508 -57207 -34272
rect -57443 -34828 -57207 -34592
rect -56443 -34508 -56207 -34272
rect -56443 -34828 -56207 -34592
rect -55443 -34508 -55207 -34272
rect -55443 -34828 -55207 -34592
rect -54443 -34508 -54207 -34272
rect -54443 -34828 -54207 -34592
rect -53443 -34508 -53207 -34272
rect -53443 -34828 -53207 -34592
rect -52443 -34508 -52207 -34272
rect -52443 -34828 -52207 -34592
rect -51443 -34508 -51207 -34272
rect -51443 -34828 -51207 -34592
rect -50443 -34508 -50207 -34272
rect -50443 -34828 -50207 -34592
rect -49443 -34508 -49207 -34272
rect -49443 -34828 -49207 -34592
rect -74783 -35168 -74547 -34932
rect -74443 -35168 -74207 -34932
rect -74103 -35168 -73867 -34932
rect -73783 -35168 -73547 -34932
rect -73443 -35168 -73207 -34932
rect -73103 -35168 -72867 -34932
rect -72783 -35168 -72547 -34932
rect -72443 -35168 -72207 -34932
rect -72103 -35168 -71867 -34932
rect -71783 -35168 -71547 -34932
rect -71443 -35168 -71207 -34932
rect -71103 -35168 -70867 -34932
rect -70783 -35168 -70547 -34932
rect -70443 -35168 -70207 -34932
rect -70103 -35168 -69867 -34932
rect -69783 -35168 -69547 -34932
rect -69443 -35168 -69207 -34932
rect -69103 -35168 -68867 -34932
rect -68783 -35168 -68547 -34932
rect -68443 -35168 -68207 -34932
rect -68103 -35168 -67867 -34932
rect -67783 -35168 -67547 -34932
rect -67443 -35168 -67207 -34932
rect -67103 -35168 -66867 -34932
rect -66783 -35168 -66547 -34932
rect -66443 -35168 -66207 -34932
rect -66103 -35168 -65867 -34932
rect -65783 -35168 -65547 -34932
rect -65443 -35168 -65207 -34932
rect -65103 -35168 -64867 -34932
rect -64783 -35168 -64547 -34932
rect -64443 -35168 -64207 -34932
rect -64103 -35168 -63867 -34932
rect -63783 -35168 -63547 -34932
rect -63443 -35168 -63207 -34932
rect -63103 -35168 -62867 -34932
rect -62783 -35168 -62547 -34932
rect -62443 -35168 -62207 -34932
rect -62103 -35168 -61867 -34932
rect -61783 -35168 -61547 -34932
rect -61443 -35168 -61207 -34932
rect -61103 -35168 -60867 -34932
rect -60783 -35168 -60547 -34932
rect -60443 -35168 -60207 -34932
rect -60103 -35168 -59867 -34932
rect -59783 -35168 -59547 -34932
rect -59443 -35168 -59207 -34932
rect -59103 -35168 -58867 -34932
rect -58783 -35168 -58547 -34932
rect -58443 -35168 -58207 -34932
rect -58103 -35168 -57867 -34932
rect -57783 -35168 -57547 -34932
rect -57443 -35168 -57207 -34932
rect -57103 -35168 -56867 -34932
rect -56783 -35168 -56547 -34932
rect -56443 -35168 -56207 -34932
rect -56103 -35168 -55867 -34932
rect -55783 -35168 -55547 -34932
rect -55443 -35168 -55207 -34932
rect -55103 -35168 -54867 -34932
rect -54783 -35168 -54547 -34932
rect -54443 -35168 -54207 -34932
rect -54103 -35168 -53867 -34932
rect -53783 -35168 -53547 -34932
rect -53443 -35168 -53207 -34932
rect -53103 -35168 -52867 -34932
rect -52783 -35168 -52547 -34932
rect -52443 -35168 -52207 -34932
rect -52103 -35168 -51867 -34932
rect -51783 -35168 -51547 -34932
rect -51443 -35168 -51207 -34932
rect -51103 -35168 -50867 -34932
rect -50783 -35168 -50547 -34932
rect -50443 -35168 -50207 -34932
rect -50103 -35168 -49867 -34932
rect -49783 -35168 -49547 -34932
rect -49443 -35168 -49207 -34932
rect -49103 -35168 -48867 -34932
rect -74443 -35508 -74207 -35272
rect -74443 -35828 -74207 -35592
rect -73443 -35508 -73207 -35272
rect -73443 -35828 -73207 -35592
rect -72443 -35508 -72207 -35272
rect -72443 -35828 -72207 -35592
rect -71443 -35508 -71207 -35272
rect -71443 -35828 -71207 -35592
rect -70443 -35508 -70207 -35272
rect -70443 -35828 -70207 -35592
rect -69443 -35508 -69207 -35272
rect -69443 -35828 -69207 -35592
rect -68443 -35508 -68207 -35272
rect -68443 -35828 -68207 -35592
rect -67443 -35508 -67207 -35272
rect -67443 -35828 -67207 -35592
rect -66443 -35508 -66207 -35272
rect -66443 -35828 -66207 -35592
rect -65443 -35508 -65207 -35272
rect -65443 -35828 -65207 -35592
rect -64443 -35508 -64207 -35272
rect -64443 -35828 -64207 -35592
rect -63443 -35508 -63207 -35272
rect -63443 -35828 -63207 -35592
rect -62443 -35508 -62207 -35272
rect -62443 -35828 -62207 -35592
rect -61443 -35508 -61207 -35272
rect -61443 -35828 -61207 -35592
rect -60443 -35508 -60207 -35272
rect -60443 -35828 -60207 -35592
rect -59443 -35508 -59207 -35272
rect -59443 -35828 -59207 -35592
rect -58443 -35508 -58207 -35272
rect -58443 -35828 -58207 -35592
rect -57443 -35508 -57207 -35272
rect -57443 -35828 -57207 -35592
rect -56443 -35508 -56207 -35272
rect -56443 -35828 -56207 -35592
rect -55443 -35508 -55207 -35272
rect -55443 -35828 -55207 -35592
rect -54443 -35508 -54207 -35272
rect -54443 -35828 -54207 -35592
rect -53443 -35508 -53207 -35272
rect -53443 -35828 -53207 -35592
rect -52443 -35508 -52207 -35272
rect -52443 -35828 -52207 -35592
rect -51443 -35508 -51207 -35272
rect -51443 -35828 -51207 -35592
rect -50443 -35508 -50207 -35272
rect -50443 -35828 -50207 -35592
rect -49443 -35508 -49207 -35272
rect -49443 -35828 -49207 -35592
rect -74783 -36168 -74547 -35932
rect -74443 -36168 -74207 -35932
rect -74103 -36168 -73867 -35932
rect -73783 -36168 -73547 -35932
rect -73443 -36168 -73207 -35932
rect -73103 -36168 -72867 -35932
rect -72783 -36168 -72547 -35932
rect -72443 -36168 -72207 -35932
rect -72103 -36168 -71867 -35932
rect -71783 -36168 -71547 -35932
rect -71443 -36168 -71207 -35932
rect -71103 -36168 -70867 -35932
rect -70783 -36168 -70547 -35932
rect -70443 -36168 -70207 -35932
rect -70103 -36168 -69867 -35932
rect -69783 -36168 -69547 -35932
rect -69443 -36168 -69207 -35932
rect -69103 -36168 -68867 -35932
rect -68783 -36168 -68547 -35932
rect -68443 -36168 -68207 -35932
rect -68103 -36168 -67867 -35932
rect -67783 -36168 -67547 -35932
rect -67443 -36168 -67207 -35932
rect -67103 -36168 -66867 -35932
rect -66783 -36168 -66547 -35932
rect -66443 -36168 -66207 -35932
rect -66103 -36168 -65867 -35932
rect -65783 -36168 -65547 -35932
rect -65443 -36168 -65207 -35932
rect -65103 -36168 -64867 -35932
rect -64783 -36168 -64547 -35932
rect -64443 -36168 -64207 -35932
rect -64103 -36168 -63867 -35932
rect -63783 -36168 -63547 -35932
rect -63443 -36168 -63207 -35932
rect -63103 -36168 -62867 -35932
rect -62783 -36168 -62547 -35932
rect -62443 -36168 -62207 -35932
rect -62103 -36168 -61867 -35932
rect -61783 -36168 -61547 -35932
rect -61443 -36168 -61207 -35932
rect -61103 -36168 -60867 -35932
rect -60783 -36168 -60547 -35932
rect -60443 -36168 -60207 -35932
rect -60103 -36168 -59867 -35932
rect -59783 -36168 -59547 -35932
rect -59443 -36168 -59207 -35932
rect -59103 -36168 -58867 -35932
rect -58783 -36168 -58547 -35932
rect -58443 -36168 -58207 -35932
rect -58103 -36168 -57867 -35932
rect -57783 -36168 -57547 -35932
rect -57443 -36168 -57207 -35932
rect -57103 -36168 -56867 -35932
rect -56783 -36168 -56547 -35932
rect -56443 -36168 -56207 -35932
rect -56103 -36168 -55867 -35932
rect -55783 -36168 -55547 -35932
rect -55443 -36168 -55207 -35932
rect -55103 -36168 -54867 -35932
rect -54783 -36168 -54547 -35932
rect -54443 -36168 -54207 -35932
rect -54103 -36168 -53867 -35932
rect -53783 -36168 -53547 -35932
rect -53443 -36168 -53207 -35932
rect -53103 -36168 -52867 -35932
rect -52783 -36168 -52547 -35932
rect -52443 -36168 -52207 -35932
rect -52103 -36168 -51867 -35932
rect -51783 -36168 -51547 -35932
rect -51443 -36168 -51207 -35932
rect -51103 -36168 -50867 -35932
rect -50783 -36168 -50547 -35932
rect -50443 -36168 -50207 -35932
rect -50103 -36168 -49867 -35932
rect -49783 -36168 -49547 -35932
rect -49443 -36168 -49207 -35932
rect -49103 -36168 -48867 -35932
rect -74443 -36508 -74207 -36272
rect -74443 -36828 -74207 -36592
rect -73443 -36508 -73207 -36272
rect -73443 -36828 -73207 -36592
rect -72443 -36508 -72207 -36272
rect -72443 -36828 -72207 -36592
rect -71443 -36508 -71207 -36272
rect -71443 -36828 -71207 -36592
rect -70443 -36508 -70207 -36272
rect -70443 -36828 -70207 -36592
rect -69443 -36508 -69207 -36272
rect -69443 -36828 -69207 -36592
rect -68443 -36508 -68207 -36272
rect -68443 -36828 -68207 -36592
rect -67443 -36508 -67207 -36272
rect -67443 -36828 -67207 -36592
rect -66443 -36508 -66207 -36272
rect -66443 -36828 -66207 -36592
rect -65443 -36508 -65207 -36272
rect -65443 -36828 -65207 -36592
rect -64443 -36508 -64207 -36272
rect -64443 -36828 -64207 -36592
rect -63443 -36508 -63207 -36272
rect -63443 -36828 -63207 -36592
rect -62443 -36508 -62207 -36272
rect -62443 -36828 -62207 -36592
rect -61443 -36508 -61207 -36272
rect -61443 -36828 -61207 -36592
rect -60443 -36508 -60207 -36272
rect -60443 -36828 -60207 -36592
rect -59443 -36508 -59207 -36272
rect -59443 -36828 -59207 -36592
rect -58443 -36508 -58207 -36272
rect -58443 -36828 -58207 -36592
rect -57443 -36508 -57207 -36272
rect -57443 -36828 -57207 -36592
rect -56443 -36508 -56207 -36272
rect -56443 -36828 -56207 -36592
rect -55443 -36508 -55207 -36272
rect -55443 -36828 -55207 -36592
rect -54443 -36508 -54207 -36272
rect -54443 -36828 -54207 -36592
rect -53443 -36508 -53207 -36272
rect -53443 -36828 -53207 -36592
rect -52443 -36508 -52207 -36272
rect -52443 -36828 -52207 -36592
rect -51443 -36508 -51207 -36272
rect -51443 -36828 -51207 -36592
rect -50443 -36508 -50207 -36272
rect -50443 -36828 -50207 -36592
rect -49443 -36508 -49207 -36272
rect -49443 -36828 -49207 -36592
rect -74783 -37168 -74547 -36932
rect -74443 -37168 -74207 -36932
rect -74103 -37168 -73867 -36932
rect -73783 -37168 -73547 -36932
rect -73443 -37168 -73207 -36932
rect -73103 -37168 -72867 -36932
rect -72783 -37168 -72547 -36932
rect -72443 -37168 -72207 -36932
rect -72103 -37168 -71867 -36932
rect -71783 -37168 -71547 -36932
rect -71443 -37168 -71207 -36932
rect -71103 -37168 -70867 -36932
rect -70783 -37168 -70547 -36932
rect -70443 -37168 -70207 -36932
rect -70103 -37168 -69867 -36932
rect -69783 -37168 -69547 -36932
rect -69443 -37168 -69207 -36932
rect -69103 -37168 -68867 -36932
rect -68783 -37168 -68547 -36932
rect -68443 -37168 -68207 -36932
rect -68103 -37168 -67867 -36932
rect -67783 -37168 -67547 -36932
rect -67443 -37168 -67207 -36932
rect -67103 -37168 -66867 -36932
rect -66783 -37168 -66547 -36932
rect -66443 -37168 -66207 -36932
rect -66103 -37168 -65867 -36932
rect -65783 -37168 -65547 -36932
rect -65443 -37168 -65207 -36932
rect -65103 -37168 -64867 -36932
rect -64783 -37168 -64547 -36932
rect -64443 -37168 -64207 -36932
rect -64103 -37168 -63867 -36932
rect -63783 -37168 -63547 -36932
rect -63443 -37168 -63207 -36932
rect -63103 -37168 -62867 -36932
rect -62783 -37168 -62547 -36932
rect -62443 -37168 -62207 -36932
rect -62103 -37168 -61867 -36932
rect -61783 -37168 -61547 -36932
rect -61443 -37168 -61207 -36932
rect -61103 -37168 -60867 -36932
rect -60783 -37168 -60547 -36932
rect -60443 -37168 -60207 -36932
rect -60103 -37168 -59867 -36932
rect -59783 -37168 -59547 -36932
rect -59443 -37168 -59207 -36932
rect -59103 -37168 -58867 -36932
rect -58783 -37168 -58547 -36932
rect -58443 -37168 -58207 -36932
rect -58103 -37168 -57867 -36932
rect -57783 -37168 -57547 -36932
rect -57443 -37168 -57207 -36932
rect -57103 -37168 -56867 -36932
rect -56783 -37168 -56547 -36932
rect -56443 -37168 -56207 -36932
rect -56103 -37168 -55867 -36932
rect -55783 -37168 -55547 -36932
rect -55443 -37168 -55207 -36932
rect -55103 -37168 -54867 -36932
rect -54783 -37168 -54547 -36932
rect -54443 -37168 -54207 -36932
rect -54103 -37168 -53867 -36932
rect -53783 -37168 -53547 -36932
rect -53443 -37168 -53207 -36932
rect -53103 -37168 -52867 -36932
rect -52783 -37168 -52547 -36932
rect -52443 -37168 -52207 -36932
rect -52103 -37168 -51867 -36932
rect -51783 -37168 -51547 -36932
rect -51443 -37168 -51207 -36932
rect -51103 -37168 -50867 -36932
rect -50783 -37168 -50547 -36932
rect -50443 -37168 -50207 -36932
rect -50103 -37168 -49867 -36932
rect -49783 -37168 -49547 -36932
rect -49443 -37168 -49207 -36932
rect -49103 -37168 -48867 -36932
rect -74443 -37508 -74207 -37272
rect -74443 -37828 -74207 -37592
rect -73443 -37508 -73207 -37272
rect -73443 -37828 -73207 -37592
rect -72443 -37508 -72207 -37272
rect -72443 -37828 -72207 -37592
rect -71443 -37508 -71207 -37272
rect -71443 -37828 -71207 -37592
rect -70443 -37508 -70207 -37272
rect -70443 -37828 -70207 -37592
rect -69443 -37508 -69207 -37272
rect -69443 -37828 -69207 -37592
rect -68443 -37508 -68207 -37272
rect -68443 -37828 -68207 -37592
rect -67443 -37508 -67207 -37272
rect -67443 -37828 -67207 -37592
rect -66443 -37508 -66207 -37272
rect -66443 -37828 -66207 -37592
rect -65443 -37508 -65207 -37272
rect -65443 -37828 -65207 -37592
rect -64443 -37508 -64207 -37272
rect -64443 -37828 -64207 -37592
rect -63443 -37508 -63207 -37272
rect -63443 -37828 -63207 -37592
rect -62443 -37508 -62207 -37272
rect -62443 -37828 -62207 -37592
rect -61443 -37508 -61207 -37272
rect -61443 -37828 -61207 -37592
rect -60443 -37508 -60207 -37272
rect -60443 -37828 -60207 -37592
rect -59443 -37508 -59207 -37272
rect -59443 -37828 -59207 -37592
rect -58443 -37508 -58207 -37272
rect -58443 -37828 -58207 -37592
rect -57443 -37508 -57207 -37272
rect -57443 -37828 -57207 -37592
rect -56443 -37508 -56207 -37272
rect -56443 -37828 -56207 -37592
rect -55443 -37508 -55207 -37272
rect -55443 -37828 -55207 -37592
rect -54443 -37508 -54207 -37272
rect -54443 -37828 -54207 -37592
rect -53443 -37508 -53207 -37272
rect -53443 -37828 -53207 -37592
rect -52443 -37508 -52207 -37272
rect -52443 -37828 -52207 -37592
rect -51443 -37508 -51207 -37272
rect -51443 -37828 -51207 -37592
rect -50443 -37508 -50207 -37272
rect -50443 -37828 -50207 -37592
rect -49443 -37508 -49207 -37272
rect -49443 -37828 -49207 -37592
rect -74783 -38168 -74547 -37932
rect -74443 -38168 -74207 -37932
rect -74103 -38168 -73867 -37932
rect -73783 -38168 -73547 -37932
rect -73443 -38168 -73207 -37932
rect -73103 -38168 -72867 -37932
rect -72783 -38168 -72547 -37932
rect -72443 -38168 -72207 -37932
rect -72103 -38168 -71867 -37932
rect -71783 -38168 -71547 -37932
rect -71443 -38168 -71207 -37932
rect -71103 -38168 -70867 -37932
rect -70783 -38168 -70547 -37932
rect -70443 -38168 -70207 -37932
rect -70103 -38168 -69867 -37932
rect -69783 -38168 -69547 -37932
rect -69443 -38168 -69207 -37932
rect -69103 -38168 -68867 -37932
rect -68783 -38168 -68547 -37932
rect -68443 -38168 -68207 -37932
rect -68103 -38168 -67867 -37932
rect -67783 -38168 -67547 -37932
rect -67443 -38168 -67207 -37932
rect -67103 -38168 -66867 -37932
rect -66783 -38168 -66547 -37932
rect -66443 -38168 -66207 -37932
rect -66103 -38168 -65867 -37932
rect -65783 -38168 -65547 -37932
rect -65443 -38168 -65207 -37932
rect -65103 -38168 -64867 -37932
rect -64783 -38168 -64547 -37932
rect -64443 -38168 -64207 -37932
rect -64103 -38168 -63867 -37932
rect -63783 -38168 -63547 -37932
rect -63443 -38168 -63207 -37932
rect -63103 -38168 -62867 -37932
rect -62783 -38168 -62547 -37932
rect -62443 -38168 -62207 -37932
rect -62103 -38168 -61867 -37932
rect -61783 -38168 -61547 -37932
rect -61443 -38168 -61207 -37932
rect -61103 -38168 -60867 -37932
rect -60783 -38168 -60547 -37932
rect -60443 -38168 -60207 -37932
rect -60103 -38168 -59867 -37932
rect -59783 -38168 -59547 -37932
rect -59443 -38168 -59207 -37932
rect -59103 -38168 -58867 -37932
rect -58783 -38168 -58547 -37932
rect -58443 -38168 -58207 -37932
rect -58103 -38168 -57867 -37932
rect -57783 -38168 -57547 -37932
rect -57443 -38168 -57207 -37932
rect -57103 -38168 -56867 -37932
rect -56783 -38168 -56547 -37932
rect -56443 -38168 -56207 -37932
rect -56103 -38168 -55867 -37932
rect -55783 -38168 -55547 -37932
rect -55443 -38168 -55207 -37932
rect -55103 -38168 -54867 -37932
rect -54783 -38168 -54547 -37932
rect -54443 -38168 -54207 -37932
rect -54103 -38168 -53867 -37932
rect -53783 -38168 -53547 -37932
rect -53443 -38168 -53207 -37932
rect -53103 -38168 -52867 -37932
rect -52783 -38168 -52547 -37932
rect -52443 -38168 -52207 -37932
rect -52103 -38168 -51867 -37932
rect -51783 -38168 -51547 -37932
rect -51443 -38168 -51207 -37932
rect -51103 -38168 -50867 -37932
rect -50783 -38168 -50547 -37932
rect -50443 -38168 -50207 -37932
rect -50103 -38168 -49867 -37932
rect -49783 -38168 -49547 -37932
rect -49443 -38168 -49207 -37932
rect -49103 -38168 -48867 -37932
rect -74443 -38508 -74207 -38272
rect -74443 -38828 -74207 -38592
rect -73443 -38508 -73207 -38272
rect -73443 -38828 -73207 -38592
rect -72443 -38508 -72207 -38272
rect -72443 -38828 -72207 -38592
rect -71443 -38508 -71207 -38272
rect -71443 -38828 -71207 -38592
rect -70443 -38508 -70207 -38272
rect -70443 -38828 -70207 -38592
rect -69443 -38508 -69207 -38272
rect -69443 -38828 -69207 -38592
rect -68443 -38508 -68207 -38272
rect -68443 -38828 -68207 -38592
rect -67443 -38508 -67207 -38272
rect -67443 -38828 -67207 -38592
rect -66443 -38508 -66207 -38272
rect -66443 -38828 -66207 -38592
rect -65443 -38508 -65207 -38272
rect -65443 -38828 -65207 -38592
rect -64443 -38508 -64207 -38272
rect -64443 -38828 -64207 -38592
rect -63443 -38508 -63207 -38272
rect -63443 -38828 -63207 -38592
rect -62443 -38508 -62207 -38272
rect -62443 -38828 -62207 -38592
rect -61443 -38508 -61207 -38272
rect -61443 -38828 -61207 -38592
rect -60443 -38508 -60207 -38272
rect -60443 -38828 -60207 -38592
rect -59443 -38508 -59207 -38272
rect -59443 -38828 -59207 -38592
rect -58443 -38508 -58207 -38272
rect -58443 -38828 -58207 -38592
rect -57443 -38508 -57207 -38272
rect -57443 -38828 -57207 -38592
rect -56443 -38508 -56207 -38272
rect -56443 -38828 -56207 -38592
rect -55443 -38508 -55207 -38272
rect -55443 -38828 -55207 -38592
rect -54443 -38508 -54207 -38272
rect -54443 -38828 -54207 -38592
rect -53443 -38508 -53207 -38272
rect -53443 -38828 -53207 -38592
rect -52443 -38508 -52207 -38272
rect -52443 -38828 -52207 -38592
rect -51443 -38508 -51207 -38272
rect -51443 -38828 -51207 -38592
rect -50443 -38508 -50207 -38272
rect -50443 -38828 -50207 -38592
rect -49443 -38508 -49207 -38272
rect -49443 -38828 -49207 -38592
rect -74783 -39168 -74547 -38932
rect -74443 -39168 -74207 -38932
rect -74103 -39168 -73867 -38932
rect -73783 -39168 -73547 -38932
rect -73443 -39168 -73207 -38932
rect -73103 -39168 -72867 -38932
rect -72783 -39168 -72547 -38932
rect -72443 -39168 -72207 -38932
rect -72103 -39168 -71867 -38932
rect -71783 -39168 -71547 -38932
rect -71443 -39168 -71207 -38932
rect -71103 -39168 -70867 -38932
rect -70783 -39168 -70547 -38932
rect -70443 -39168 -70207 -38932
rect -70103 -39168 -69867 -38932
rect -69783 -39168 -69547 -38932
rect -69443 -39168 -69207 -38932
rect -69103 -39168 -68867 -38932
rect -68783 -39168 -68547 -38932
rect -68443 -39168 -68207 -38932
rect -68103 -39168 -67867 -38932
rect -67783 -39168 -67547 -38932
rect -67443 -39168 -67207 -38932
rect -67103 -39168 -66867 -38932
rect -66783 -39168 -66547 -38932
rect -66443 -39168 -66207 -38932
rect -66103 -39168 -65867 -38932
rect -65783 -39168 -65547 -38932
rect -65443 -39168 -65207 -38932
rect -65103 -39168 -64867 -38932
rect -64783 -39168 -64547 -38932
rect -64443 -39168 -64207 -38932
rect -64103 -39168 -63867 -38932
rect -63783 -39168 -63547 -38932
rect -63443 -39168 -63207 -38932
rect -63103 -39168 -62867 -38932
rect -62783 -39168 -62547 -38932
rect -62443 -39168 -62207 -38932
rect -62103 -39168 -61867 -38932
rect -61783 -39168 -61547 -38932
rect -61443 -39168 -61207 -38932
rect -61103 -39168 -60867 -38932
rect -60783 -39168 -60547 -38932
rect -60443 -39168 -60207 -38932
rect -60103 -39168 -59867 -38932
rect -59783 -39168 -59547 -38932
rect -59443 -39168 -59207 -38932
rect -59103 -39168 -58867 -38932
rect -58783 -39168 -58547 -38932
rect -58443 -39168 -58207 -38932
rect -58103 -39168 -57867 -38932
rect -57783 -39168 -57547 -38932
rect -57443 -39168 -57207 -38932
rect -57103 -39168 -56867 -38932
rect -56783 -39168 -56547 -38932
rect -56443 -39168 -56207 -38932
rect -56103 -39168 -55867 -38932
rect -55783 -39168 -55547 -38932
rect -55443 -39168 -55207 -38932
rect -55103 -39168 -54867 -38932
rect -54783 -39168 -54547 -38932
rect -54443 -39168 -54207 -38932
rect -54103 -39168 -53867 -38932
rect -53783 -39168 -53547 -38932
rect -53443 -39168 -53207 -38932
rect -53103 -39168 -52867 -38932
rect -52783 -39168 -52547 -38932
rect -52443 -39168 -52207 -38932
rect -52103 -39168 -51867 -38932
rect -51783 -39168 -51547 -38932
rect -51443 -39168 -51207 -38932
rect -51103 -39168 -50867 -38932
rect -50783 -39168 -50547 -38932
rect -50443 -39168 -50207 -38932
rect -50103 -39168 -49867 -38932
rect -49783 -39168 -49547 -38932
rect -49443 -39168 -49207 -38932
rect -49103 -39168 -48867 -38932
rect -74443 -39508 -74207 -39272
rect -74443 -39828 -74207 -39592
rect -73443 -39508 -73207 -39272
rect -73443 -39828 -73207 -39592
rect -72443 -39508 -72207 -39272
rect -72443 -39828 -72207 -39592
rect -71443 -39508 -71207 -39272
rect -71443 -39828 -71207 -39592
rect -70443 -39508 -70207 -39272
rect -70443 -39828 -70207 -39592
rect -69443 -39508 -69207 -39272
rect -69443 -39828 -69207 -39592
rect -68443 -39508 -68207 -39272
rect -68443 -39828 -68207 -39592
rect -67443 -39508 -67207 -39272
rect -67443 -39828 -67207 -39592
rect -66443 -39508 -66207 -39272
rect -66443 -39828 -66207 -39592
rect -65443 -39508 -65207 -39272
rect -65443 -39828 -65207 -39592
rect -64443 -39508 -64207 -39272
rect -64443 -39828 -64207 -39592
rect -63443 -39508 -63207 -39272
rect -63443 -39828 -63207 -39592
rect -62443 -39508 -62207 -39272
rect -62443 -39828 -62207 -39592
rect -61443 -39508 -61207 -39272
rect -61443 -39828 -61207 -39592
rect -60443 -39508 -60207 -39272
rect -60443 -39828 -60207 -39592
rect -59443 -39508 -59207 -39272
rect -59443 -39828 -59207 -39592
rect -58443 -39508 -58207 -39272
rect -58443 -39828 -58207 -39592
rect -57443 -39508 -57207 -39272
rect -57443 -39828 -57207 -39592
rect -56443 -39508 -56207 -39272
rect -56443 -39828 -56207 -39592
rect -55443 -39508 -55207 -39272
rect -55443 -39828 -55207 -39592
rect -54443 -39508 -54207 -39272
rect -54443 -39828 -54207 -39592
rect -53443 -39508 -53207 -39272
rect -53443 -39828 -53207 -39592
rect -52443 -39508 -52207 -39272
rect -52443 -39828 -52207 -39592
rect -51443 -39508 -51207 -39272
rect -51443 -39828 -51207 -39592
rect -50443 -39508 -50207 -39272
rect -50443 -39828 -50207 -39592
rect -49443 -39508 -49207 -39272
rect -49443 -39828 -49207 -39592
rect -74783 -40168 -74547 -39932
rect -74443 -40168 -74207 -39932
rect -74103 -40168 -73867 -39932
rect -73783 -40168 -73547 -39932
rect -73443 -40168 -73207 -39932
rect -73103 -40168 -72867 -39932
rect -72783 -40168 -72547 -39932
rect -72443 -40168 -72207 -39932
rect -72103 -40168 -71867 -39932
rect -71783 -40168 -71547 -39932
rect -71443 -40168 -71207 -39932
rect -71103 -40168 -70867 -39932
rect -70783 -40168 -70547 -39932
rect -70443 -40168 -70207 -39932
rect -70103 -40168 -69867 -39932
rect -69783 -40168 -69547 -39932
rect -69443 -40168 -69207 -39932
rect -69103 -40168 -68867 -39932
rect -68783 -40168 -68547 -39932
rect -68443 -40168 -68207 -39932
rect -68103 -40168 -67867 -39932
rect -67783 -40168 -67547 -39932
rect -67443 -40168 -67207 -39932
rect -67103 -40168 -66867 -39932
rect -66783 -40168 -66547 -39932
rect -66443 -40168 -66207 -39932
rect -66103 -40168 -65867 -39932
rect -65783 -40168 -65547 -39932
rect -65443 -40168 -65207 -39932
rect -65103 -40168 -64867 -39932
rect -64783 -40168 -64547 -39932
rect -64443 -40168 -64207 -39932
rect -64103 -40168 -63867 -39932
rect -63783 -40168 -63547 -39932
rect -63443 -40168 -63207 -39932
rect -63103 -40168 -62867 -39932
rect -62783 -40168 -62547 -39932
rect -62443 -40168 -62207 -39932
rect -62103 -40168 -61867 -39932
rect -61783 -40168 -61547 -39932
rect -61443 -40168 -61207 -39932
rect -61103 -40168 -60867 -39932
rect -60783 -40168 -60547 -39932
rect -60443 -40168 -60207 -39932
rect -60103 -40168 -59867 -39932
rect -59783 -40168 -59547 -39932
rect -59443 -40168 -59207 -39932
rect -59103 -40168 -58867 -39932
rect -58783 -40168 -58547 -39932
rect -58443 -40168 -58207 -39932
rect -58103 -40168 -57867 -39932
rect -57783 -40168 -57547 -39932
rect -57443 -40168 -57207 -39932
rect -57103 -40168 -56867 -39932
rect -56783 -40168 -56547 -39932
rect -56443 -40168 -56207 -39932
rect -56103 -40168 -55867 -39932
rect -55783 -40168 -55547 -39932
rect -55443 -40168 -55207 -39932
rect -55103 -40168 -54867 -39932
rect -54783 -40168 -54547 -39932
rect -54443 -40168 -54207 -39932
rect -54103 -40168 -53867 -39932
rect -53783 -40168 -53547 -39932
rect -53443 -40168 -53207 -39932
rect -53103 -40168 -52867 -39932
rect -52783 -40168 -52547 -39932
rect -52443 -40168 -52207 -39932
rect -52103 -40168 -51867 -39932
rect -51783 -40168 -51547 -39932
rect -51443 -40168 -51207 -39932
rect -51103 -40168 -50867 -39932
rect -50783 -40168 -50547 -39932
rect -50443 -40168 -50207 -39932
rect -50103 -40168 -49867 -39932
rect -49783 -40168 -49547 -39932
rect -49443 -40168 -49207 -39932
rect -49103 -40168 -48867 -39932
rect -74443 -40508 -74207 -40272
rect -74443 -40828 -74207 -40592
rect -73443 -40508 -73207 -40272
rect -73443 -40828 -73207 -40592
rect -72443 -40508 -72207 -40272
rect -72443 -40828 -72207 -40592
rect -71443 -40508 -71207 -40272
rect -71443 -40828 -71207 -40592
rect -70443 -40508 -70207 -40272
rect -70443 -40828 -70207 -40592
rect -69443 -40508 -69207 -40272
rect -69443 -40828 -69207 -40592
rect -68443 -40508 -68207 -40272
rect -68443 -40828 -68207 -40592
rect -67443 -40508 -67207 -40272
rect -67443 -40828 -67207 -40592
rect -66443 -40508 -66207 -40272
rect -66443 -40828 -66207 -40592
rect -65443 -40508 -65207 -40272
rect -65443 -40828 -65207 -40592
rect -64443 -40508 -64207 -40272
rect -64443 -40828 -64207 -40592
rect -63443 -40508 -63207 -40272
rect -63443 -40828 -63207 -40592
rect -62443 -40508 -62207 -40272
rect -62443 -40828 -62207 -40592
rect -61443 -40508 -61207 -40272
rect -61443 -40828 -61207 -40592
rect -60443 -40508 -60207 -40272
rect -60443 -40828 -60207 -40592
rect -59443 -40508 -59207 -40272
rect -59443 -40828 -59207 -40592
rect -58443 -40508 -58207 -40272
rect -58443 -40828 -58207 -40592
rect -57443 -40508 -57207 -40272
rect -57443 -40828 -57207 -40592
rect -56443 -40508 -56207 -40272
rect -56443 -40828 -56207 -40592
rect -55443 -40508 -55207 -40272
rect -55443 -40828 -55207 -40592
rect -54443 -40508 -54207 -40272
rect -54443 -40828 -54207 -40592
rect -53443 -40508 -53207 -40272
rect -53443 -40828 -53207 -40592
rect -52443 -40508 -52207 -40272
rect -52443 -40828 -52207 -40592
rect -51443 -40508 -51207 -40272
rect -51443 -40828 -51207 -40592
rect -50443 -40508 -50207 -40272
rect -50443 -40828 -50207 -40592
rect -49443 -40508 -49207 -40272
rect -49443 -40828 -49207 -40592
rect -74783 -41168 -74547 -40932
rect -74443 -41168 -74207 -40932
rect -74103 -41168 -73867 -40932
rect -73783 -41168 -73547 -40932
rect -73443 -41168 -73207 -40932
rect -73103 -41168 -72867 -40932
rect -72783 -41168 -72547 -40932
rect -72443 -41168 -72207 -40932
rect -72103 -41168 -71867 -40932
rect -71783 -41168 -71547 -40932
rect -71443 -41168 -71207 -40932
rect -71103 -41168 -70867 -40932
rect -70783 -41168 -70547 -40932
rect -70443 -41168 -70207 -40932
rect -70103 -41168 -69867 -40932
rect -69783 -41168 -69547 -40932
rect -69443 -41168 -69207 -40932
rect -69103 -41168 -68867 -40932
rect -68783 -41168 -68547 -40932
rect -68443 -41168 -68207 -40932
rect -68103 -41168 -67867 -40932
rect -67783 -41168 -67547 -40932
rect -67443 -41168 -67207 -40932
rect -67103 -41168 -66867 -40932
rect -66783 -41168 -66547 -40932
rect -66443 -41168 -66207 -40932
rect -66103 -41168 -65867 -40932
rect -65783 -41168 -65547 -40932
rect -65443 -41168 -65207 -40932
rect -65103 -41168 -64867 -40932
rect -64783 -41168 -64547 -40932
rect -64443 -41168 -64207 -40932
rect -64103 -41168 -63867 -40932
rect -63783 -41168 -63547 -40932
rect -63443 -41168 -63207 -40932
rect -63103 -41168 -62867 -40932
rect -62783 -41168 -62547 -40932
rect -62443 -41168 -62207 -40932
rect -62103 -41168 -61867 -40932
rect -61783 -41168 -61547 -40932
rect -61443 -41168 -61207 -40932
rect -61103 -41168 -60867 -40932
rect -60783 -41168 -60547 -40932
rect -60443 -41168 -60207 -40932
rect -60103 -41168 -59867 -40932
rect -59783 -41168 -59547 -40932
rect -59443 -41168 -59207 -40932
rect -59103 -41168 -58867 -40932
rect -58783 -41168 -58547 -40932
rect -58443 -41168 -58207 -40932
rect -58103 -41168 -57867 -40932
rect -57783 -41168 -57547 -40932
rect -57443 -41168 -57207 -40932
rect -57103 -41168 -56867 -40932
rect -56783 -41168 -56547 -40932
rect -56443 -41168 -56207 -40932
rect -56103 -41168 -55867 -40932
rect -55783 -41168 -55547 -40932
rect -55443 -41168 -55207 -40932
rect -55103 -41168 -54867 -40932
rect -54783 -41168 -54547 -40932
rect -54443 -41168 -54207 -40932
rect -54103 -41168 -53867 -40932
rect -53783 -41168 -53547 -40932
rect -53443 -41168 -53207 -40932
rect -53103 -41168 -52867 -40932
rect -52783 -41168 -52547 -40932
rect -52443 -41168 -52207 -40932
rect -52103 -41168 -51867 -40932
rect -51783 -41168 -51547 -40932
rect -51443 -41168 -51207 -40932
rect -51103 -41168 -50867 -40932
rect -50783 -41168 -50547 -40932
rect -50443 -41168 -50207 -40932
rect -50103 -41168 -49867 -40932
rect -49783 -41168 -49547 -40932
rect -49443 -41168 -49207 -40932
rect -49103 -41168 -48867 -40932
rect -74443 -41508 -74207 -41272
rect -74443 -41828 -74207 -41592
rect -73443 -41508 -73207 -41272
rect -73443 -41828 -73207 -41592
rect -72443 -41508 -72207 -41272
rect -72443 -41828 -72207 -41592
rect -71443 -41508 -71207 -41272
rect -71443 -41828 -71207 -41592
rect -70443 -41508 -70207 -41272
rect -70443 -41828 -70207 -41592
rect -69443 -41508 -69207 -41272
rect -69443 -41828 -69207 -41592
rect -68443 -41508 -68207 -41272
rect -68443 -41828 -68207 -41592
rect -67443 -41508 -67207 -41272
rect -67443 -41828 -67207 -41592
rect -66443 -41508 -66207 -41272
rect -66443 -41828 -66207 -41592
rect -65443 -41508 -65207 -41272
rect -65443 -41828 -65207 -41592
rect -64443 -41508 -64207 -41272
rect -64443 -41828 -64207 -41592
rect -63443 -41508 -63207 -41272
rect -63443 -41828 -63207 -41592
rect -62443 -41508 -62207 -41272
rect -62443 -41828 -62207 -41592
rect -61443 -41508 -61207 -41272
rect -61443 -41828 -61207 -41592
rect -60443 -41508 -60207 -41272
rect -60443 -41828 -60207 -41592
rect -59443 -41508 -59207 -41272
rect -59443 -41828 -59207 -41592
rect -58443 -41508 -58207 -41272
rect -58443 -41828 -58207 -41592
rect -57443 -41508 -57207 -41272
rect -57443 -41828 -57207 -41592
rect -56443 -41508 -56207 -41272
rect -56443 -41828 -56207 -41592
rect -55443 -41508 -55207 -41272
rect -55443 -41828 -55207 -41592
rect -54443 -41508 -54207 -41272
rect -54443 -41828 -54207 -41592
rect -53443 -41508 -53207 -41272
rect -53443 -41828 -53207 -41592
rect -52443 -41508 -52207 -41272
rect -52443 -41828 -52207 -41592
rect -51443 -41508 -51207 -41272
rect -51443 -41828 -51207 -41592
rect -50443 -41508 -50207 -41272
rect -50443 -41828 -50207 -41592
rect -49443 -41508 -49207 -41272
rect -49443 -41828 -49207 -41592
rect -74783 -42168 -74547 -41932
rect -74443 -42168 -74207 -41932
rect -74103 -42168 -73867 -41932
rect -73783 -42168 -73547 -41932
rect -73443 -42168 -73207 -41932
rect -73103 -42168 -72867 -41932
rect -72783 -42168 -72547 -41932
rect -72443 -42168 -72207 -41932
rect -72103 -42168 -71867 -41932
rect -71783 -42168 -71547 -41932
rect -71443 -42168 -71207 -41932
rect -71103 -42168 -70867 -41932
rect -70783 -42168 -70547 -41932
rect -70443 -42168 -70207 -41932
rect -70103 -42168 -69867 -41932
rect -69783 -42168 -69547 -41932
rect -69443 -42168 -69207 -41932
rect -69103 -42168 -68867 -41932
rect -68783 -42168 -68547 -41932
rect -68443 -42168 -68207 -41932
rect -68103 -42168 -67867 -41932
rect -67783 -42168 -67547 -41932
rect -67443 -42168 -67207 -41932
rect -67103 -42168 -66867 -41932
rect -66783 -42168 -66547 -41932
rect -66443 -42168 -66207 -41932
rect -66103 -42168 -65867 -41932
rect -65783 -42168 -65547 -41932
rect -65443 -42168 -65207 -41932
rect -65103 -42168 -64867 -41932
rect -64783 -42168 -64547 -41932
rect -64443 -42168 -64207 -41932
rect -64103 -42168 -63867 -41932
rect -63783 -42168 -63547 -41932
rect -63443 -42168 -63207 -41932
rect -63103 -42168 -62867 -41932
rect -62783 -42168 -62547 -41932
rect -62443 -42168 -62207 -41932
rect -62103 -42168 -61867 -41932
rect -61783 -42168 -61547 -41932
rect -61443 -42168 -61207 -41932
rect -61103 -42168 -60867 -41932
rect -60783 -42168 -60547 -41932
rect -60443 -42168 -60207 -41932
rect -60103 -42168 -59867 -41932
rect -59783 -42168 -59547 -41932
rect -59443 -42168 -59207 -41932
rect -59103 -42168 -58867 -41932
rect -58783 -42168 -58547 -41932
rect -58443 -42168 -58207 -41932
rect -58103 -42168 -57867 -41932
rect -57783 -42168 -57547 -41932
rect -57443 -42168 -57207 -41932
rect -57103 -42168 -56867 -41932
rect -56783 -42168 -56547 -41932
rect -56443 -42168 -56207 -41932
rect -56103 -42168 -55867 -41932
rect -55783 -42168 -55547 -41932
rect -55443 -42168 -55207 -41932
rect -55103 -42168 -54867 -41932
rect -54783 -42168 -54547 -41932
rect -54443 -42168 -54207 -41932
rect -54103 -42168 -53867 -41932
rect -53783 -42168 -53547 -41932
rect -53443 -42168 -53207 -41932
rect -53103 -42168 -52867 -41932
rect -52783 -42168 -52547 -41932
rect -52443 -42168 -52207 -41932
rect -52103 -42168 -51867 -41932
rect -51783 -42168 -51547 -41932
rect -51443 -42168 -51207 -41932
rect -51103 -42168 -50867 -41932
rect -50783 -42168 -50547 -41932
rect -50443 -42168 -50207 -41932
rect -50103 -42168 -49867 -41932
rect -49783 -42168 -49547 -41932
rect -49443 -42168 -49207 -41932
rect -49103 -42168 -48867 -41932
rect -74443 -42508 -74207 -42272
rect -74443 -42828 -74207 -42592
rect -73443 -42508 -73207 -42272
rect -73443 -42828 -73207 -42592
rect -72443 -42508 -72207 -42272
rect -72443 -42828 -72207 -42592
rect -71443 -42508 -71207 -42272
rect -71443 -42828 -71207 -42592
rect -70443 -42508 -70207 -42272
rect -70443 -42828 -70207 -42592
rect -69443 -42508 -69207 -42272
rect -69443 -42828 -69207 -42592
rect -68443 -42508 -68207 -42272
rect -68443 -42828 -68207 -42592
rect -67443 -42508 -67207 -42272
rect -67443 -42828 -67207 -42592
rect -66443 -42508 -66207 -42272
rect -66443 -42828 -66207 -42592
rect -65443 -42508 -65207 -42272
rect -65443 -42828 -65207 -42592
rect -64443 -42508 -64207 -42272
rect -64443 -42828 -64207 -42592
rect -63443 -42508 -63207 -42272
rect -63443 -42828 -63207 -42592
rect -62443 -42508 -62207 -42272
rect -62443 -42828 -62207 -42592
rect -61443 -42508 -61207 -42272
rect -61443 -42828 -61207 -42592
rect -60443 -42508 -60207 -42272
rect -60443 -42828 -60207 -42592
rect -59443 -42508 -59207 -42272
rect -59443 -42828 -59207 -42592
rect -58443 -42508 -58207 -42272
rect -58443 -42828 -58207 -42592
rect -57443 -42508 -57207 -42272
rect -57443 -42828 -57207 -42592
rect -56443 -42508 -56207 -42272
rect -56443 -42828 -56207 -42592
rect -55443 -42508 -55207 -42272
rect -55443 -42828 -55207 -42592
rect -54443 -42508 -54207 -42272
rect -54443 -42828 -54207 -42592
rect -53443 -42508 -53207 -42272
rect -53443 -42828 -53207 -42592
rect -52443 -42508 -52207 -42272
rect -52443 -42828 -52207 -42592
rect -51443 -42508 -51207 -42272
rect -51443 -42828 -51207 -42592
rect -50443 -42508 -50207 -42272
rect -50443 -42828 -50207 -42592
rect -49443 -42508 -49207 -42272
rect -49443 -42828 -49207 -42592
rect -74783 -43168 -74547 -42932
rect -74443 -43168 -74207 -42932
rect -74103 -43168 -73867 -42932
rect -73783 -43168 -73547 -42932
rect -73443 -43168 -73207 -42932
rect -73103 -43168 -72867 -42932
rect -72783 -43168 -72547 -42932
rect -72443 -43168 -72207 -42932
rect -72103 -43168 -71867 -42932
rect -71783 -43168 -71547 -42932
rect -71443 -43168 -71207 -42932
rect -71103 -43168 -70867 -42932
rect -70783 -43168 -70547 -42932
rect -70443 -43168 -70207 -42932
rect -70103 -43168 -69867 -42932
rect -69783 -43168 -69547 -42932
rect -69443 -43168 -69207 -42932
rect -69103 -43168 -68867 -42932
rect -68783 -43168 -68547 -42932
rect -68443 -43168 -68207 -42932
rect -68103 -43168 -67867 -42932
rect -67783 -43168 -67547 -42932
rect -67443 -43168 -67207 -42932
rect -67103 -43168 -66867 -42932
rect -66783 -43168 -66547 -42932
rect -66443 -43168 -66207 -42932
rect -66103 -43168 -65867 -42932
rect -65783 -43168 -65547 -42932
rect -65443 -43168 -65207 -42932
rect -65103 -43168 -64867 -42932
rect -64783 -43168 -64547 -42932
rect -64443 -43168 -64207 -42932
rect -64103 -43168 -63867 -42932
rect -63783 -43168 -63547 -42932
rect -63443 -43168 -63207 -42932
rect -63103 -43168 -62867 -42932
rect -62783 -43168 -62547 -42932
rect -62443 -43168 -62207 -42932
rect -62103 -43168 -61867 -42932
rect -61783 -43168 -61547 -42932
rect -61443 -43168 -61207 -42932
rect -61103 -43168 -60867 -42932
rect -60783 -43168 -60547 -42932
rect -60443 -43168 -60207 -42932
rect -60103 -43168 -59867 -42932
rect -59783 -43168 -59547 -42932
rect -59443 -43168 -59207 -42932
rect -59103 -43168 -58867 -42932
rect -58783 -43168 -58547 -42932
rect -58443 -43168 -58207 -42932
rect -58103 -43168 -57867 -42932
rect -57783 -43168 -57547 -42932
rect -57443 -43168 -57207 -42932
rect -57103 -43168 -56867 -42932
rect -56783 -43168 -56547 -42932
rect -56443 -43168 -56207 -42932
rect -56103 -43168 -55867 -42932
rect -55783 -43168 -55547 -42932
rect -55443 -43168 -55207 -42932
rect -55103 -43168 -54867 -42932
rect -54783 -43168 -54547 -42932
rect -54443 -43168 -54207 -42932
rect -54103 -43168 -53867 -42932
rect -53783 -43168 -53547 -42932
rect -53443 -43168 -53207 -42932
rect -53103 -43168 -52867 -42932
rect -52783 -43168 -52547 -42932
rect -52443 -43168 -52207 -42932
rect -52103 -43168 -51867 -42932
rect -51783 -43168 -51547 -42932
rect -51443 -43168 -51207 -42932
rect -51103 -43168 -50867 -42932
rect -50783 -43168 -50547 -42932
rect -50443 -43168 -50207 -42932
rect -50103 -43168 -49867 -42932
rect -49783 -43168 -49547 -42932
rect -49443 -43168 -49207 -42932
rect -49103 -43168 -48867 -42932
rect -74443 -43508 -74207 -43272
rect -74443 -43828 -74207 -43592
rect -73443 -43508 -73207 -43272
rect -73443 -43828 -73207 -43592
rect -72443 -43508 -72207 -43272
rect -72443 -43828 -72207 -43592
rect -71443 -43508 -71207 -43272
rect -71443 -43828 -71207 -43592
rect -70443 -43508 -70207 -43272
rect -70443 -43828 -70207 -43592
rect -69443 -43508 -69207 -43272
rect -69443 -43828 -69207 -43592
rect -68443 -43508 -68207 -43272
rect -68443 -43828 -68207 -43592
rect -67443 -43508 -67207 -43272
rect -67443 -43828 -67207 -43592
rect -66443 -43508 -66207 -43272
rect -66443 -43828 -66207 -43592
rect -65443 -43508 -65207 -43272
rect -65443 -43828 -65207 -43592
rect -64443 -43508 -64207 -43272
rect -64443 -43828 -64207 -43592
rect -63443 -43508 -63207 -43272
rect -63443 -43828 -63207 -43592
rect -62443 -43508 -62207 -43272
rect -62443 -43828 -62207 -43592
rect -61443 -43508 -61207 -43272
rect -61443 -43828 -61207 -43592
rect -60443 -43508 -60207 -43272
rect -60443 -43828 -60207 -43592
rect -59443 -43508 -59207 -43272
rect -59443 -43828 -59207 -43592
rect -58443 -43508 -58207 -43272
rect -58443 -43828 -58207 -43592
rect -57443 -43508 -57207 -43272
rect -57443 -43828 -57207 -43592
rect -56443 -43508 -56207 -43272
rect -56443 -43828 -56207 -43592
rect -55443 -43508 -55207 -43272
rect -55443 -43828 -55207 -43592
rect -54443 -43508 -54207 -43272
rect -54443 -43828 -54207 -43592
rect -53443 -43508 -53207 -43272
rect -53443 -43828 -53207 -43592
rect -52443 -43508 -52207 -43272
rect -52443 -43828 -52207 -43592
rect -51443 -43508 -51207 -43272
rect -51443 -43828 -51207 -43592
rect -50443 -43508 -50207 -43272
rect -50443 -43828 -50207 -43592
rect -49443 -43508 -49207 -43272
rect -49443 -43828 -49207 -43592
rect -74783 -44168 -74547 -43932
rect -74443 -44168 -74207 -43932
rect -74103 -44168 -73867 -43932
rect -73783 -44168 -73547 -43932
rect -73443 -44168 -73207 -43932
rect -73103 -44168 -72867 -43932
rect -72783 -44168 -72547 -43932
rect -72443 -44168 -72207 -43932
rect -72103 -44168 -71867 -43932
rect -71783 -44168 -71547 -43932
rect -71443 -44168 -71207 -43932
rect -71103 -44168 -70867 -43932
rect -70783 -44168 -70547 -43932
rect -70443 -44168 -70207 -43932
rect -70103 -44168 -69867 -43932
rect -69783 -44168 -69547 -43932
rect -69443 -44168 -69207 -43932
rect -69103 -44168 -68867 -43932
rect -68783 -44168 -68547 -43932
rect -68443 -44168 -68207 -43932
rect -68103 -44168 -67867 -43932
rect -67783 -44168 -67547 -43932
rect -67443 -44168 -67207 -43932
rect -67103 -44168 -66867 -43932
rect -66783 -44168 -66547 -43932
rect -66443 -44168 -66207 -43932
rect -66103 -44168 -65867 -43932
rect -65783 -44168 -65547 -43932
rect -65443 -44168 -65207 -43932
rect -65103 -44168 -64867 -43932
rect -64783 -44168 -64547 -43932
rect -64443 -44168 -64207 -43932
rect -64103 -44168 -63867 -43932
rect -63783 -44168 -63547 -43932
rect -63443 -44168 -63207 -43932
rect -63103 -44168 -62867 -43932
rect -62783 -44168 -62547 -43932
rect -62443 -44168 -62207 -43932
rect -62103 -44168 -61867 -43932
rect -61783 -44168 -61547 -43932
rect -61443 -44168 -61207 -43932
rect -61103 -44168 -60867 -43932
rect -60783 -44168 -60547 -43932
rect -60443 -44168 -60207 -43932
rect -60103 -44168 -59867 -43932
rect -59783 -44168 -59547 -43932
rect -59443 -44168 -59207 -43932
rect -59103 -44168 -58867 -43932
rect -58783 -44168 -58547 -43932
rect -58443 -44168 -58207 -43932
rect -58103 -44168 -57867 -43932
rect -57783 -44168 -57547 -43932
rect -57443 -44168 -57207 -43932
rect -57103 -44168 -56867 -43932
rect -56783 -44168 -56547 -43932
rect -56443 -44168 -56207 -43932
rect -56103 -44168 -55867 -43932
rect -55783 -44168 -55547 -43932
rect -55443 -44168 -55207 -43932
rect -55103 -44168 -54867 -43932
rect -54783 -44168 -54547 -43932
rect -54443 -44168 -54207 -43932
rect -54103 -44168 -53867 -43932
rect -53783 -44168 -53547 -43932
rect -53443 -44168 -53207 -43932
rect -53103 -44168 -52867 -43932
rect -52783 -44168 -52547 -43932
rect -52443 -44168 -52207 -43932
rect -52103 -44168 -51867 -43932
rect -51783 -44168 -51547 -43932
rect -51443 -44168 -51207 -43932
rect -51103 -44168 -50867 -43932
rect -50783 -44168 -50547 -43932
rect -50443 -44168 -50207 -43932
rect -50103 -44168 -49867 -43932
rect -49783 -44168 -49547 -43932
rect -49443 -44168 -49207 -43932
rect -49103 -44168 -48867 -43932
rect -74443 -44508 -74207 -44272
rect -74443 -44828 -74207 -44592
rect -73443 -44508 -73207 -44272
rect -73443 -44828 -73207 -44592
rect -72443 -44508 -72207 -44272
rect -72443 -44828 -72207 -44592
rect -71443 -44508 -71207 -44272
rect -71443 -44828 -71207 -44592
rect -70443 -44508 -70207 -44272
rect -70443 -44828 -70207 -44592
rect -69443 -44508 -69207 -44272
rect -69443 -44828 -69207 -44592
rect -68443 -44508 -68207 -44272
rect -68443 -44828 -68207 -44592
rect -67443 -44508 -67207 -44272
rect -67443 -44828 -67207 -44592
rect -66443 -44508 -66207 -44272
rect -66443 -44828 -66207 -44592
rect -65443 -44508 -65207 -44272
rect -65443 -44828 -65207 -44592
rect -64443 -44508 -64207 -44272
rect -64443 -44828 -64207 -44592
rect -63443 -44508 -63207 -44272
rect -63443 -44828 -63207 -44592
rect -62443 -44508 -62207 -44272
rect -62443 -44828 -62207 -44592
rect -61443 -44508 -61207 -44272
rect -61443 -44828 -61207 -44592
rect -60443 -44508 -60207 -44272
rect -60443 -44828 -60207 -44592
rect -59443 -44508 -59207 -44272
rect -59443 -44828 -59207 -44592
rect -58443 -44508 -58207 -44272
rect -58443 -44828 -58207 -44592
rect -57443 -44508 -57207 -44272
rect -57443 -44828 -57207 -44592
rect -56443 -44508 -56207 -44272
rect -56443 -44828 -56207 -44592
rect -55443 -44508 -55207 -44272
rect -55443 -44828 -55207 -44592
rect -54443 -44508 -54207 -44272
rect -54443 -44828 -54207 -44592
rect -53443 -44508 -53207 -44272
rect -53443 -44828 -53207 -44592
rect -52443 -44508 -52207 -44272
rect -52443 -44828 -52207 -44592
rect -51443 -44508 -51207 -44272
rect -51443 -44828 -51207 -44592
rect -50443 -44508 -50207 -44272
rect -50443 -44828 -50207 -44592
rect -49443 -44508 -49207 -44272
rect -49443 -44828 -49207 -44592
rect -46198 -44428 -36362 -32672
rect -4198 -44428 5638 -32672
rect 8657 -32508 8893 -32272
rect 8657 -32828 8893 -32592
rect 9657 -32508 9893 -32272
rect 9657 -32828 9893 -32592
rect 10657 -32508 10893 -32272
rect 10657 -32828 10893 -32592
rect 11657 -32508 11893 -32272
rect 11657 -32828 11893 -32592
rect 12657 -32508 12893 -32272
rect 12657 -32828 12893 -32592
rect 13657 -32508 13893 -32272
rect 13657 -32828 13893 -32592
rect 14657 -32508 14893 -32272
rect 14657 -32828 14893 -32592
rect 15657 -32508 15893 -32272
rect 15657 -32828 15893 -32592
rect 16657 -32508 16893 -32272
rect 16657 -32828 16893 -32592
rect 17657 -32508 17893 -32272
rect 17657 -32828 17893 -32592
rect 18657 -32508 18893 -32272
rect 18657 -32828 18893 -32592
rect 19657 -32508 19893 -32272
rect 19657 -32828 19893 -32592
rect 20657 -32508 20893 -32272
rect 20657 -32828 20893 -32592
rect 21657 -32508 21893 -32272
rect 21657 -32828 21893 -32592
rect 22657 -32508 22893 -32272
rect 22657 -32828 22893 -32592
rect 23657 -32508 23893 -32272
rect 23657 -32828 23893 -32592
rect 24657 -32508 24893 -32272
rect 24657 -32828 24893 -32592
rect 25657 -32508 25893 -32272
rect 25657 -32828 25893 -32592
rect 26657 -32508 26893 -32272
rect 26657 -32828 26893 -32592
rect 27657 -32508 27893 -32272
rect 27657 -32828 27893 -32592
rect 28657 -32508 28893 -32272
rect 28657 -32828 28893 -32592
rect 29657 -32508 29893 -32272
rect 29657 -32828 29893 -32592
rect 30657 -32508 30893 -32272
rect 30657 -32828 30893 -32592
rect 31657 -32508 31893 -32272
rect 31657 -32828 31893 -32592
rect 32657 -32508 32893 -32272
rect 32657 -32828 32893 -32592
rect 33657 -32508 33893 -32272
rect 33657 -32828 33893 -32592
rect 8317 -33168 8553 -32932
rect 8657 -33168 8893 -32932
rect 8997 -33168 9233 -32932
rect 9317 -33168 9553 -32932
rect 9657 -33168 9893 -32932
rect 9997 -33168 10233 -32932
rect 10317 -33168 10553 -32932
rect 10657 -33168 10893 -32932
rect 10997 -33168 11233 -32932
rect 11317 -33168 11553 -32932
rect 11657 -33168 11893 -32932
rect 11997 -33168 12233 -32932
rect 12317 -33168 12553 -32932
rect 12657 -33168 12893 -32932
rect 12997 -33168 13233 -32932
rect 13317 -33168 13553 -32932
rect 13657 -33168 13893 -32932
rect 13997 -33168 14233 -32932
rect 14317 -33168 14553 -32932
rect 14657 -33168 14893 -32932
rect 14997 -33168 15233 -32932
rect 15317 -33168 15553 -32932
rect 15657 -33168 15893 -32932
rect 15997 -33168 16233 -32932
rect 16317 -33168 16553 -32932
rect 16657 -33168 16893 -32932
rect 16997 -33168 17233 -32932
rect 17317 -33168 17553 -32932
rect 17657 -33168 17893 -32932
rect 17997 -33168 18233 -32932
rect 18317 -33168 18553 -32932
rect 18657 -33168 18893 -32932
rect 18997 -33168 19233 -32932
rect 19317 -33168 19553 -32932
rect 19657 -33168 19893 -32932
rect 19997 -33168 20233 -32932
rect 20317 -33168 20553 -32932
rect 20657 -33168 20893 -32932
rect 20997 -33168 21233 -32932
rect 21317 -33168 21553 -32932
rect 21657 -33168 21893 -32932
rect 21997 -33168 22233 -32932
rect 22317 -33168 22553 -32932
rect 22657 -33168 22893 -32932
rect 22997 -33168 23233 -32932
rect 23317 -33168 23553 -32932
rect 23657 -33168 23893 -32932
rect 23997 -33168 24233 -32932
rect 24317 -33168 24553 -32932
rect 24657 -33168 24893 -32932
rect 24997 -33168 25233 -32932
rect 25317 -33168 25553 -32932
rect 25657 -33168 25893 -32932
rect 25997 -33168 26233 -32932
rect 26317 -33168 26553 -32932
rect 26657 -33168 26893 -32932
rect 26997 -33168 27233 -32932
rect 27317 -33168 27553 -32932
rect 27657 -33168 27893 -32932
rect 27997 -33168 28233 -32932
rect 28317 -33168 28553 -32932
rect 28657 -33168 28893 -32932
rect 28997 -33168 29233 -32932
rect 29317 -33168 29553 -32932
rect 29657 -33168 29893 -32932
rect 29997 -33168 30233 -32932
rect 30317 -33168 30553 -32932
rect 30657 -33168 30893 -32932
rect 30997 -33168 31233 -32932
rect 31317 -33168 31553 -32932
rect 31657 -33168 31893 -32932
rect 31997 -33168 32233 -32932
rect 32317 -33168 32553 -32932
rect 32657 -33168 32893 -32932
rect 32997 -33168 33233 -32932
rect 33317 -33168 33553 -32932
rect 33657 -33168 33893 -32932
rect 33997 -33168 34233 -32932
rect 8657 -33508 8893 -33272
rect 8657 -33828 8893 -33592
rect 9657 -33508 9893 -33272
rect 9657 -33828 9893 -33592
rect 10657 -33508 10893 -33272
rect 10657 -33828 10893 -33592
rect 11657 -33508 11893 -33272
rect 11657 -33828 11893 -33592
rect 12657 -33508 12893 -33272
rect 12657 -33828 12893 -33592
rect 13657 -33508 13893 -33272
rect 13657 -33828 13893 -33592
rect 14657 -33508 14893 -33272
rect 14657 -33828 14893 -33592
rect 15657 -33508 15893 -33272
rect 15657 -33828 15893 -33592
rect 16657 -33508 16893 -33272
rect 16657 -33828 16893 -33592
rect 17657 -33508 17893 -33272
rect 17657 -33828 17893 -33592
rect 18657 -33508 18893 -33272
rect 18657 -33828 18893 -33592
rect 19657 -33508 19893 -33272
rect 19657 -33828 19893 -33592
rect 20657 -33508 20893 -33272
rect 20657 -33828 20893 -33592
rect 21657 -33508 21893 -33272
rect 21657 -33828 21893 -33592
rect 22657 -33508 22893 -33272
rect 22657 -33828 22893 -33592
rect 23657 -33508 23893 -33272
rect 23657 -33828 23893 -33592
rect 24657 -33508 24893 -33272
rect 24657 -33828 24893 -33592
rect 25657 -33508 25893 -33272
rect 25657 -33828 25893 -33592
rect 26657 -33508 26893 -33272
rect 26657 -33828 26893 -33592
rect 27657 -33508 27893 -33272
rect 27657 -33828 27893 -33592
rect 28657 -33508 28893 -33272
rect 28657 -33828 28893 -33592
rect 29657 -33508 29893 -33272
rect 29657 -33828 29893 -33592
rect 30657 -33508 30893 -33272
rect 30657 -33828 30893 -33592
rect 31657 -33508 31893 -33272
rect 31657 -33828 31893 -33592
rect 32657 -33508 32893 -33272
rect 32657 -33828 32893 -33592
rect 33657 -33508 33893 -33272
rect 33657 -33828 33893 -33592
rect 8317 -34168 8553 -33932
rect 8657 -34168 8893 -33932
rect 8997 -34168 9233 -33932
rect 9317 -34168 9553 -33932
rect 9657 -34168 9893 -33932
rect 9997 -34168 10233 -33932
rect 10317 -34168 10553 -33932
rect 10657 -34168 10893 -33932
rect 10997 -34168 11233 -33932
rect 11317 -34168 11553 -33932
rect 11657 -34168 11893 -33932
rect 11997 -34168 12233 -33932
rect 12317 -34168 12553 -33932
rect 12657 -34168 12893 -33932
rect 12997 -34168 13233 -33932
rect 13317 -34168 13553 -33932
rect 13657 -34168 13893 -33932
rect 13997 -34168 14233 -33932
rect 14317 -34168 14553 -33932
rect 14657 -34168 14893 -33932
rect 14997 -34168 15233 -33932
rect 15317 -34168 15553 -33932
rect 15657 -34168 15893 -33932
rect 15997 -34168 16233 -33932
rect 16317 -34168 16553 -33932
rect 16657 -34168 16893 -33932
rect 16997 -34168 17233 -33932
rect 17317 -34168 17553 -33932
rect 17657 -34168 17893 -33932
rect 17997 -34168 18233 -33932
rect 18317 -34168 18553 -33932
rect 18657 -34168 18893 -33932
rect 18997 -34168 19233 -33932
rect 19317 -34168 19553 -33932
rect 19657 -34168 19893 -33932
rect 19997 -34168 20233 -33932
rect 20317 -34168 20553 -33932
rect 20657 -34168 20893 -33932
rect 20997 -34168 21233 -33932
rect 21317 -34168 21553 -33932
rect 21657 -34168 21893 -33932
rect 21997 -34168 22233 -33932
rect 22317 -34168 22553 -33932
rect 22657 -34168 22893 -33932
rect 22997 -34168 23233 -33932
rect 23317 -34168 23553 -33932
rect 23657 -34168 23893 -33932
rect 23997 -34168 24233 -33932
rect 24317 -34168 24553 -33932
rect 24657 -34168 24893 -33932
rect 24997 -34168 25233 -33932
rect 25317 -34168 25553 -33932
rect 25657 -34168 25893 -33932
rect 25997 -34168 26233 -33932
rect 26317 -34168 26553 -33932
rect 26657 -34168 26893 -33932
rect 26997 -34168 27233 -33932
rect 27317 -34168 27553 -33932
rect 27657 -34168 27893 -33932
rect 27997 -34168 28233 -33932
rect 28317 -34168 28553 -33932
rect 28657 -34168 28893 -33932
rect 28997 -34168 29233 -33932
rect 29317 -34168 29553 -33932
rect 29657 -34168 29893 -33932
rect 29997 -34168 30233 -33932
rect 30317 -34168 30553 -33932
rect 30657 -34168 30893 -33932
rect 30997 -34168 31233 -33932
rect 31317 -34168 31553 -33932
rect 31657 -34168 31893 -33932
rect 31997 -34168 32233 -33932
rect 32317 -34168 32553 -33932
rect 32657 -34168 32893 -33932
rect 32997 -34168 33233 -33932
rect 33317 -34168 33553 -33932
rect 33657 -34168 33893 -33932
rect 33997 -34168 34233 -33932
rect 8657 -34508 8893 -34272
rect 8657 -34828 8893 -34592
rect 9657 -34508 9893 -34272
rect 9657 -34828 9893 -34592
rect 10657 -34508 10893 -34272
rect 10657 -34828 10893 -34592
rect 11657 -34508 11893 -34272
rect 11657 -34828 11893 -34592
rect 12657 -34508 12893 -34272
rect 12657 -34828 12893 -34592
rect 13657 -34508 13893 -34272
rect 13657 -34828 13893 -34592
rect 14657 -34508 14893 -34272
rect 14657 -34828 14893 -34592
rect 15657 -34508 15893 -34272
rect 15657 -34828 15893 -34592
rect 16657 -34508 16893 -34272
rect 16657 -34828 16893 -34592
rect 17657 -34508 17893 -34272
rect 17657 -34828 17893 -34592
rect 18657 -34508 18893 -34272
rect 18657 -34828 18893 -34592
rect 19657 -34508 19893 -34272
rect 19657 -34828 19893 -34592
rect 20657 -34508 20893 -34272
rect 20657 -34828 20893 -34592
rect 21657 -34508 21893 -34272
rect 21657 -34828 21893 -34592
rect 22657 -34508 22893 -34272
rect 22657 -34828 22893 -34592
rect 23657 -34508 23893 -34272
rect 23657 -34828 23893 -34592
rect 24657 -34508 24893 -34272
rect 24657 -34828 24893 -34592
rect 25657 -34508 25893 -34272
rect 25657 -34828 25893 -34592
rect 26657 -34508 26893 -34272
rect 26657 -34828 26893 -34592
rect 27657 -34508 27893 -34272
rect 27657 -34828 27893 -34592
rect 28657 -34508 28893 -34272
rect 28657 -34828 28893 -34592
rect 29657 -34508 29893 -34272
rect 29657 -34828 29893 -34592
rect 30657 -34508 30893 -34272
rect 30657 -34828 30893 -34592
rect 31657 -34508 31893 -34272
rect 31657 -34828 31893 -34592
rect 32657 -34508 32893 -34272
rect 32657 -34828 32893 -34592
rect 33657 -34508 33893 -34272
rect 33657 -34828 33893 -34592
rect 8317 -35168 8553 -34932
rect 8657 -35168 8893 -34932
rect 8997 -35168 9233 -34932
rect 9317 -35168 9553 -34932
rect 9657 -35168 9893 -34932
rect 9997 -35168 10233 -34932
rect 10317 -35168 10553 -34932
rect 10657 -35168 10893 -34932
rect 10997 -35168 11233 -34932
rect 11317 -35168 11553 -34932
rect 11657 -35168 11893 -34932
rect 11997 -35168 12233 -34932
rect 12317 -35168 12553 -34932
rect 12657 -35168 12893 -34932
rect 12997 -35168 13233 -34932
rect 13317 -35168 13553 -34932
rect 13657 -35168 13893 -34932
rect 13997 -35168 14233 -34932
rect 14317 -35168 14553 -34932
rect 14657 -35168 14893 -34932
rect 14997 -35168 15233 -34932
rect 15317 -35168 15553 -34932
rect 15657 -35168 15893 -34932
rect 15997 -35168 16233 -34932
rect 16317 -35168 16553 -34932
rect 16657 -35168 16893 -34932
rect 16997 -35168 17233 -34932
rect 17317 -35168 17553 -34932
rect 17657 -35168 17893 -34932
rect 17997 -35168 18233 -34932
rect 18317 -35168 18553 -34932
rect 18657 -35168 18893 -34932
rect 18997 -35168 19233 -34932
rect 19317 -35168 19553 -34932
rect 19657 -35168 19893 -34932
rect 19997 -35168 20233 -34932
rect 20317 -35168 20553 -34932
rect 20657 -35168 20893 -34932
rect 20997 -35168 21233 -34932
rect 21317 -35168 21553 -34932
rect 21657 -35168 21893 -34932
rect 21997 -35168 22233 -34932
rect 22317 -35168 22553 -34932
rect 22657 -35168 22893 -34932
rect 22997 -35168 23233 -34932
rect 23317 -35168 23553 -34932
rect 23657 -35168 23893 -34932
rect 23997 -35168 24233 -34932
rect 24317 -35168 24553 -34932
rect 24657 -35168 24893 -34932
rect 24997 -35168 25233 -34932
rect 25317 -35168 25553 -34932
rect 25657 -35168 25893 -34932
rect 25997 -35168 26233 -34932
rect 26317 -35168 26553 -34932
rect 26657 -35168 26893 -34932
rect 26997 -35168 27233 -34932
rect 27317 -35168 27553 -34932
rect 27657 -35168 27893 -34932
rect 27997 -35168 28233 -34932
rect 28317 -35168 28553 -34932
rect 28657 -35168 28893 -34932
rect 28997 -35168 29233 -34932
rect 29317 -35168 29553 -34932
rect 29657 -35168 29893 -34932
rect 29997 -35168 30233 -34932
rect 30317 -35168 30553 -34932
rect 30657 -35168 30893 -34932
rect 30997 -35168 31233 -34932
rect 31317 -35168 31553 -34932
rect 31657 -35168 31893 -34932
rect 31997 -35168 32233 -34932
rect 32317 -35168 32553 -34932
rect 32657 -35168 32893 -34932
rect 32997 -35168 33233 -34932
rect 33317 -35168 33553 -34932
rect 33657 -35168 33893 -34932
rect 33997 -35168 34233 -34932
rect 8657 -35508 8893 -35272
rect 8657 -35828 8893 -35592
rect 9657 -35508 9893 -35272
rect 9657 -35828 9893 -35592
rect 10657 -35508 10893 -35272
rect 10657 -35828 10893 -35592
rect 11657 -35508 11893 -35272
rect 11657 -35828 11893 -35592
rect 12657 -35508 12893 -35272
rect 12657 -35828 12893 -35592
rect 13657 -35508 13893 -35272
rect 13657 -35828 13893 -35592
rect 14657 -35508 14893 -35272
rect 14657 -35828 14893 -35592
rect 15657 -35508 15893 -35272
rect 15657 -35828 15893 -35592
rect 16657 -35508 16893 -35272
rect 16657 -35828 16893 -35592
rect 17657 -35508 17893 -35272
rect 17657 -35828 17893 -35592
rect 18657 -35508 18893 -35272
rect 18657 -35828 18893 -35592
rect 19657 -35508 19893 -35272
rect 19657 -35828 19893 -35592
rect 20657 -35508 20893 -35272
rect 20657 -35828 20893 -35592
rect 21657 -35508 21893 -35272
rect 21657 -35828 21893 -35592
rect 22657 -35508 22893 -35272
rect 22657 -35828 22893 -35592
rect 23657 -35508 23893 -35272
rect 23657 -35828 23893 -35592
rect 24657 -35508 24893 -35272
rect 24657 -35828 24893 -35592
rect 25657 -35508 25893 -35272
rect 25657 -35828 25893 -35592
rect 26657 -35508 26893 -35272
rect 26657 -35828 26893 -35592
rect 27657 -35508 27893 -35272
rect 27657 -35828 27893 -35592
rect 28657 -35508 28893 -35272
rect 28657 -35828 28893 -35592
rect 29657 -35508 29893 -35272
rect 29657 -35828 29893 -35592
rect 30657 -35508 30893 -35272
rect 30657 -35828 30893 -35592
rect 31657 -35508 31893 -35272
rect 31657 -35828 31893 -35592
rect 32657 -35508 32893 -35272
rect 32657 -35828 32893 -35592
rect 33657 -35508 33893 -35272
rect 33657 -35828 33893 -35592
rect 8317 -36168 8553 -35932
rect 8657 -36168 8893 -35932
rect 8997 -36168 9233 -35932
rect 9317 -36168 9553 -35932
rect 9657 -36168 9893 -35932
rect 9997 -36168 10233 -35932
rect 10317 -36168 10553 -35932
rect 10657 -36168 10893 -35932
rect 10997 -36168 11233 -35932
rect 11317 -36168 11553 -35932
rect 11657 -36168 11893 -35932
rect 11997 -36168 12233 -35932
rect 12317 -36168 12553 -35932
rect 12657 -36168 12893 -35932
rect 12997 -36168 13233 -35932
rect 13317 -36168 13553 -35932
rect 13657 -36168 13893 -35932
rect 13997 -36168 14233 -35932
rect 14317 -36168 14553 -35932
rect 14657 -36168 14893 -35932
rect 14997 -36168 15233 -35932
rect 15317 -36168 15553 -35932
rect 15657 -36168 15893 -35932
rect 15997 -36168 16233 -35932
rect 16317 -36168 16553 -35932
rect 16657 -36168 16893 -35932
rect 16997 -36168 17233 -35932
rect 17317 -36168 17553 -35932
rect 17657 -36168 17893 -35932
rect 17997 -36168 18233 -35932
rect 18317 -36168 18553 -35932
rect 18657 -36168 18893 -35932
rect 18997 -36168 19233 -35932
rect 19317 -36168 19553 -35932
rect 19657 -36168 19893 -35932
rect 19997 -36168 20233 -35932
rect 20317 -36168 20553 -35932
rect 20657 -36168 20893 -35932
rect 20997 -36168 21233 -35932
rect 21317 -36168 21553 -35932
rect 21657 -36168 21893 -35932
rect 21997 -36168 22233 -35932
rect 22317 -36168 22553 -35932
rect 22657 -36168 22893 -35932
rect 22997 -36168 23233 -35932
rect 23317 -36168 23553 -35932
rect 23657 -36168 23893 -35932
rect 23997 -36168 24233 -35932
rect 24317 -36168 24553 -35932
rect 24657 -36168 24893 -35932
rect 24997 -36168 25233 -35932
rect 25317 -36168 25553 -35932
rect 25657 -36168 25893 -35932
rect 25997 -36168 26233 -35932
rect 26317 -36168 26553 -35932
rect 26657 -36168 26893 -35932
rect 26997 -36168 27233 -35932
rect 27317 -36168 27553 -35932
rect 27657 -36168 27893 -35932
rect 27997 -36168 28233 -35932
rect 28317 -36168 28553 -35932
rect 28657 -36168 28893 -35932
rect 28997 -36168 29233 -35932
rect 29317 -36168 29553 -35932
rect 29657 -36168 29893 -35932
rect 29997 -36168 30233 -35932
rect 30317 -36168 30553 -35932
rect 30657 -36168 30893 -35932
rect 30997 -36168 31233 -35932
rect 31317 -36168 31553 -35932
rect 31657 -36168 31893 -35932
rect 31997 -36168 32233 -35932
rect 32317 -36168 32553 -35932
rect 32657 -36168 32893 -35932
rect 32997 -36168 33233 -35932
rect 33317 -36168 33553 -35932
rect 33657 -36168 33893 -35932
rect 33997 -36168 34233 -35932
rect 8657 -36508 8893 -36272
rect 8657 -36828 8893 -36592
rect 9657 -36508 9893 -36272
rect 9657 -36828 9893 -36592
rect 10657 -36508 10893 -36272
rect 10657 -36828 10893 -36592
rect 11657 -36508 11893 -36272
rect 11657 -36828 11893 -36592
rect 12657 -36508 12893 -36272
rect 12657 -36828 12893 -36592
rect 13657 -36508 13893 -36272
rect 13657 -36828 13893 -36592
rect 14657 -36508 14893 -36272
rect 14657 -36828 14893 -36592
rect 15657 -36508 15893 -36272
rect 15657 -36828 15893 -36592
rect 16657 -36508 16893 -36272
rect 16657 -36828 16893 -36592
rect 17657 -36508 17893 -36272
rect 17657 -36828 17893 -36592
rect 18657 -36508 18893 -36272
rect 18657 -36828 18893 -36592
rect 19657 -36508 19893 -36272
rect 19657 -36828 19893 -36592
rect 20657 -36508 20893 -36272
rect 20657 -36828 20893 -36592
rect 21657 -36508 21893 -36272
rect 21657 -36828 21893 -36592
rect 22657 -36508 22893 -36272
rect 22657 -36828 22893 -36592
rect 23657 -36508 23893 -36272
rect 23657 -36828 23893 -36592
rect 24657 -36508 24893 -36272
rect 24657 -36828 24893 -36592
rect 25657 -36508 25893 -36272
rect 25657 -36828 25893 -36592
rect 26657 -36508 26893 -36272
rect 26657 -36828 26893 -36592
rect 27657 -36508 27893 -36272
rect 27657 -36828 27893 -36592
rect 28657 -36508 28893 -36272
rect 28657 -36828 28893 -36592
rect 29657 -36508 29893 -36272
rect 29657 -36828 29893 -36592
rect 30657 -36508 30893 -36272
rect 30657 -36828 30893 -36592
rect 31657 -36508 31893 -36272
rect 31657 -36828 31893 -36592
rect 32657 -36508 32893 -36272
rect 32657 -36828 32893 -36592
rect 33657 -36508 33893 -36272
rect 33657 -36828 33893 -36592
rect 8317 -37168 8553 -36932
rect 8657 -37168 8893 -36932
rect 8997 -37168 9233 -36932
rect 9317 -37168 9553 -36932
rect 9657 -37168 9893 -36932
rect 9997 -37168 10233 -36932
rect 10317 -37168 10553 -36932
rect 10657 -37168 10893 -36932
rect 10997 -37168 11233 -36932
rect 11317 -37168 11553 -36932
rect 11657 -37168 11893 -36932
rect 11997 -37168 12233 -36932
rect 12317 -37168 12553 -36932
rect 12657 -37168 12893 -36932
rect 12997 -37168 13233 -36932
rect 13317 -37168 13553 -36932
rect 13657 -37168 13893 -36932
rect 13997 -37168 14233 -36932
rect 14317 -37168 14553 -36932
rect 14657 -37168 14893 -36932
rect 14997 -37168 15233 -36932
rect 15317 -37168 15553 -36932
rect 15657 -37168 15893 -36932
rect 15997 -37168 16233 -36932
rect 16317 -37168 16553 -36932
rect 16657 -37168 16893 -36932
rect 16997 -37168 17233 -36932
rect 17317 -37168 17553 -36932
rect 17657 -37168 17893 -36932
rect 17997 -37168 18233 -36932
rect 18317 -37168 18553 -36932
rect 18657 -37168 18893 -36932
rect 18997 -37168 19233 -36932
rect 19317 -37168 19553 -36932
rect 19657 -37168 19893 -36932
rect 19997 -37168 20233 -36932
rect 20317 -37168 20553 -36932
rect 20657 -37168 20893 -36932
rect 20997 -37168 21233 -36932
rect 21317 -37168 21553 -36932
rect 21657 -37168 21893 -36932
rect 21997 -37168 22233 -36932
rect 22317 -37168 22553 -36932
rect 22657 -37168 22893 -36932
rect 22997 -37168 23233 -36932
rect 23317 -37168 23553 -36932
rect 23657 -37168 23893 -36932
rect 23997 -37168 24233 -36932
rect 24317 -37168 24553 -36932
rect 24657 -37168 24893 -36932
rect 24997 -37168 25233 -36932
rect 25317 -37168 25553 -36932
rect 25657 -37168 25893 -36932
rect 25997 -37168 26233 -36932
rect 26317 -37168 26553 -36932
rect 26657 -37168 26893 -36932
rect 26997 -37168 27233 -36932
rect 27317 -37168 27553 -36932
rect 27657 -37168 27893 -36932
rect 27997 -37168 28233 -36932
rect 28317 -37168 28553 -36932
rect 28657 -37168 28893 -36932
rect 28997 -37168 29233 -36932
rect 29317 -37168 29553 -36932
rect 29657 -37168 29893 -36932
rect 29997 -37168 30233 -36932
rect 30317 -37168 30553 -36932
rect 30657 -37168 30893 -36932
rect 30997 -37168 31233 -36932
rect 31317 -37168 31553 -36932
rect 31657 -37168 31893 -36932
rect 31997 -37168 32233 -36932
rect 32317 -37168 32553 -36932
rect 32657 -37168 32893 -36932
rect 32997 -37168 33233 -36932
rect 33317 -37168 33553 -36932
rect 33657 -37168 33893 -36932
rect 33997 -37168 34233 -36932
rect 8657 -37508 8893 -37272
rect 8657 -37828 8893 -37592
rect 9657 -37508 9893 -37272
rect 9657 -37828 9893 -37592
rect 10657 -37508 10893 -37272
rect 10657 -37828 10893 -37592
rect 11657 -37508 11893 -37272
rect 11657 -37828 11893 -37592
rect 12657 -37508 12893 -37272
rect 12657 -37828 12893 -37592
rect 13657 -37508 13893 -37272
rect 13657 -37828 13893 -37592
rect 14657 -37508 14893 -37272
rect 14657 -37828 14893 -37592
rect 15657 -37508 15893 -37272
rect 15657 -37828 15893 -37592
rect 16657 -37508 16893 -37272
rect 16657 -37828 16893 -37592
rect 17657 -37508 17893 -37272
rect 17657 -37828 17893 -37592
rect 18657 -37508 18893 -37272
rect 18657 -37828 18893 -37592
rect 19657 -37508 19893 -37272
rect 19657 -37828 19893 -37592
rect 20657 -37508 20893 -37272
rect 20657 -37828 20893 -37592
rect 21657 -37508 21893 -37272
rect 21657 -37828 21893 -37592
rect 22657 -37508 22893 -37272
rect 22657 -37828 22893 -37592
rect 23657 -37508 23893 -37272
rect 23657 -37828 23893 -37592
rect 24657 -37508 24893 -37272
rect 24657 -37828 24893 -37592
rect 25657 -37508 25893 -37272
rect 25657 -37828 25893 -37592
rect 26657 -37508 26893 -37272
rect 26657 -37828 26893 -37592
rect 27657 -37508 27893 -37272
rect 27657 -37828 27893 -37592
rect 28657 -37508 28893 -37272
rect 28657 -37828 28893 -37592
rect 29657 -37508 29893 -37272
rect 29657 -37828 29893 -37592
rect 30657 -37508 30893 -37272
rect 30657 -37828 30893 -37592
rect 31657 -37508 31893 -37272
rect 31657 -37828 31893 -37592
rect 32657 -37508 32893 -37272
rect 32657 -37828 32893 -37592
rect 33657 -37508 33893 -37272
rect 33657 -37828 33893 -37592
rect 8317 -38168 8553 -37932
rect 8657 -38168 8893 -37932
rect 8997 -38168 9233 -37932
rect 9317 -38168 9553 -37932
rect 9657 -38168 9893 -37932
rect 9997 -38168 10233 -37932
rect 10317 -38168 10553 -37932
rect 10657 -38168 10893 -37932
rect 10997 -38168 11233 -37932
rect 11317 -38168 11553 -37932
rect 11657 -38168 11893 -37932
rect 11997 -38168 12233 -37932
rect 12317 -38168 12553 -37932
rect 12657 -38168 12893 -37932
rect 12997 -38168 13233 -37932
rect 13317 -38168 13553 -37932
rect 13657 -38168 13893 -37932
rect 13997 -38168 14233 -37932
rect 14317 -38168 14553 -37932
rect 14657 -38168 14893 -37932
rect 14997 -38168 15233 -37932
rect 15317 -38168 15553 -37932
rect 15657 -38168 15893 -37932
rect 15997 -38168 16233 -37932
rect 16317 -38168 16553 -37932
rect 16657 -38168 16893 -37932
rect 16997 -38168 17233 -37932
rect 17317 -38168 17553 -37932
rect 17657 -38168 17893 -37932
rect 17997 -38168 18233 -37932
rect 18317 -38168 18553 -37932
rect 18657 -38168 18893 -37932
rect 18997 -38168 19233 -37932
rect 19317 -38168 19553 -37932
rect 19657 -38168 19893 -37932
rect 19997 -38168 20233 -37932
rect 20317 -38168 20553 -37932
rect 20657 -38168 20893 -37932
rect 20997 -38168 21233 -37932
rect 21317 -38168 21553 -37932
rect 21657 -38168 21893 -37932
rect 21997 -38168 22233 -37932
rect 22317 -38168 22553 -37932
rect 22657 -38168 22893 -37932
rect 22997 -38168 23233 -37932
rect 23317 -38168 23553 -37932
rect 23657 -38168 23893 -37932
rect 23997 -38168 24233 -37932
rect 24317 -38168 24553 -37932
rect 24657 -38168 24893 -37932
rect 24997 -38168 25233 -37932
rect 25317 -38168 25553 -37932
rect 25657 -38168 25893 -37932
rect 25997 -38168 26233 -37932
rect 26317 -38168 26553 -37932
rect 26657 -38168 26893 -37932
rect 26997 -38168 27233 -37932
rect 27317 -38168 27553 -37932
rect 27657 -38168 27893 -37932
rect 27997 -38168 28233 -37932
rect 28317 -38168 28553 -37932
rect 28657 -38168 28893 -37932
rect 28997 -38168 29233 -37932
rect 29317 -38168 29553 -37932
rect 29657 -38168 29893 -37932
rect 29997 -38168 30233 -37932
rect 30317 -38168 30553 -37932
rect 30657 -38168 30893 -37932
rect 30997 -38168 31233 -37932
rect 31317 -38168 31553 -37932
rect 31657 -38168 31893 -37932
rect 31997 -38168 32233 -37932
rect 32317 -38168 32553 -37932
rect 32657 -38168 32893 -37932
rect 32997 -38168 33233 -37932
rect 33317 -38168 33553 -37932
rect 33657 -38168 33893 -37932
rect 33997 -38168 34233 -37932
rect 8657 -38508 8893 -38272
rect 8657 -38828 8893 -38592
rect 9657 -38508 9893 -38272
rect 9657 -38828 9893 -38592
rect 10657 -38508 10893 -38272
rect 10657 -38828 10893 -38592
rect 11657 -38508 11893 -38272
rect 11657 -38828 11893 -38592
rect 12657 -38508 12893 -38272
rect 12657 -38828 12893 -38592
rect 13657 -38508 13893 -38272
rect 13657 -38828 13893 -38592
rect 14657 -38508 14893 -38272
rect 14657 -38828 14893 -38592
rect 15657 -38508 15893 -38272
rect 15657 -38828 15893 -38592
rect 16657 -38508 16893 -38272
rect 16657 -38828 16893 -38592
rect 17657 -38508 17893 -38272
rect 17657 -38828 17893 -38592
rect 18657 -38508 18893 -38272
rect 18657 -38828 18893 -38592
rect 19657 -38508 19893 -38272
rect 19657 -38828 19893 -38592
rect 20657 -38508 20893 -38272
rect 20657 -38828 20893 -38592
rect 21657 -38508 21893 -38272
rect 21657 -38828 21893 -38592
rect 22657 -38508 22893 -38272
rect 22657 -38828 22893 -38592
rect 23657 -38508 23893 -38272
rect 23657 -38828 23893 -38592
rect 24657 -38508 24893 -38272
rect 24657 -38828 24893 -38592
rect 25657 -38508 25893 -38272
rect 25657 -38828 25893 -38592
rect 26657 -38508 26893 -38272
rect 26657 -38828 26893 -38592
rect 27657 -38508 27893 -38272
rect 27657 -38828 27893 -38592
rect 28657 -38508 28893 -38272
rect 28657 -38828 28893 -38592
rect 29657 -38508 29893 -38272
rect 29657 -38828 29893 -38592
rect 30657 -38508 30893 -38272
rect 30657 -38828 30893 -38592
rect 31657 -38508 31893 -38272
rect 31657 -38828 31893 -38592
rect 32657 -38508 32893 -38272
rect 32657 -38828 32893 -38592
rect 33657 -38508 33893 -38272
rect 33657 -38828 33893 -38592
rect 8317 -39168 8553 -38932
rect 8657 -39168 8893 -38932
rect 8997 -39168 9233 -38932
rect 9317 -39168 9553 -38932
rect 9657 -39168 9893 -38932
rect 9997 -39168 10233 -38932
rect 10317 -39168 10553 -38932
rect 10657 -39168 10893 -38932
rect 10997 -39168 11233 -38932
rect 11317 -39168 11553 -38932
rect 11657 -39168 11893 -38932
rect 11997 -39168 12233 -38932
rect 12317 -39168 12553 -38932
rect 12657 -39168 12893 -38932
rect 12997 -39168 13233 -38932
rect 13317 -39168 13553 -38932
rect 13657 -39168 13893 -38932
rect 13997 -39168 14233 -38932
rect 14317 -39168 14553 -38932
rect 14657 -39168 14893 -38932
rect 14997 -39168 15233 -38932
rect 15317 -39168 15553 -38932
rect 15657 -39168 15893 -38932
rect 15997 -39168 16233 -38932
rect 16317 -39168 16553 -38932
rect 16657 -39168 16893 -38932
rect 16997 -39168 17233 -38932
rect 17317 -39168 17553 -38932
rect 17657 -39168 17893 -38932
rect 17997 -39168 18233 -38932
rect 18317 -39168 18553 -38932
rect 18657 -39168 18893 -38932
rect 18997 -39168 19233 -38932
rect 19317 -39168 19553 -38932
rect 19657 -39168 19893 -38932
rect 19997 -39168 20233 -38932
rect 20317 -39168 20553 -38932
rect 20657 -39168 20893 -38932
rect 20997 -39168 21233 -38932
rect 21317 -39168 21553 -38932
rect 21657 -39168 21893 -38932
rect 21997 -39168 22233 -38932
rect 22317 -39168 22553 -38932
rect 22657 -39168 22893 -38932
rect 22997 -39168 23233 -38932
rect 23317 -39168 23553 -38932
rect 23657 -39168 23893 -38932
rect 23997 -39168 24233 -38932
rect 24317 -39168 24553 -38932
rect 24657 -39168 24893 -38932
rect 24997 -39168 25233 -38932
rect 25317 -39168 25553 -38932
rect 25657 -39168 25893 -38932
rect 25997 -39168 26233 -38932
rect 26317 -39168 26553 -38932
rect 26657 -39168 26893 -38932
rect 26997 -39168 27233 -38932
rect 27317 -39168 27553 -38932
rect 27657 -39168 27893 -38932
rect 27997 -39168 28233 -38932
rect 28317 -39168 28553 -38932
rect 28657 -39168 28893 -38932
rect 28997 -39168 29233 -38932
rect 29317 -39168 29553 -38932
rect 29657 -39168 29893 -38932
rect 29997 -39168 30233 -38932
rect 30317 -39168 30553 -38932
rect 30657 -39168 30893 -38932
rect 30997 -39168 31233 -38932
rect 31317 -39168 31553 -38932
rect 31657 -39168 31893 -38932
rect 31997 -39168 32233 -38932
rect 32317 -39168 32553 -38932
rect 32657 -39168 32893 -38932
rect 32997 -39168 33233 -38932
rect 33317 -39168 33553 -38932
rect 33657 -39168 33893 -38932
rect 33997 -39168 34233 -38932
rect 8657 -39508 8893 -39272
rect 8657 -39828 8893 -39592
rect 9657 -39508 9893 -39272
rect 9657 -39828 9893 -39592
rect 10657 -39508 10893 -39272
rect 10657 -39828 10893 -39592
rect 11657 -39508 11893 -39272
rect 11657 -39828 11893 -39592
rect 12657 -39508 12893 -39272
rect 12657 -39828 12893 -39592
rect 13657 -39508 13893 -39272
rect 13657 -39828 13893 -39592
rect 14657 -39508 14893 -39272
rect 14657 -39828 14893 -39592
rect 15657 -39508 15893 -39272
rect 15657 -39828 15893 -39592
rect 16657 -39508 16893 -39272
rect 16657 -39828 16893 -39592
rect 17657 -39508 17893 -39272
rect 17657 -39828 17893 -39592
rect 18657 -39508 18893 -39272
rect 18657 -39828 18893 -39592
rect 19657 -39508 19893 -39272
rect 19657 -39828 19893 -39592
rect 20657 -39508 20893 -39272
rect 20657 -39828 20893 -39592
rect 21657 -39508 21893 -39272
rect 21657 -39828 21893 -39592
rect 22657 -39508 22893 -39272
rect 22657 -39828 22893 -39592
rect 23657 -39508 23893 -39272
rect 23657 -39828 23893 -39592
rect 24657 -39508 24893 -39272
rect 24657 -39828 24893 -39592
rect 25657 -39508 25893 -39272
rect 25657 -39828 25893 -39592
rect 26657 -39508 26893 -39272
rect 26657 -39828 26893 -39592
rect 27657 -39508 27893 -39272
rect 27657 -39828 27893 -39592
rect 28657 -39508 28893 -39272
rect 28657 -39828 28893 -39592
rect 29657 -39508 29893 -39272
rect 29657 -39828 29893 -39592
rect 30657 -39508 30893 -39272
rect 30657 -39828 30893 -39592
rect 31657 -39508 31893 -39272
rect 31657 -39828 31893 -39592
rect 32657 -39508 32893 -39272
rect 32657 -39828 32893 -39592
rect 33657 -39508 33893 -39272
rect 33657 -39828 33893 -39592
rect 8317 -40168 8553 -39932
rect 8657 -40168 8893 -39932
rect 8997 -40168 9233 -39932
rect 9317 -40168 9553 -39932
rect 9657 -40168 9893 -39932
rect 9997 -40168 10233 -39932
rect 10317 -40168 10553 -39932
rect 10657 -40168 10893 -39932
rect 10997 -40168 11233 -39932
rect 11317 -40168 11553 -39932
rect 11657 -40168 11893 -39932
rect 11997 -40168 12233 -39932
rect 12317 -40168 12553 -39932
rect 12657 -40168 12893 -39932
rect 12997 -40168 13233 -39932
rect 13317 -40168 13553 -39932
rect 13657 -40168 13893 -39932
rect 13997 -40168 14233 -39932
rect 14317 -40168 14553 -39932
rect 14657 -40168 14893 -39932
rect 14997 -40168 15233 -39932
rect 15317 -40168 15553 -39932
rect 15657 -40168 15893 -39932
rect 15997 -40168 16233 -39932
rect 16317 -40168 16553 -39932
rect 16657 -40168 16893 -39932
rect 16997 -40168 17233 -39932
rect 17317 -40168 17553 -39932
rect 17657 -40168 17893 -39932
rect 17997 -40168 18233 -39932
rect 18317 -40168 18553 -39932
rect 18657 -40168 18893 -39932
rect 18997 -40168 19233 -39932
rect 19317 -40168 19553 -39932
rect 19657 -40168 19893 -39932
rect 19997 -40168 20233 -39932
rect 20317 -40168 20553 -39932
rect 20657 -40168 20893 -39932
rect 20997 -40168 21233 -39932
rect 21317 -40168 21553 -39932
rect 21657 -40168 21893 -39932
rect 21997 -40168 22233 -39932
rect 22317 -40168 22553 -39932
rect 22657 -40168 22893 -39932
rect 22997 -40168 23233 -39932
rect 23317 -40168 23553 -39932
rect 23657 -40168 23893 -39932
rect 23997 -40168 24233 -39932
rect 24317 -40168 24553 -39932
rect 24657 -40168 24893 -39932
rect 24997 -40168 25233 -39932
rect 25317 -40168 25553 -39932
rect 25657 -40168 25893 -39932
rect 25997 -40168 26233 -39932
rect 26317 -40168 26553 -39932
rect 26657 -40168 26893 -39932
rect 26997 -40168 27233 -39932
rect 27317 -40168 27553 -39932
rect 27657 -40168 27893 -39932
rect 27997 -40168 28233 -39932
rect 28317 -40168 28553 -39932
rect 28657 -40168 28893 -39932
rect 28997 -40168 29233 -39932
rect 29317 -40168 29553 -39932
rect 29657 -40168 29893 -39932
rect 29997 -40168 30233 -39932
rect 30317 -40168 30553 -39932
rect 30657 -40168 30893 -39932
rect 30997 -40168 31233 -39932
rect 31317 -40168 31553 -39932
rect 31657 -40168 31893 -39932
rect 31997 -40168 32233 -39932
rect 32317 -40168 32553 -39932
rect 32657 -40168 32893 -39932
rect 32997 -40168 33233 -39932
rect 33317 -40168 33553 -39932
rect 33657 -40168 33893 -39932
rect 33997 -40168 34233 -39932
rect 8657 -40508 8893 -40272
rect 8657 -40828 8893 -40592
rect 9657 -40508 9893 -40272
rect 9657 -40828 9893 -40592
rect 10657 -40508 10893 -40272
rect 10657 -40828 10893 -40592
rect 11657 -40508 11893 -40272
rect 11657 -40828 11893 -40592
rect 12657 -40508 12893 -40272
rect 12657 -40828 12893 -40592
rect 13657 -40508 13893 -40272
rect 13657 -40828 13893 -40592
rect 14657 -40508 14893 -40272
rect 14657 -40828 14893 -40592
rect 15657 -40508 15893 -40272
rect 15657 -40828 15893 -40592
rect 16657 -40508 16893 -40272
rect 16657 -40828 16893 -40592
rect 17657 -40508 17893 -40272
rect 17657 -40828 17893 -40592
rect 18657 -40508 18893 -40272
rect 18657 -40828 18893 -40592
rect 19657 -40508 19893 -40272
rect 19657 -40828 19893 -40592
rect 20657 -40508 20893 -40272
rect 20657 -40828 20893 -40592
rect 21657 -40508 21893 -40272
rect 21657 -40828 21893 -40592
rect 22657 -40508 22893 -40272
rect 22657 -40828 22893 -40592
rect 23657 -40508 23893 -40272
rect 23657 -40828 23893 -40592
rect 24657 -40508 24893 -40272
rect 24657 -40828 24893 -40592
rect 25657 -40508 25893 -40272
rect 25657 -40828 25893 -40592
rect 26657 -40508 26893 -40272
rect 26657 -40828 26893 -40592
rect 27657 -40508 27893 -40272
rect 27657 -40828 27893 -40592
rect 28657 -40508 28893 -40272
rect 28657 -40828 28893 -40592
rect 29657 -40508 29893 -40272
rect 29657 -40828 29893 -40592
rect 30657 -40508 30893 -40272
rect 30657 -40828 30893 -40592
rect 31657 -40508 31893 -40272
rect 31657 -40828 31893 -40592
rect 32657 -40508 32893 -40272
rect 32657 -40828 32893 -40592
rect 33657 -40508 33893 -40272
rect 33657 -40828 33893 -40592
rect 8317 -41168 8553 -40932
rect 8657 -41168 8893 -40932
rect 8997 -41168 9233 -40932
rect 9317 -41168 9553 -40932
rect 9657 -41168 9893 -40932
rect 9997 -41168 10233 -40932
rect 10317 -41168 10553 -40932
rect 10657 -41168 10893 -40932
rect 10997 -41168 11233 -40932
rect 11317 -41168 11553 -40932
rect 11657 -41168 11893 -40932
rect 11997 -41168 12233 -40932
rect 12317 -41168 12553 -40932
rect 12657 -41168 12893 -40932
rect 12997 -41168 13233 -40932
rect 13317 -41168 13553 -40932
rect 13657 -41168 13893 -40932
rect 13997 -41168 14233 -40932
rect 14317 -41168 14553 -40932
rect 14657 -41168 14893 -40932
rect 14997 -41168 15233 -40932
rect 15317 -41168 15553 -40932
rect 15657 -41168 15893 -40932
rect 15997 -41168 16233 -40932
rect 16317 -41168 16553 -40932
rect 16657 -41168 16893 -40932
rect 16997 -41168 17233 -40932
rect 17317 -41168 17553 -40932
rect 17657 -41168 17893 -40932
rect 17997 -41168 18233 -40932
rect 18317 -41168 18553 -40932
rect 18657 -41168 18893 -40932
rect 18997 -41168 19233 -40932
rect 19317 -41168 19553 -40932
rect 19657 -41168 19893 -40932
rect 19997 -41168 20233 -40932
rect 20317 -41168 20553 -40932
rect 20657 -41168 20893 -40932
rect 20997 -41168 21233 -40932
rect 21317 -41168 21553 -40932
rect 21657 -41168 21893 -40932
rect 21997 -41168 22233 -40932
rect 22317 -41168 22553 -40932
rect 22657 -41168 22893 -40932
rect 22997 -41168 23233 -40932
rect 23317 -41168 23553 -40932
rect 23657 -41168 23893 -40932
rect 23997 -41168 24233 -40932
rect 24317 -41168 24553 -40932
rect 24657 -41168 24893 -40932
rect 24997 -41168 25233 -40932
rect 25317 -41168 25553 -40932
rect 25657 -41168 25893 -40932
rect 25997 -41168 26233 -40932
rect 26317 -41168 26553 -40932
rect 26657 -41168 26893 -40932
rect 26997 -41168 27233 -40932
rect 27317 -41168 27553 -40932
rect 27657 -41168 27893 -40932
rect 27997 -41168 28233 -40932
rect 28317 -41168 28553 -40932
rect 28657 -41168 28893 -40932
rect 28997 -41168 29233 -40932
rect 29317 -41168 29553 -40932
rect 29657 -41168 29893 -40932
rect 29997 -41168 30233 -40932
rect 30317 -41168 30553 -40932
rect 30657 -41168 30893 -40932
rect 30997 -41168 31233 -40932
rect 31317 -41168 31553 -40932
rect 31657 -41168 31893 -40932
rect 31997 -41168 32233 -40932
rect 32317 -41168 32553 -40932
rect 32657 -41168 32893 -40932
rect 32997 -41168 33233 -40932
rect 33317 -41168 33553 -40932
rect 33657 -41168 33893 -40932
rect 33997 -41168 34233 -40932
rect 8657 -41508 8893 -41272
rect 8657 -41828 8893 -41592
rect 9657 -41508 9893 -41272
rect 9657 -41828 9893 -41592
rect 10657 -41508 10893 -41272
rect 10657 -41828 10893 -41592
rect 11657 -41508 11893 -41272
rect 11657 -41828 11893 -41592
rect 12657 -41508 12893 -41272
rect 12657 -41828 12893 -41592
rect 13657 -41508 13893 -41272
rect 13657 -41828 13893 -41592
rect 14657 -41508 14893 -41272
rect 14657 -41828 14893 -41592
rect 15657 -41508 15893 -41272
rect 15657 -41828 15893 -41592
rect 16657 -41508 16893 -41272
rect 16657 -41828 16893 -41592
rect 17657 -41508 17893 -41272
rect 17657 -41828 17893 -41592
rect 18657 -41508 18893 -41272
rect 18657 -41828 18893 -41592
rect 19657 -41508 19893 -41272
rect 19657 -41828 19893 -41592
rect 20657 -41508 20893 -41272
rect 20657 -41828 20893 -41592
rect 21657 -41508 21893 -41272
rect 21657 -41828 21893 -41592
rect 22657 -41508 22893 -41272
rect 22657 -41828 22893 -41592
rect 23657 -41508 23893 -41272
rect 23657 -41828 23893 -41592
rect 24657 -41508 24893 -41272
rect 24657 -41828 24893 -41592
rect 25657 -41508 25893 -41272
rect 25657 -41828 25893 -41592
rect 26657 -41508 26893 -41272
rect 26657 -41828 26893 -41592
rect 27657 -41508 27893 -41272
rect 27657 -41828 27893 -41592
rect 28657 -41508 28893 -41272
rect 28657 -41828 28893 -41592
rect 29657 -41508 29893 -41272
rect 29657 -41828 29893 -41592
rect 30657 -41508 30893 -41272
rect 30657 -41828 30893 -41592
rect 31657 -41508 31893 -41272
rect 31657 -41828 31893 -41592
rect 32657 -41508 32893 -41272
rect 32657 -41828 32893 -41592
rect 33657 -41508 33893 -41272
rect 33657 -41828 33893 -41592
rect 8317 -42168 8553 -41932
rect 8657 -42168 8893 -41932
rect 8997 -42168 9233 -41932
rect 9317 -42168 9553 -41932
rect 9657 -42168 9893 -41932
rect 9997 -42168 10233 -41932
rect 10317 -42168 10553 -41932
rect 10657 -42168 10893 -41932
rect 10997 -42168 11233 -41932
rect 11317 -42168 11553 -41932
rect 11657 -42168 11893 -41932
rect 11997 -42168 12233 -41932
rect 12317 -42168 12553 -41932
rect 12657 -42168 12893 -41932
rect 12997 -42168 13233 -41932
rect 13317 -42168 13553 -41932
rect 13657 -42168 13893 -41932
rect 13997 -42168 14233 -41932
rect 14317 -42168 14553 -41932
rect 14657 -42168 14893 -41932
rect 14997 -42168 15233 -41932
rect 15317 -42168 15553 -41932
rect 15657 -42168 15893 -41932
rect 15997 -42168 16233 -41932
rect 16317 -42168 16553 -41932
rect 16657 -42168 16893 -41932
rect 16997 -42168 17233 -41932
rect 17317 -42168 17553 -41932
rect 17657 -42168 17893 -41932
rect 17997 -42168 18233 -41932
rect 18317 -42168 18553 -41932
rect 18657 -42168 18893 -41932
rect 18997 -42168 19233 -41932
rect 19317 -42168 19553 -41932
rect 19657 -42168 19893 -41932
rect 19997 -42168 20233 -41932
rect 20317 -42168 20553 -41932
rect 20657 -42168 20893 -41932
rect 20997 -42168 21233 -41932
rect 21317 -42168 21553 -41932
rect 21657 -42168 21893 -41932
rect 21997 -42168 22233 -41932
rect 22317 -42168 22553 -41932
rect 22657 -42168 22893 -41932
rect 22997 -42168 23233 -41932
rect 23317 -42168 23553 -41932
rect 23657 -42168 23893 -41932
rect 23997 -42168 24233 -41932
rect 24317 -42168 24553 -41932
rect 24657 -42168 24893 -41932
rect 24997 -42168 25233 -41932
rect 25317 -42168 25553 -41932
rect 25657 -42168 25893 -41932
rect 25997 -42168 26233 -41932
rect 26317 -42168 26553 -41932
rect 26657 -42168 26893 -41932
rect 26997 -42168 27233 -41932
rect 27317 -42168 27553 -41932
rect 27657 -42168 27893 -41932
rect 27997 -42168 28233 -41932
rect 28317 -42168 28553 -41932
rect 28657 -42168 28893 -41932
rect 28997 -42168 29233 -41932
rect 29317 -42168 29553 -41932
rect 29657 -42168 29893 -41932
rect 29997 -42168 30233 -41932
rect 30317 -42168 30553 -41932
rect 30657 -42168 30893 -41932
rect 30997 -42168 31233 -41932
rect 31317 -42168 31553 -41932
rect 31657 -42168 31893 -41932
rect 31997 -42168 32233 -41932
rect 32317 -42168 32553 -41932
rect 32657 -42168 32893 -41932
rect 32997 -42168 33233 -41932
rect 33317 -42168 33553 -41932
rect 33657 -42168 33893 -41932
rect 33997 -42168 34233 -41932
rect 8657 -42508 8893 -42272
rect 8657 -42828 8893 -42592
rect 9657 -42508 9893 -42272
rect 9657 -42828 9893 -42592
rect 10657 -42508 10893 -42272
rect 10657 -42828 10893 -42592
rect 11657 -42508 11893 -42272
rect 11657 -42828 11893 -42592
rect 12657 -42508 12893 -42272
rect 12657 -42828 12893 -42592
rect 13657 -42508 13893 -42272
rect 13657 -42828 13893 -42592
rect 14657 -42508 14893 -42272
rect 14657 -42828 14893 -42592
rect 15657 -42508 15893 -42272
rect 15657 -42828 15893 -42592
rect 16657 -42508 16893 -42272
rect 16657 -42828 16893 -42592
rect 17657 -42508 17893 -42272
rect 17657 -42828 17893 -42592
rect 18657 -42508 18893 -42272
rect 18657 -42828 18893 -42592
rect 19657 -42508 19893 -42272
rect 19657 -42828 19893 -42592
rect 20657 -42508 20893 -42272
rect 20657 -42828 20893 -42592
rect 21657 -42508 21893 -42272
rect 21657 -42828 21893 -42592
rect 22657 -42508 22893 -42272
rect 22657 -42828 22893 -42592
rect 23657 -42508 23893 -42272
rect 23657 -42828 23893 -42592
rect 24657 -42508 24893 -42272
rect 24657 -42828 24893 -42592
rect 25657 -42508 25893 -42272
rect 25657 -42828 25893 -42592
rect 26657 -42508 26893 -42272
rect 26657 -42828 26893 -42592
rect 27657 -42508 27893 -42272
rect 27657 -42828 27893 -42592
rect 28657 -42508 28893 -42272
rect 28657 -42828 28893 -42592
rect 29657 -42508 29893 -42272
rect 29657 -42828 29893 -42592
rect 30657 -42508 30893 -42272
rect 30657 -42828 30893 -42592
rect 31657 -42508 31893 -42272
rect 31657 -42828 31893 -42592
rect 32657 -42508 32893 -42272
rect 32657 -42828 32893 -42592
rect 33657 -42508 33893 -42272
rect 33657 -42828 33893 -42592
rect 8317 -43168 8553 -42932
rect 8657 -43168 8893 -42932
rect 8997 -43168 9233 -42932
rect 9317 -43168 9553 -42932
rect 9657 -43168 9893 -42932
rect 9997 -43168 10233 -42932
rect 10317 -43168 10553 -42932
rect 10657 -43168 10893 -42932
rect 10997 -43168 11233 -42932
rect 11317 -43168 11553 -42932
rect 11657 -43168 11893 -42932
rect 11997 -43168 12233 -42932
rect 12317 -43168 12553 -42932
rect 12657 -43168 12893 -42932
rect 12997 -43168 13233 -42932
rect 13317 -43168 13553 -42932
rect 13657 -43168 13893 -42932
rect 13997 -43168 14233 -42932
rect 14317 -43168 14553 -42932
rect 14657 -43168 14893 -42932
rect 14997 -43168 15233 -42932
rect 15317 -43168 15553 -42932
rect 15657 -43168 15893 -42932
rect 15997 -43168 16233 -42932
rect 16317 -43168 16553 -42932
rect 16657 -43168 16893 -42932
rect 16997 -43168 17233 -42932
rect 17317 -43168 17553 -42932
rect 17657 -43168 17893 -42932
rect 17997 -43168 18233 -42932
rect 18317 -43168 18553 -42932
rect 18657 -43168 18893 -42932
rect 18997 -43168 19233 -42932
rect 19317 -43168 19553 -42932
rect 19657 -43168 19893 -42932
rect 19997 -43168 20233 -42932
rect 20317 -43168 20553 -42932
rect 20657 -43168 20893 -42932
rect 20997 -43168 21233 -42932
rect 21317 -43168 21553 -42932
rect 21657 -43168 21893 -42932
rect 21997 -43168 22233 -42932
rect 22317 -43168 22553 -42932
rect 22657 -43168 22893 -42932
rect 22997 -43168 23233 -42932
rect 23317 -43168 23553 -42932
rect 23657 -43168 23893 -42932
rect 23997 -43168 24233 -42932
rect 24317 -43168 24553 -42932
rect 24657 -43168 24893 -42932
rect 24997 -43168 25233 -42932
rect 25317 -43168 25553 -42932
rect 25657 -43168 25893 -42932
rect 25997 -43168 26233 -42932
rect 26317 -43168 26553 -42932
rect 26657 -43168 26893 -42932
rect 26997 -43168 27233 -42932
rect 27317 -43168 27553 -42932
rect 27657 -43168 27893 -42932
rect 27997 -43168 28233 -42932
rect 28317 -43168 28553 -42932
rect 28657 -43168 28893 -42932
rect 28997 -43168 29233 -42932
rect 29317 -43168 29553 -42932
rect 29657 -43168 29893 -42932
rect 29997 -43168 30233 -42932
rect 30317 -43168 30553 -42932
rect 30657 -43168 30893 -42932
rect 30997 -43168 31233 -42932
rect 31317 -43168 31553 -42932
rect 31657 -43168 31893 -42932
rect 31997 -43168 32233 -42932
rect 32317 -43168 32553 -42932
rect 32657 -43168 32893 -42932
rect 32997 -43168 33233 -42932
rect 33317 -43168 33553 -42932
rect 33657 -43168 33893 -42932
rect 33997 -43168 34233 -42932
rect 8657 -43508 8893 -43272
rect 8657 -43828 8893 -43592
rect 9657 -43508 9893 -43272
rect 9657 -43828 9893 -43592
rect 10657 -43508 10893 -43272
rect 10657 -43828 10893 -43592
rect 11657 -43508 11893 -43272
rect 11657 -43828 11893 -43592
rect 12657 -43508 12893 -43272
rect 12657 -43828 12893 -43592
rect 13657 -43508 13893 -43272
rect 13657 -43828 13893 -43592
rect 14657 -43508 14893 -43272
rect 14657 -43828 14893 -43592
rect 15657 -43508 15893 -43272
rect 15657 -43828 15893 -43592
rect 16657 -43508 16893 -43272
rect 16657 -43828 16893 -43592
rect 17657 -43508 17893 -43272
rect 17657 -43828 17893 -43592
rect 18657 -43508 18893 -43272
rect 18657 -43828 18893 -43592
rect 19657 -43508 19893 -43272
rect 19657 -43828 19893 -43592
rect 20657 -43508 20893 -43272
rect 20657 -43828 20893 -43592
rect 21657 -43508 21893 -43272
rect 21657 -43828 21893 -43592
rect 22657 -43508 22893 -43272
rect 22657 -43828 22893 -43592
rect 23657 -43508 23893 -43272
rect 23657 -43828 23893 -43592
rect 24657 -43508 24893 -43272
rect 24657 -43828 24893 -43592
rect 25657 -43508 25893 -43272
rect 25657 -43828 25893 -43592
rect 26657 -43508 26893 -43272
rect 26657 -43828 26893 -43592
rect 27657 -43508 27893 -43272
rect 27657 -43828 27893 -43592
rect 28657 -43508 28893 -43272
rect 28657 -43828 28893 -43592
rect 29657 -43508 29893 -43272
rect 29657 -43828 29893 -43592
rect 30657 -43508 30893 -43272
rect 30657 -43828 30893 -43592
rect 31657 -43508 31893 -43272
rect 31657 -43828 31893 -43592
rect 32657 -43508 32893 -43272
rect 32657 -43828 32893 -43592
rect 33657 -43508 33893 -43272
rect 33657 -43828 33893 -43592
rect 8317 -44168 8553 -43932
rect 8657 -44168 8893 -43932
rect 8997 -44168 9233 -43932
rect 9317 -44168 9553 -43932
rect 9657 -44168 9893 -43932
rect 9997 -44168 10233 -43932
rect 10317 -44168 10553 -43932
rect 10657 -44168 10893 -43932
rect 10997 -44168 11233 -43932
rect 11317 -44168 11553 -43932
rect 11657 -44168 11893 -43932
rect 11997 -44168 12233 -43932
rect 12317 -44168 12553 -43932
rect 12657 -44168 12893 -43932
rect 12997 -44168 13233 -43932
rect 13317 -44168 13553 -43932
rect 13657 -44168 13893 -43932
rect 13997 -44168 14233 -43932
rect 14317 -44168 14553 -43932
rect 14657 -44168 14893 -43932
rect 14997 -44168 15233 -43932
rect 15317 -44168 15553 -43932
rect 15657 -44168 15893 -43932
rect 15997 -44168 16233 -43932
rect 16317 -44168 16553 -43932
rect 16657 -44168 16893 -43932
rect 16997 -44168 17233 -43932
rect 17317 -44168 17553 -43932
rect 17657 -44168 17893 -43932
rect 17997 -44168 18233 -43932
rect 18317 -44168 18553 -43932
rect 18657 -44168 18893 -43932
rect 18997 -44168 19233 -43932
rect 19317 -44168 19553 -43932
rect 19657 -44168 19893 -43932
rect 19997 -44168 20233 -43932
rect 20317 -44168 20553 -43932
rect 20657 -44168 20893 -43932
rect 20997 -44168 21233 -43932
rect 21317 -44168 21553 -43932
rect 21657 -44168 21893 -43932
rect 21997 -44168 22233 -43932
rect 22317 -44168 22553 -43932
rect 22657 -44168 22893 -43932
rect 22997 -44168 23233 -43932
rect 23317 -44168 23553 -43932
rect 23657 -44168 23893 -43932
rect 23997 -44168 24233 -43932
rect 24317 -44168 24553 -43932
rect 24657 -44168 24893 -43932
rect 24997 -44168 25233 -43932
rect 25317 -44168 25553 -43932
rect 25657 -44168 25893 -43932
rect 25997 -44168 26233 -43932
rect 26317 -44168 26553 -43932
rect 26657 -44168 26893 -43932
rect 26997 -44168 27233 -43932
rect 27317 -44168 27553 -43932
rect 27657 -44168 27893 -43932
rect 27997 -44168 28233 -43932
rect 28317 -44168 28553 -43932
rect 28657 -44168 28893 -43932
rect 28997 -44168 29233 -43932
rect 29317 -44168 29553 -43932
rect 29657 -44168 29893 -43932
rect 29997 -44168 30233 -43932
rect 30317 -44168 30553 -43932
rect 30657 -44168 30893 -43932
rect 30997 -44168 31233 -43932
rect 31317 -44168 31553 -43932
rect 31657 -44168 31893 -43932
rect 31997 -44168 32233 -43932
rect 32317 -44168 32553 -43932
rect 32657 -44168 32893 -43932
rect 32997 -44168 33233 -43932
rect 33317 -44168 33553 -43932
rect 33657 -44168 33893 -43932
rect 33997 -44168 34233 -43932
rect 8657 -44508 8893 -44272
rect 8657 -44828 8893 -44592
rect 9657 -44508 9893 -44272
rect 9657 -44828 9893 -44592
rect 10657 -44508 10893 -44272
rect 10657 -44828 10893 -44592
rect 11657 -44508 11893 -44272
rect 11657 -44828 11893 -44592
rect 12657 -44508 12893 -44272
rect 12657 -44828 12893 -44592
rect 13657 -44508 13893 -44272
rect 13657 -44828 13893 -44592
rect 14657 -44508 14893 -44272
rect 14657 -44828 14893 -44592
rect 15657 -44508 15893 -44272
rect 15657 -44828 15893 -44592
rect 16657 -44508 16893 -44272
rect 16657 -44828 16893 -44592
rect 17657 -44508 17893 -44272
rect 17657 -44828 17893 -44592
rect 18657 -44508 18893 -44272
rect 18657 -44828 18893 -44592
rect 19657 -44508 19893 -44272
rect 19657 -44828 19893 -44592
rect 20657 -44508 20893 -44272
rect 20657 -44828 20893 -44592
rect 21657 -44508 21893 -44272
rect 21657 -44828 21893 -44592
rect 22657 -44508 22893 -44272
rect 22657 -44828 22893 -44592
rect 23657 -44508 23893 -44272
rect 23657 -44828 23893 -44592
rect 24657 -44508 24893 -44272
rect 24657 -44828 24893 -44592
rect 25657 -44508 25893 -44272
rect 25657 -44828 25893 -44592
rect 26657 -44508 26893 -44272
rect 26657 -44828 26893 -44592
rect 27657 -44508 27893 -44272
rect 27657 -44828 27893 -44592
rect 28657 -44508 28893 -44272
rect 28657 -44828 28893 -44592
rect 29657 -44508 29893 -44272
rect 29657 -44828 29893 -44592
rect 30657 -44508 30893 -44272
rect 30657 -44828 30893 -44592
rect 31657 -44508 31893 -44272
rect 31657 -44828 31893 -44592
rect 32657 -44508 32893 -44272
rect 32657 -44828 32893 -44592
rect 33657 -44508 33893 -44272
rect 33657 -44828 33893 -44592
rect -74783 -45168 -74547 -44932
rect -74443 -45168 -74207 -44932
rect -74103 -45168 -73867 -44932
rect -73783 -45168 -73547 -44932
rect -73443 -45168 -73207 -44932
rect -73103 -45168 -72867 -44932
rect -72783 -45168 -72547 -44932
rect -72443 -45168 -72207 -44932
rect -72103 -45168 -71867 -44932
rect -71783 -45168 -71547 -44932
rect -71443 -45168 -71207 -44932
rect -71103 -45168 -70867 -44932
rect -70783 -45168 -70547 -44932
rect -70443 -45168 -70207 -44932
rect -70103 -45168 -69867 -44932
rect -69783 -45168 -69547 -44932
rect -69443 -45168 -69207 -44932
rect -69103 -45168 -68867 -44932
rect -68783 -45168 -68547 -44932
rect -68443 -45168 -68207 -44932
rect -68103 -45168 -67867 -44932
rect -67783 -45168 -67547 -44932
rect -67443 -45168 -67207 -44932
rect -67103 -45168 -66867 -44932
rect -66783 -45168 -66547 -44932
rect -66443 -45168 -66207 -44932
rect -66103 -45168 -65867 -44932
rect -65783 -45168 -65547 -44932
rect -65443 -45168 -65207 -44932
rect -65103 -45168 -64867 -44932
rect -64783 -45168 -64547 -44932
rect -64443 -45168 -64207 -44932
rect -64103 -45168 -63867 -44932
rect -63783 -45168 -63547 -44932
rect -63443 -45168 -63207 -44932
rect -63103 -45168 -62867 -44932
rect -62783 -45168 -62547 -44932
rect -62443 -45168 -62207 -44932
rect -62103 -45168 -61867 -44932
rect -61783 -45168 -61547 -44932
rect -61443 -45168 -61207 -44932
rect -61103 -45168 -60867 -44932
rect -60783 -45168 -60547 -44932
rect -60443 -45168 -60207 -44932
rect -60103 -45168 -59867 -44932
rect -59783 -45168 -59547 -44932
rect -59443 -45168 -59207 -44932
rect -59103 -45168 -58867 -44932
rect -58783 -45168 -58547 -44932
rect -58443 -45168 -58207 -44932
rect -58103 -45168 -57867 -44932
rect -57783 -45168 -57547 -44932
rect -57443 -45168 -57207 -44932
rect -57103 -45168 -56867 -44932
rect -56783 -45168 -56547 -44932
rect -56443 -45168 -56207 -44932
rect -56103 -45168 -55867 -44932
rect -55783 -45168 -55547 -44932
rect -55443 -45168 -55207 -44932
rect -55103 -45168 -54867 -44932
rect -54783 -45168 -54547 -44932
rect -54443 -45168 -54207 -44932
rect -54103 -45168 -53867 -44932
rect -53783 -45168 -53547 -44932
rect -53443 -45168 -53207 -44932
rect -53103 -45168 -52867 -44932
rect -52783 -45168 -52547 -44932
rect -52443 -45168 -52207 -44932
rect -52103 -45168 -51867 -44932
rect -51783 -45168 -51547 -44932
rect -51443 -45168 -51207 -44932
rect -51103 -45168 -50867 -44932
rect -50783 -45168 -50547 -44932
rect -50443 -45168 -50207 -44932
rect -50103 -45168 -49867 -44932
rect -49783 -45168 -49547 -44932
rect -49443 -45168 -49207 -44932
rect -49103 -45168 -48867 -44932
rect 8317 -45168 8553 -44932
rect 8657 -45168 8893 -44932
rect 8997 -45168 9233 -44932
rect 9317 -45168 9553 -44932
rect 9657 -45168 9893 -44932
rect 9997 -45168 10233 -44932
rect 10317 -45168 10553 -44932
rect 10657 -45168 10893 -44932
rect 10997 -45168 11233 -44932
rect 11317 -45168 11553 -44932
rect 11657 -45168 11893 -44932
rect 11997 -45168 12233 -44932
rect 12317 -45168 12553 -44932
rect 12657 -45168 12893 -44932
rect 12997 -45168 13233 -44932
rect 13317 -45168 13553 -44932
rect 13657 -45168 13893 -44932
rect 13997 -45168 14233 -44932
rect 14317 -45168 14553 -44932
rect 14657 -45168 14893 -44932
rect 14997 -45168 15233 -44932
rect 15317 -45168 15553 -44932
rect 15657 -45168 15893 -44932
rect 15997 -45168 16233 -44932
rect 16317 -45168 16553 -44932
rect 16657 -45168 16893 -44932
rect 16997 -45168 17233 -44932
rect 17317 -45168 17553 -44932
rect 17657 -45168 17893 -44932
rect 17997 -45168 18233 -44932
rect 18317 -45168 18553 -44932
rect 18657 -45168 18893 -44932
rect 18997 -45168 19233 -44932
rect 19317 -45168 19553 -44932
rect 19657 -45168 19893 -44932
rect 19997 -45168 20233 -44932
rect 20317 -45168 20553 -44932
rect 20657 -45168 20893 -44932
rect 20997 -45168 21233 -44932
rect 21317 -45168 21553 -44932
rect 21657 -45168 21893 -44932
rect 21997 -45168 22233 -44932
rect 22317 -45168 22553 -44932
rect 22657 -45168 22893 -44932
rect 22997 -45168 23233 -44932
rect 23317 -45168 23553 -44932
rect 23657 -45168 23893 -44932
rect 23997 -45168 24233 -44932
rect 24317 -45168 24553 -44932
rect 24657 -45168 24893 -44932
rect 24997 -45168 25233 -44932
rect 25317 -45168 25553 -44932
rect 25657 -45168 25893 -44932
rect 25997 -45168 26233 -44932
rect 26317 -45168 26553 -44932
rect 26657 -45168 26893 -44932
rect 26997 -45168 27233 -44932
rect 27317 -45168 27553 -44932
rect 27657 -45168 27893 -44932
rect 27997 -45168 28233 -44932
rect 28317 -45168 28553 -44932
rect 28657 -45168 28893 -44932
rect 28997 -45168 29233 -44932
rect 29317 -45168 29553 -44932
rect 29657 -45168 29893 -44932
rect 29997 -45168 30233 -44932
rect 30317 -45168 30553 -44932
rect 30657 -45168 30893 -44932
rect 30997 -45168 31233 -44932
rect 31317 -45168 31553 -44932
rect 31657 -45168 31893 -44932
rect 31997 -45168 32233 -44932
rect 32317 -45168 32553 -44932
rect 32657 -45168 32893 -44932
rect 32997 -45168 33233 -44932
rect 33317 -45168 33553 -44932
rect 33657 -45168 33893 -44932
rect 33997 -45168 34233 -44932
rect -74443 -45508 -74207 -45272
rect -74443 -45828 -74207 -45592
rect -73443 -45508 -73207 -45272
rect -73443 -45828 -73207 -45592
rect -72443 -45508 -72207 -45272
rect -72443 -45828 -72207 -45592
rect -71443 -45508 -71207 -45272
rect -71443 -45828 -71207 -45592
rect -70443 -45508 -70207 -45272
rect -70443 -45828 -70207 -45592
rect -69443 -45508 -69207 -45272
rect -69443 -45828 -69207 -45592
rect -68443 -45508 -68207 -45272
rect -68443 -45828 -68207 -45592
rect -67443 -45508 -67207 -45272
rect -67443 -45828 -67207 -45592
rect -66443 -45508 -66207 -45272
rect -66443 -45828 -66207 -45592
rect -65443 -45508 -65207 -45272
rect -65443 -45828 -65207 -45592
rect -64443 -45508 -64207 -45272
rect -64443 -45828 -64207 -45592
rect -63443 -45508 -63207 -45272
rect -63443 -45828 -63207 -45592
rect -62443 -45508 -62207 -45272
rect -62443 -45828 -62207 -45592
rect -61443 -45508 -61207 -45272
rect -61443 -45828 -61207 -45592
rect -60443 -45508 -60207 -45272
rect -60443 -45828 -60207 -45592
rect -59443 -45508 -59207 -45272
rect -59443 -45828 -59207 -45592
rect -58443 -45508 -58207 -45272
rect -58443 -45828 -58207 -45592
rect -57443 -45508 -57207 -45272
rect -57443 -45828 -57207 -45592
rect -56443 -45508 -56207 -45272
rect -56443 -45828 -56207 -45592
rect -55443 -45508 -55207 -45272
rect -55443 -45828 -55207 -45592
rect -54443 -45508 -54207 -45272
rect -54443 -45828 -54207 -45592
rect -53443 -45508 -53207 -45272
rect -53443 -45828 -53207 -45592
rect -52443 -45508 -52207 -45272
rect -52443 -45828 -52207 -45592
rect -51443 -45508 -51207 -45272
rect -51443 -45828 -51207 -45592
rect -50443 -45508 -50207 -45272
rect -50443 -45828 -50207 -45592
rect -49443 -45508 -49207 -45272
rect -49443 -45828 -49207 -45592
rect 8657 -45508 8893 -45272
rect 8657 -45828 8893 -45592
rect 9657 -45508 9893 -45272
rect 9657 -45828 9893 -45592
rect 10657 -45508 10893 -45272
rect 10657 -45828 10893 -45592
rect 11657 -45508 11893 -45272
rect 11657 -45828 11893 -45592
rect 12657 -45508 12893 -45272
rect 12657 -45828 12893 -45592
rect 13657 -45508 13893 -45272
rect 13657 -45828 13893 -45592
rect 14657 -45508 14893 -45272
rect 14657 -45828 14893 -45592
rect 15657 -45508 15893 -45272
rect 15657 -45828 15893 -45592
rect 16657 -45508 16893 -45272
rect 16657 -45828 16893 -45592
rect 17657 -45508 17893 -45272
rect 17657 -45828 17893 -45592
rect 18657 -45508 18893 -45272
rect 18657 -45828 18893 -45592
rect 19657 -45508 19893 -45272
rect 19657 -45828 19893 -45592
rect 20657 -45508 20893 -45272
rect 20657 -45828 20893 -45592
rect 21657 -45508 21893 -45272
rect 21657 -45828 21893 -45592
rect 22657 -45508 22893 -45272
rect 22657 -45828 22893 -45592
rect 23657 -45508 23893 -45272
rect 23657 -45828 23893 -45592
rect 24657 -45508 24893 -45272
rect 24657 -45828 24893 -45592
rect 25657 -45508 25893 -45272
rect 25657 -45828 25893 -45592
rect 26657 -45508 26893 -45272
rect 26657 -45828 26893 -45592
rect 27657 -45508 27893 -45272
rect 27657 -45828 27893 -45592
rect 28657 -45508 28893 -45272
rect 28657 -45828 28893 -45592
rect 29657 -45508 29893 -45272
rect 29657 -45828 29893 -45592
rect 30657 -45508 30893 -45272
rect 30657 -45828 30893 -45592
rect 31657 -45508 31893 -45272
rect 31657 -45828 31893 -45592
rect 32657 -45508 32893 -45272
rect 32657 -45828 32893 -45592
rect 33657 -45508 33893 -45272
rect 33657 -45828 33893 -45592
rect -74783 -46168 -74547 -45932
rect -74443 -46168 -74207 -45932
rect -74103 -46168 -73867 -45932
rect -73783 -46168 -73547 -45932
rect -73443 -46168 -73207 -45932
rect -73103 -46168 -72867 -45932
rect -72783 -46168 -72547 -45932
rect -72443 -46168 -72207 -45932
rect -72103 -46168 -71867 -45932
rect -71783 -46168 -71547 -45932
rect -71443 -46168 -71207 -45932
rect -71103 -46168 -70867 -45932
rect -70783 -46168 -70547 -45932
rect -70443 -46168 -70207 -45932
rect -70103 -46168 -69867 -45932
rect -69783 -46168 -69547 -45932
rect -69443 -46168 -69207 -45932
rect -69103 -46168 -68867 -45932
rect -68783 -46168 -68547 -45932
rect -68443 -46168 -68207 -45932
rect -68103 -46168 -67867 -45932
rect -67783 -46168 -67547 -45932
rect -67443 -46168 -67207 -45932
rect -67103 -46168 -66867 -45932
rect -66783 -46168 -66547 -45932
rect -66443 -46168 -66207 -45932
rect -66103 -46168 -65867 -45932
rect -65783 -46168 -65547 -45932
rect -65443 -46168 -65207 -45932
rect -65103 -46168 -64867 -45932
rect -64783 -46168 -64547 -45932
rect -64443 -46168 -64207 -45932
rect -64103 -46168 -63867 -45932
rect -63783 -46168 -63547 -45932
rect -63443 -46168 -63207 -45932
rect -63103 -46168 -62867 -45932
rect -62783 -46168 -62547 -45932
rect -62443 -46168 -62207 -45932
rect -62103 -46168 -61867 -45932
rect -61783 -46168 -61547 -45932
rect -61443 -46168 -61207 -45932
rect -61103 -46168 -60867 -45932
rect -60783 -46168 -60547 -45932
rect -60443 -46168 -60207 -45932
rect -60103 -46168 -59867 -45932
rect -59783 -46168 -59547 -45932
rect -59443 -46168 -59207 -45932
rect -59103 -46168 -58867 -45932
rect -58783 -46168 -58547 -45932
rect -58443 -46168 -58207 -45932
rect -58103 -46168 -57867 -45932
rect -57783 -46168 -57547 -45932
rect -57443 -46168 -57207 -45932
rect -57103 -46168 -56867 -45932
rect -56783 -46168 -56547 -45932
rect -56443 -46168 -56207 -45932
rect -56103 -46168 -55867 -45932
rect -55783 -46168 -55547 -45932
rect -55443 -46168 -55207 -45932
rect -55103 -46168 -54867 -45932
rect -54783 -46168 -54547 -45932
rect -54443 -46168 -54207 -45932
rect -54103 -46168 -53867 -45932
rect -53783 -46168 -53547 -45932
rect -53443 -46168 -53207 -45932
rect -53103 -46168 -52867 -45932
rect -52783 -46168 -52547 -45932
rect -52443 -46168 -52207 -45932
rect -52103 -46168 -51867 -45932
rect -51783 -46168 -51547 -45932
rect -51443 -46168 -51207 -45932
rect -51103 -46168 -50867 -45932
rect -50783 -46168 -50547 -45932
rect -50443 -46168 -50207 -45932
rect -50103 -46168 -49867 -45932
rect -49783 -46168 -49547 -45932
rect -49443 -46168 -49207 -45932
rect -49103 -46168 -48867 -45932
rect 8317 -46168 8553 -45932
rect 8657 -46168 8893 -45932
rect 8997 -46168 9233 -45932
rect 9317 -46168 9553 -45932
rect 9657 -46168 9893 -45932
rect 9997 -46168 10233 -45932
rect 10317 -46168 10553 -45932
rect 10657 -46168 10893 -45932
rect 10997 -46168 11233 -45932
rect 11317 -46168 11553 -45932
rect 11657 -46168 11893 -45932
rect 11997 -46168 12233 -45932
rect 12317 -46168 12553 -45932
rect 12657 -46168 12893 -45932
rect 12997 -46168 13233 -45932
rect 13317 -46168 13553 -45932
rect 13657 -46168 13893 -45932
rect 13997 -46168 14233 -45932
rect 14317 -46168 14553 -45932
rect 14657 -46168 14893 -45932
rect 14997 -46168 15233 -45932
rect 15317 -46168 15553 -45932
rect 15657 -46168 15893 -45932
rect 15997 -46168 16233 -45932
rect 16317 -46168 16553 -45932
rect 16657 -46168 16893 -45932
rect 16997 -46168 17233 -45932
rect 17317 -46168 17553 -45932
rect 17657 -46168 17893 -45932
rect 17997 -46168 18233 -45932
rect 18317 -46168 18553 -45932
rect 18657 -46168 18893 -45932
rect 18997 -46168 19233 -45932
rect 19317 -46168 19553 -45932
rect 19657 -46168 19893 -45932
rect 19997 -46168 20233 -45932
rect 20317 -46168 20553 -45932
rect 20657 -46168 20893 -45932
rect 20997 -46168 21233 -45932
rect 21317 -46168 21553 -45932
rect 21657 -46168 21893 -45932
rect 21997 -46168 22233 -45932
rect 22317 -46168 22553 -45932
rect 22657 -46168 22893 -45932
rect 22997 -46168 23233 -45932
rect 23317 -46168 23553 -45932
rect 23657 -46168 23893 -45932
rect 23997 -46168 24233 -45932
rect 24317 -46168 24553 -45932
rect 24657 -46168 24893 -45932
rect 24997 -46168 25233 -45932
rect 25317 -46168 25553 -45932
rect 25657 -46168 25893 -45932
rect 25997 -46168 26233 -45932
rect 26317 -46168 26553 -45932
rect 26657 -46168 26893 -45932
rect 26997 -46168 27233 -45932
rect 27317 -46168 27553 -45932
rect 27657 -46168 27893 -45932
rect 27997 -46168 28233 -45932
rect 28317 -46168 28553 -45932
rect 28657 -46168 28893 -45932
rect 28997 -46168 29233 -45932
rect 29317 -46168 29553 -45932
rect 29657 -46168 29893 -45932
rect 29997 -46168 30233 -45932
rect 30317 -46168 30553 -45932
rect 30657 -46168 30893 -45932
rect 30997 -46168 31233 -45932
rect 31317 -46168 31553 -45932
rect 31657 -46168 31893 -45932
rect 31997 -46168 32233 -45932
rect 32317 -46168 32553 -45932
rect 32657 -46168 32893 -45932
rect 32997 -46168 33233 -45932
rect 33317 -46168 33553 -45932
rect 33657 -46168 33893 -45932
rect 33997 -46168 34233 -45932
rect -74443 -46508 -74207 -46272
rect -73443 -46508 -73207 -46272
rect -72443 -46508 -72207 -46272
rect -71443 -46508 -71207 -46272
rect -70443 -46508 -70207 -46272
rect -69443 -46508 -69207 -46272
rect -68443 -46508 -68207 -46272
rect -67443 -46508 -67207 -46272
rect -66443 -46508 -66207 -46272
rect -65443 -46508 -65207 -46272
rect -64443 -46508 -64207 -46272
rect -63443 -46508 -63207 -46272
rect -62443 -46508 -62207 -46272
rect -61443 -46508 -61207 -46272
rect -60443 -46508 -60207 -46272
rect -59443 -46508 -59207 -46272
rect -58443 -46508 -58207 -46272
rect -57443 -46508 -57207 -46272
rect -56443 -46508 -56207 -46272
rect -55443 -46508 -55207 -46272
rect -54443 -46508 -54207 -46272
rect -53443 -46508 -53207 -46272
rect -52443 -46508 -52207 -46272
rect -51443 -46508 -51207 -46272
rect -50443 -46508 -50207 -46272
rect -49443 -46508 -49207 -46272
rect 8657 -46508 8893 -46272
rect 9657 -46508 9893 -46272
rect 10657 -46508 10893 -46272
rect 11657 -46508 11893 -46272
rect 12657 -46508 12893 -46272
rect 13657 -46508 13893 -46272
rect 14657 -46508 14893 -46272
rect 15657 -46508 15893 -46272
rect 16657 -46508 16893 -46272
rect 17657 -46508 17893 -46272
rect 18657 -46508 18893 -46272
rect 19657 -46508 19893 -46272
rect 20657 -46508 20893 -46272
rect 21657 -46508 21893 -46272
rect 22657 -46508 22893 -46272
rect 23657 -46508 23893 -46272
rect 24657 -46508 24893 -46272
rect 25657 -46508 25893 -46272
rect 26657 -46508 26893 -46272
rect 27657 -46508 27893 -46272
rect 28657 -46508 28893 -46272
rect 29657 -46508 29893 -46272
rect 30657 -46508 30893 -46272
rect 31657 -46508 31893 -46272
rect 32657 -46508 32893 -46272
rect 33657 -46508 33893 -46272
<< metal5 >>
rect -74485 38508 -74165 38550
rect -74485 38272 -74443 38508
rect -74207 38272 -74165 38508
rect -74485 38210 -74165 38272
rect -73485 38508 -73165 38550
rect -73485 38272 -73443 38508
rect -73207 38272 -73165 38508
rect -73485 38210 -73165 38272
rect -72485 38508 -72165 38550
rect -72485 38272 -72443 38508
rect -72207 38272 -72165 38508
rect -72485 38210 -72165 38272
rect -71485 38508 -71165 38550
rect -71485 38272 -71443 38508
rect -71207 38272 -71165 38508
rect -71485 38210 -71165 38272
rect -70485 38508 -70165 38550
rect -70485 38272 -70443 38508
rect -70207 38272 -70165 38508
rect -70485 38210 -70165 38272
rect -69485 38508 -69165 38550
rect -69485 38272 -69443 38508
rect -69207 38272 -69165 38508
rect -69485 38210 -69165 38272
rect -68485 38508 -68165 38550
rect -68485 38272 -68443 38508
rect -68207 38272 -68165 38508
rect -68485 38210 -68165 38272
rect -67485 38508 -67165 38550
rect -67485 38272 -67443 38508
rect -67207 38272 -67165 38508
rect -67485 38210 -67165 38272
rect -66485 38508 -66165 38550
rect -66485 38272 -66443 38508
rect -66207 38272 -66165 38508
rect -66485 38210 -66165 38272
rect -65485 38508 -65165 38550
rect -65485 38272 -65443 38508
rect -65207 38272 -65165 38508
rect -65485 38210 -65165 38272
rect -64485 38508 -64165 38550
rect -64485 38272 -64443 38508
rect -64207 38272 -64165 38508
rect -64485 38210 -64165 38272
rect -63485 38508 -63165 38550
rect -63485 38272 -63443 38508
rect -63207 38272 -63165 38508
rect -63485 38210 -63165 38272
rect -62485 38508 -62165 38550
rect -62485 38272 -62443 38508
rect -62207 38272 -62165 38508
rect -62485 38210 -62165 38272
rect -61485 38508 -61165 38550
rect -61485 38272 -61443 38508
rect -61207 38272 -61165 38508
rect -61485 38210 -61165 38272
rect -60485 38508 -60165 38550
rect -60485 38272 -60443 38508
rect -60207 38272 -60165 38508
rect -60485 38210 -60165 38272
rect -59485 38508 -59165 38550
rect -59485 38272 -59443 38508
rect -59207 38272 -59165 38508
rect -59485 38210 -59165 38272
rect 9994 38508 10314 38550
rect 9994 38272 10036 38508
rect 10272 38272 10314 38508
rect 9994 38210 10314 38272
rect 10994 38508 11314 38550
rect 10994 38272 11036 38508
rect 11272 38272 11314 38508
rect 10994 38210 11314 38272
rect 11994 38508 12314 38550
rect 11994 38272 12036 38508
rect 12272 38272 12314 38508
rect 11994 38210 12314 38272
rect 12994 38508 13314 38550
rect 12994 38272 13036 38508
rect 13272 38272 13314 38508
rect 12994 38210 13314 38272
rect 13994 38508 14314 38550
rect 13994 38272 14036 38508
rect 14272 38272 14314 38508
rect 13994 38210 14314 38272
rect 14994 38508 15314 38550
rect 14994 38272 15036 38508
rect 15272 38272 15314 38508
rect 14994 38210 15314 38272
rect 15994 38508 16314 38550
rect 15994 38272 16036 38508
rect 16272 38272 16314 38508
rect 15994 38210 16314 38272
rect 16994 38508 17314 38550
rect 16994 38272 17036 38508
rect 17272 38272 17314 38508
rect 16994 38210 17314 38272
rect 17994 38508 18314 38550
rect 17994 38272 18036 38508
rect 18272 38272 18314 38508
rect 17994 38210 18314 38272
rect 18994 38508 19314 38550
rect 18994 38272 19036 38508
rect 19272 38272 19314 38508
rect 18994 38210 19314 38272
rect 19994 38508 20314 38550
rect 19994 38272 20036 38508
rect 20272 38272 20314 38508
rect 19994 38210 20314 38272
rect 20994 38508 21314 38550
rect 20994 38272 21036 38508
rect 21272 38272 21314 38508
rect 20994 38210 21314 38272
rect 21994 38508 22314 38550
rect 21994 38272 22036 38508
rect 22272 38272 22314 38508
rect 21994 38210 22314 38272
rect 22994 38508 23314 38550
rect 22994 38272 23036 38508
rect 23272 38272 23314 38508
rect 22994 38210 23314 38272
rect 23994 38508 24314 38550
rect 23994 38272 24036 38508
rect 24272 38272 24314 38508
rect 23994 38210 24314 38272
rect 24994 38508 25314 38550
rect 24994 38272 25036 38508
rect 25272 38272 25314 38508
rect 24994 38210 25314 38272
rect 25994 38508 26314 38550
rect 25994 38272 26036 38508
rect 26272 38272 26314 38508
rect 25994 38210 26314 38272
rect 26994 38508 27314 38550
rect 26994 38272 27036 38508
rect 27272 38272 27314 38508
rect 26994 38210 27314 38272
rect 27994 38508 28314 38550
rect 27994 38272 28036 38508
rect 28272 38272 28314 38508
rect 27994 38210 28314 38272
rect 28994 38508 29314 38550
rect 28994 38272 29036 38508
rect 29272 38272 29314 38508
rect 28994 38210 29314 38272
rect 29994 38508 30314 38550
rect 29994 38272 30036 38508
rect 30272 38272 30314 38508
rect 29994 38210 30314 38272
rect 30994 38508 31314 38550
rect 30994 38272 31036 38508
rect 31272 38272 31314 38508
rect 30994 38210 31314 38272
rect 31994 38508 32314 38550
rect 31994 38272 32036 38508
rect 32272 38272 32314 38508
rect 31994 38210 32314 38272
rect 32994 38508 33314 38550
rect 32994 38272 33036 38508
rect 33272 38272 33314 38508
rect 32994 38210 33314 38272
rect 33994 38508 34314 38550
rect 33994 38272 34036 38508
rect 34272 38272 34314 38508
rect 33994 38210 34314 38272
rect -74825 38168 -58825 38210
rect -74825 37932 -74783 38168
rect -74547 37932 -74443 38168
rect -74207 37932 -74103 38168
rect -73867 37932 -73783 38168
rect -73547 37932 -73443 38168
rect -73207 37932 -73103 38168
rect -72867 37932 -72783 38168
rect -72547 37932 -72443 38168
rect -72207 37932 -72103 38168
rect -71867 37932 -71783 38168
rect -71547 37932 -71443 38168
rect -71207 37932 -71103 38168
rect -70867 37932 -70783 38168
rect -70547 37932 -70443 38168
rect -70207 37932 -70103 38168
rect -69867 37932 -69783 38168
rect -69547 37932 -69443 38168
rect -69207 37932 -69103 38168
rect -68867 37932 -68783 38168
rect -68547 37932 -68443 38168
rect -68207 37932 -68103 38168
rect -67867 37932 -67783 38168
rect -67547 37932 -67443 38168
rect -67207 37932 -67103 38168
rect -66867 37932 -66783 38168
rect -66547 37932 -66443 38168
rect -66207 37932 -66103 38168
rect -65867 37932 -65783 38168
rect -65547 37932 -65443 38168
rect -65207 37932 -65103 38168
rect -64867 37932 -64783 38168
rect -64547 37932 -64443 38168
rect -64207 37932 -64103 38168
rect -63867 37932 -63783 38168
rect -63547 37932 -63443 38168
rect -63207 37932 -63103 38168
rect -62867 37932 -62783 38168
rect -62547 37932 -62443 38168
rect -62207 37932 -62103 38168
rect -61867 37932 -61783 38168
rect -61547 37932 -61443 38168
rect -61207 37932 -61103 38168
rect -60867 37932 -60783 38168
rect -60547 37932 -60443 38168
rect -60207 37932 -60103 38168
rect -59867 37932 -59783 38168
rect -59547 37932 -59443 38168
rect -59207 37932 -59103 38168
rect -58867 37932 -58825 38168
rect -74825 37890 -58825 37932
rect 9654 38168 34654 38210
rect 9654 37932 9696 38168
rect 9932 37932 10036 38168
rect 10272 37932 10376 38168
rect 10612 37932 10696 38168
rect 10932 37932 11036 38168
rect 11272 37932 11376 38168
rect 11612 37932 11696 38168
rect 11932 37932 12036 38168
rect 12272 37932 12376 38168
rect 12612 37932 12696 38168
rect 12932 37932 13036 38168
rect 13272 37932 13376 38168
rect 13612 37932 13696 38168
rect 13932 37932 14036 38168
rect 14272 37932 14376 38168
rect 14612 37932 14696 38168
rect 14932 37932 15036 38168
rect 15272 37932 15376 38168
rect 15612 37932 15696 38168
rect 15932 37932 16036 38168
rect 16272 37932 16376 38168
rect 16612 37932 16696 38168
rect 16932 37932 17036 38168
rect 17272 37932 17376 38168
rect 17612 37932 17696 38168
rect 17932 37932 18036 38168
rect 18272 37932 18376 38168
rect 18612 37932 18696 38168
rect 18932 37932 19036 38168
rect 19272 37932 19376 38168
rect 19612 37932 19696 38168
rect 19932 37932 20036 38168
rect 20272 37932 20376 38168
rect 20612 37932 20696 38168
rect 20932 37932 21036 38168
rect 21272 37932 21376 38168
rect 21612 37932 21696 38168
rect 21932 37932 22036 38168
rect 22272 37932 22376 38168
rect 22612 37932 22696 38168
rect 22932 37932 23036 38168
rect 23272 37932 23376 38168
rect 23612 37932 23696 38168
rect 23932 37932 24036 38168
rect 24272 37932 24376 38168
rect 24612 37932 24696 38168
rect 24932 37932 25036 38168
rect 25272 37932 25376 38168
rect 25612 37932 25696 38168
rect 25932 37932 26036 38168
rect 26272 37932 26376 38168
rect 26612 37932 26696 38168
rect 26932 37932 27036 38168
rect 27272 37932 27376 38168
rect 27612 37932 27696 38168
rect 27932 37932 28036 38168
rect 28272 37932 28376 38168
rect 28612 37932 28696 38168
rect 28932 37932 29036 38168
rect 29272 37932 29376 38168
rect 29612 37932 29696 38168
rect 29932 37932 30036 38168
rect 30272 37932 30376 38168
rect 30612 37932 30696 38168
rect 30932 37932 31036 38168
rect 31272 37932 31376 38168
rect 31612 37932 31696 38168
rect 31932 37932 32036 38168
rect 32272 37932 32376 38168
rect 32612 37932 32696 38168
rect 32932 37932 33036 38168
rect 33272 37932 33376 38168
rect 33612 37932 33696 38168
rect 33932 37932 34036 38168
rect 34272 37932 34376 38168
rect 34612 37932 34654 38168
rect 9654 37890 34654 37932
rect -74485 37828 -74165 37890
rect -74485 37592 -74443 37828
rect -74207 37592 -74165 37828
rect -74485 37508 -74165 37592
rect -74485 37272 -74443 37508
rect -74207 37272 -74165 37508
rect -74485 37210 -74165 37272
rect -73485 37828 -73165 37890
rect -73485 37592 -73443 37828
rect -73207 37592 -73165 37828
rect -73485 37508 -73165 37592
rect -73485 37272 -73443 37508
rect -73207 37272 -73165 37508
rect -73485 37210 -73165 37272
rect -72485 37828 -72165 37890
rect -72485 37592 -72443 37828
rect -72207 37592 -72165 37828
rect -72485 37508 -72165 37592
rect -72485 37272 -72443 37508
rect -72207 37272 -72165 37508
rect -72485 37210 -72165 37272
rect -71485 37828 -71165 37890
rect -71485 37592 -71443 37828
rect -71207 37592 -71165 37828
rect -71485 37508 -71165 37592
rect -71485 37272 -71443 37508
rect -71207 37272 -71165 37508
rect -71485 37210 -71165 37272
rect -70485 37828 -70165 37890
rect -70485 37592 -70443 37828
rect -70207 37592 -70165 37828
rect -70485 37508 -70165 37592
rect -70485 37272 -70443 37508
rect -70207 37272 -70165 37508
rect -70485 37210 -70165 37272
rect -69485 37828 -69165 37890
rect -69485 37592 -69443 37828
rect -69207 37592 -69165 37828
rect -69485 37508 -69165 37592
rect -69485 37272 -69443 37508
rect -69207 37272 -69165 37508
rect -69485 37210 -69165 37272
rect -68485 37828 -68165 37890
rect -68485 37592 -68443 37828
rect -68207 37592 -68165 37828
rect -68485 37508 -68165 37592
rect -68485 37272 -68443 37508
rect -68207 37272 -68165 37508
rect -68485 37210 -68165 37272
rect -67485 37828 -67165 37890
rect -67485 37592 -67443 37828
rect -67207 37592 -67165 37828
rect -67485 37508 -67165 37592
rect -67485 37272 -67443 37508
rect -67207 37272 -67165 37508
rect -67485 37210 -67165 37272
rect -66485 37828 -66165 37890
rect -66485 37592 -66443 37828
rect -66207 37592 -66165 37828
rect -66485 37508 -66165 37592
rect -66485 37272 -66443 37508
rect -66207 37272 -66165 37508
rect -66485 37210 -66165 37272
rect -65485 37828 -65165 37890
rect -65485 37592 -65443 37828
rect -65207 37592 -65165 37828
rect -65485 37508 -65165 37592
rect -65485 37272 -65443 37508
rect -65207 37272 -65165 37508
rect -65485 37210 -65165 37272
rect -64485 37828 -64165 37890
rect -64485 37592 -64443 37828
rect -64207 37592 -64165 37828
rect -64485 37508 -64165 37592
rect -64485 37272 -64443 37508
rect -64207 37272 -64165 37508
rect -64485 37210 -64165 37272
rect -63485 37828 -63165 37890
rect -63485 37592 -63443 37828
rect -63207 37592 -63165 37828
rect -63485 37508 -63165 37592
rect -63485 37272 -63443 37508
rect -63207 37272 -63165 37508
rect -63485 37210 -63165 37272
rect -62485 37828 -62165 37890
rect -62485 37592 -62443 37828
rect -62207 37592 -62165 37828
rect -62485 37508 -62165 37592
rect -62485 37272 -62443 37508
rect -62207 37272 -62165 37508
rect -62485 37210 -62165 37272
rect -61485 37828 -61165 37890
rect -61485 37592 -61443 37828
rect -61207 37592 -61165 37828
rect -61485 37508 -61165 37592
rect -61485 37272 -61443 37508
rect -61207 37272 -61165 37508
rect -61485 37210 -61165 37272
rect -60485 37828 -60165 37890
rect -60485 37592 -60443 37828
rect -60207 37592 -60165 37828
rect -60485 37508 -60165 37592
rect -60485 37272 -60443 37508
rect -60207 37272 -60165 37508
rect -60485 37210 -60165 37272
rect -59485 37828 -59165 37890
rect -59485 37592 -59443 37828
rect -59207 37592 -59165 37828
rect -59485 37508 -59165 37592
rect -59485 37272 -59443 37508
rect -59207 37272 -59165 37508
rect -59485 37210 -59165 37272
rect 9994 37828 10314 37890
rect 9994 37592 10036 37828
rect 10272 37592 10314 37828
rect 9994 37508 10314 37592
rect 9994 37272 10036 37508
rect 10272 37272 10314 37508
rect 9994 37210 10314 37272
rect 10994 37828 11314 37890
rect 10994 37592 11036 37828
rect 11272 37592 11314 37828
rect 10994 37508 11314 37592
rect 10994 37272 11036 37508
rect 11272 37272 11314 37508
rect 10994 37210 11314 37272
rect 11994 37828 12314 37890
rect 11994 37592 12036 37828
rect 12272 37592 12314 37828
rect 11994 37508 12314 37592
rect 11994 37272 12036 37508
rect 12272 37272 12314 37508
rect 11994 37210 12314 37272
rect 12994 37828 13314 37890
rect 12994 37592 13036 37828
rect 13272 37592 13314 37828
rect 12994 37508 13314 37592
rect 12994 37272 13036 37508
rect 13272 37272 13314 37508
rect 12994 37210 13314 37272
rect 13994 37828 14314 37890
rect 13994 37592 14036 37828
rect 14272 37592 14314 37828
rect 13994 37508 14314 37592
rect 13994 37272 14036 37508
rect 14272 37272 14314 37508
rect 13994 37210 14314 37272
rect 14994 37828 15314 37890
rect 14994 37592 15036 37828
rect 15272 37592 15314 37828
rect 14994 37508 15314 37592
rect 14994 37272 15036 37508
rect 15272 37272 15314 37508
rect 14994 37210 15314 37272
rect 15994 37828 16314 37890
rect 15994 37592 16036 37828
rect 16272 37592 16314 37828
rect 15994 37508 16314 37592
rect 15994 37272 16036 37508
rect 16272 37272 16314 37508
rect 15994 37210 16314 37272
rect 16994 37828 17314 37890
rect 16994 37592 17036 37828
rect 17272 37592 17314 37828
rect 16994 37508 17314 37592
rect 16994 37272 17036 37508
rect 17272 37272 17314 37508
rect 16994 37210 17314 37272
rect 17994 37828 18314 37890
rect 17994 37592 18036 37828
rect 18272 37592 18314 37828
rect 17994 37508 18314 37592
rect 17994 37272 18036 37508
rect 18272 37272 18314 37508
rect 17994 37210 18314 37272
rect 18994 37828 19314 37890
rect 18994 37592 19036 37828
rect 19272 37592 19314 37828
rect 18994 37508 19314 37592
rect 18994 37272 19036 37508
rect 19272 37272 19314 37508
rect 18994 37210 19314 37272
rect 19994 37828 20314 37890
rect 19994 37592 20036 37828
rect 20272 37592 20314 37828
rect 19994 37508 20314 37592
rect 19994 37272 20036 37508
rect 20272 37272 20314 37508
rect 19994 37210 20314 37272
rect 20994 37828 21314 37890
rect 20994 37592 21036 37828
rect 21272 37592 21314 37828
rect 20994 37508 21314 37592
rect 20994 37272 21036 37508
rect 21272 37272 21314 37508
rect 20994 37210 21314 37272
rect 21994 37828 22314 37890
rect 21994 37592 22036 37828
rect 22272 37592 22314 37828
rect 21994 37508 22314 37592
rect 21994 37272 22036 37508
rect 22272 37272 22314 37508
rect 21994 37210 22314 37272
rect 22994 37828 23314 37890
rect 22994 37592 23036 37828
rect 23272 37592 23314 37828
rect 22994 37508 23314 37592
rect 22994 37272 23036 37508
rect 23272 37272 23314 37508
rect 22994 37210 23314 37272
rect 23994 37828 24314 37890
rect 23994 37592 24036 37828
rect 24272 37592 24314 37828
rect 23994 37508 24314 37592
rect 23994 37272 24036 37508
rect 24272 37272 24314 37508
rect 23994 37210 24314 37272
rect 24994 37828 25314 37890
rect 24994 37592 25036 37828
rect 25272 37592 25314 37828
rect 24994 37508 25314 37592
rect 24994 37272 25036 37508
rect 25272 37272 25314 37508
rect 24994 37210 25314 37272
rect 25994 37828 26314 37890
rect 25994 37592 26036 37828
rect 26272 37592 26314 37828
rect 25994 37508 26314 37592
rect 25994 37272 26036 37508
rect 26272 37272 26314 37508
rect 25994 37210 26314 37272
rect 26994 37828 27314 37890
rect 26994 37592 27036 37828
rect 27272 37592 27314 37828
rect 26994 37508 27314 37592
rect 26994 37272 27036 37508
rect 27272 37272 27314 37508
rect 26994 37210 27314 37272
rect 27994 37828 28314 37890
rect 27994 37592 28036 37828
rect 28272 37592 28314 37828
rect 27994 37508 28314 37592
rect 27994 37272 28036 37508
rect 28272 37272 28314 37508
rect 27994 37210 28314 37272
rect 28994 37828 29314 37890
rect 28994 37592 29036 37828
rect 29272 37592 29314 37828
rect 28994 37508 29314 37592
rect 28994 37272 29036 37508
rect 29272 37272 29314 37508
rect 28994 37210 29314 37272
rect 29994 37828 30314 37890
rect 29994 37592 30036 37828
rect 30272 37592 30314 37828
rect 29994 37508 30314 37592
rect 29994 37272 30036 37508
rect 30272 37272 30314 37508
rect 29994 37210 30314 37272
rect 30994 37828 31314 37890
rect 30994 37592 31036 37828
rect 31272 37592 31314 37828
rect 30994 37508 31314 37592
rect 30994 37272 31036 37508
rect 31272 37272 31314 37508
rect 30994 37210 31314 37272
rect 31994 37828 32314 37890
rect 31994 37592 32036 37828
rect 32272 37592 32314 37828
rect 31994 37508 32314 37592
rect 31994 37272 32036 37508
rect 32272 37272 32314 37508
rect 31994 37210 32314 37272
rect 32994 37828 33314 37890
rect 32994 37592 33036 37828
rect 33272 37592 33314 37828
rect 32994 37508 33314 37592
rect 32994 37272 33036 37508
rect 33272 37272 33314 37508
rect 32994 37210 33314 37272
rect 33994 37828 34314 37890
rect 33994 37592 34036 37828
rect 34272 37592 34314 37828
rect 33994 37508 34314 37592
rect 33994 37272 34036 37508
rect 34272 37272 34314 37508
rect 33994 37210 34314 37272
rect -74825 37168 -58825 37210
rect -74825 36932 -74783 37168
rect -74547 36932 -74443 37168
rect -74207 36932 -74103 37168
rect -73867 36932 -73783 37168
rect -73547 36932 -73443 37168
rect -73207 36932 -73103 37168
rect -72867 36932 -72783 37168
rect -72547 36932 -72443 37168
rect -72207 36932 -72103 37168
rect -71867 36932 -71783 37168
rect -71547 36932 -71443 37168
rect -71207 36932 -71103 37168
rect -70867 36932 -70783 37168
rect -70547 36932 -70443 37168
rect -70207 36932 -70103 37168
rect -69867 36932 -69783 37168
rect -69547 36932 -69443 37168
rect -69207 36932 -69103 37168
rect -68867 36932 -68783 37168
rect -68547 36932 -68443 37168
rect -68207 36932 -68103 37168
rect -67867 36932 -67783 37168
rect -67547 36932 -67443 37168
rect -67207 36932 -67103 37168
rect -66867 36932 -66783 37168
rect -66547 36932 -66443 37168
rect -66207 36932 -66103 37168
rect -65867 36932 -65783 37168
rect -65547 36932 -65443 37168
rect -65207 36932 -65103 37168
rect -64867 36932 -64783 37168
rect -64547 36932 -64443 37168
rect -64207 36932 -64103 37168
rect -63867 36932 -63783 37168
rect -63547 36932 -63443 37168
rect -63207 36932 -63103 37168
rect -62867 36932 -62783 37168
rect -62547 36932 -62443 37168
rect -62207 36932 -62103 37168
rect -61867 36932 -61783 37168
rect -61547 36932 -61443 37168
rect -61207 36932 -61103 37168
rect -60867 36932 -60783 37168
rect -60547 36932 -60443 37168
rect -60207 36932 -60103 37168
rect -59867 36932 -59783 37168
rect -59547 36932 -59443 37168
rect -59207 36932 -59103 37168
rect -58867 36932 -58825 37168
rect -74825 36890 -58825 36932
rect 9654 37168 34654 37210
rect 9654 36932 9696 37168
rect 9932 36932 10036 37168
rect 10272 36932 10376 37168
rect 10612 36932 10696 37168
rect 10932 36932 11036 37168
rect 11272 36932 11376 37168
rect 11612 36932 11696 37168
rect 11932 36932 12036 37168
rect 12272 36932 12376 37168
rect 12612 36932 12696 37168
rect 12932 36932 13036 37168
rect 13272 36932 13376 37168
rect 13612 36932 13696 37168
rect 13932 36932 14036 37168
rect 14272 36932 14376 37168
rect 14612 36932 14696 37168
rect 14932 36932 15036 37168
rect 15272 36932 15376 37168
rect 15612 36932 15696 37168
rect 15932 36932 16036 37168
rect 16272 36932 16376 37168
rect 16612 36932 16696 37168
rect 16932 36932 17036 37168
rect 17272 36932 17376 37168
rect 17612 36932 17696 37168
rect 17932 36932 18036 37168
rect 18272 36932 18376 37168
rect 18612 36932 18696 37168
rect 18932 36932 19036 37168
rect 19272 36932 19376 37168
rect 19612 36932 19696 37168
rect 19932 36932 20036 37168
rect 20272 36932 20376 37168
rect 20612 36932 20696 37168
rect 20932 36932 21036 37168
rect 21272 36932 21376 37168
rect 21612 36932 21696 37168
rect 21932 36932 22036 37168
rect 22272 36932 22376 37168
rect 22612 36932 22696 37168
rect 22932 36932 23036 37168
rect 23272 36932 23376 37168
rect 23612 36932 23696 37168
rect 23932 36932 24036 37168
rect 24272 36932 24376 37168
rect 24612 36932 24696 37168
rect 24932 36932 25036 37168
rect 25272 36932 25376 37168
rect 25612 36932 25696 37168
rect 25932 36932 26036 37168
rect 26272 36932 26376 37168
rect 26612 36932 26696 37168
rect 26932 36932 27036 37168
rect 27272 36932 27376 37168
rect 27612 36932 27696 37168
rect 27932 36932 28036 37168
rect 28272 36932 28376 37168
rect 28612 36932 28696 37168
rect 28932 36932 29036 37168
rect 29272 36932 29376 37168
rect 29612 36932 29696 37168
rect 29932 36932 30036 37168
rect 30272 36932 30376 37168
rect 30612 36932 30696 37168
rect 30932 36932 31036 37168
rect 31272 36932 31376 37168
rect 31612 36932 31696 37168
rect 31932 36932 32036 37168
rect 32272 36932 32376 37168
rect 32612 36932 32696 37168
rect 32932 36932 33036 37168
rect 33272 36932 33376 37168
rect 33612 36932 33696 37168
rect 33932 36932 34036 37168
rect 34272 36932 34376 37168
rect 34612 36932 34654 37168
rect 9654 36890 34654 36932
rect -74485 36828 -74165 36890
rect -74485 36592 -74443 36828
rect -74207 36592 -74165 36828
rect -74485 36508 -74165 36592
rect -74485 36272 -74443 36508
rect -74207 36272 -74165 36508
rect -74485 36210 -74165 36272
rect -73485 36828 -73165 36890
rect -73485 36592 -73443 36828
rect -73207 36592 -73165 36828
rect -73485 36508 -73165 36592
rect -73485 36272 -73443 36508
rect -73207 36272 -73165 36508
rect -73485 36210 -73165 36272
rect -72485 36828 -72165 36890
rect -72485 36592 -72443 36828
rect -72207 36592 -72165 36828
rect -72485 36508 -72165 36592
rect -72485 36272 -72443 36508
rect -72207 36272 -72165 36508
rect -72485 36210 -72165 36272
rect -71485 36828 -71165 36890
rect -71485 36592 -71443 36828
rect -71207 36592 -71165 36828
rect -71485 36508 -71165 36592
rect -71485 36272 -71443 36508
rect -71207 36272 -71165 36508
rect -71485 36210 -71165 36272
rect -70485 36828 -70165 36890
rect -70485 36592 -70443 36828
rect -70207 36592 -70165 36828
rect -70485 36508 -70165 36592
rect -70485 36272 -70443 36508
rect -70207 36272 -70165 36508
rect -70485 36210 -70165 36272
rect -69485 36828 -69165 36890
rect -69485 36592 -69443 36828
rect -69207 36592 -69165 36828
rect -69485 36508 -69165 36592
rect -69485 36272 -69443 36508
rect -69207 36272 -69165 36508
rect -69485 36210 -69165 36272
rect -68485 36828 -68165 36890
rect -68485 36592 -68443 36828
rect -68207 36592 -68165 36828
rect -68485 36508 -68165 36592
rect -68485 36272 -68443 36508
rect -68207 36272 -68165 36508
rect -68485 36210 -68165 36272
rect -67485 36828 -67165 36890
rect -67485 36592 -67443 36828
rect -67207 36592 -67165 36828
rect -67485 36508 -67165 36592
rect -67485 36272 -67443 36508
rect -67207 36272 -67165 36508
rect -67485 36210 -67165 36272
rect -66485 36828 -66165 36890
rect -66485 36592 -66443 36828
rect -66207 36592 -66165 36828
rect -66485 36508 -66165 36592
rect -66485 36272 -66443 36508
rect -66207 36272 -66165 36508
rect -66485 36210 -66165 36272
rect -65485 36828 -65165 36890
rect -65485 36592 -65443 36828
rect -65207 36592 -65165 36828
rect -65485 36508 -65165 36592
rect -65485 36272 -65443 36508
rect -65207 36272 -65165 36508
rect -65485 36210 -65165 36272
rect -64485 36828 -64165 36890
rect -64485 36592 -64443 36828
rect -64207 36592 -64165 36828
rect -64485 36508 -64165 36592
rect -64485 36272 -64443 36508
rect -64207 36272 -64165 36508
rect -64485 36210 -64165 36272
rect -63485 36828 -63165 36890
rect -63485 36592 -63443 36828
rect -63207 36592 -63165 36828
rect -63485 36508 -63165 36592
rect -63485 36272 -63443 36508
rect -63207 36272 -63165 36508
rect -63485 36210 -63165 36272
rect -62485 36828 -62165 36890
rect -62485 36592 -62443 36828
rect -62207 36592 -62165 36828
rect -62485 36508 -62165 36592
rect -62485 36272 -62443 36508
rect -62207 36272 -62165 36508
rect -62485 36210 -62165 36272
rect -61485 36828 -61165 36890
rect -61485 36592 -61443 36828
rect -61207 36592 -61165 36828
rect -61485 36508 -61165 36592
rect -61485 36272 -61443 36508
rect -61207 36272 -61165 36508
rect -61485 36210 -61165 36272
rect -60485 36828 -60165 36890
rect -60485 36592 -60443 36828
rect -60207 36592 -60165 36828
rect -60485 36508 -60165 36592
rect -60485 36272 -60443 36508
rect -60207 36272 -60165 36508
rect -60485 36210 -60165 36272
rect -59485 36828 -59165 36890
rect -59485 36592 -59443 36828
rect -59207 36592 -59165 36828
rect -59485 36508 -59165 36592
rect -59485 36272 -59443 36508
rect -59207 36272 -59165 36508
rect -59485 36210 -59165 36272
rect 9994 36828 10314 36890
rect 9994 36592 10036 36828
rect 10272 36592 10314 36828
rect 9994 36508 10314 36592
rect 9994 36272 10036 36508
rect 10272 36272 10314 36508
rect 9994 36210 10314 36272
rect 10994 36828 11314 36890
rect 10994 36592 11036 36828
rect 11272 36592 11314 36828
rect 10994 36508 11314 36592
rect 10994 36272 11036 36508
rect 11272 36272 11314 36508
rect 10994 36210 11314 36272
rect 11994 36828 12314 36890
rect 11994 36592 12036 36828
rect 12272 36592 12314 36828
rect 11994 36508 12314 36592
rect 11994 36272 12036 36508
rect 12272 36272 12314 36508
rect 11994 36210 12314 36272
rect 12994 36828 13314 36890
rect 12994 36592 13036 36828
rect 13272 36592 13314 36828
rect 12994 36508 13314 36592
rect 12994 36272 13036 36508
rect 13272 36272 13314 36508
rect 12994 36210 13314 36272
rect 13994 36828 14314 36890
rect 13994 36592 14036 36828
rect 14272 36592 14314 36828
rect 13994 36508 14314 36592
rect 13994 36272 14036 36508
rect 14272 36272 14314 36508
rect 13994 36210 14314 36272
rect 14994 36828 15314 36890
rect 14994 36592 15036 36828
rect 15272 36592 15314 36828
rect 14994 36508 15314 36592
rect 14994 36272 15036 36508
rect 15272 36272 15314 36508
rect 14994 36210 15314 36272
rect 15994 36828 16314 36890
rect 15994 36592 16036 36828
rect 16272 36592 16314 36828
rect 15994 36508 16314 36592
rect 15994 36272 16036 36508
rect 16272 36272 16314 36508
rect 15994 36210 16314 36272
rect 16994 36828 17314 36890
rect 16994 36592 17036 36828
rect 17272 36592 17314 36828
rect 16994 36508 17314 36592
rect 16994 36272 17036 36508
rect 17272 36272 17314 36508
rect 16994 36210 17314 36272
rect 17994 36828 18314 36890
rect 17994 36592 18036 36828
rect 18272 36592 18314 36828
rect 17994 36508 18314 36592
rect 17994 36272 18036 36508
rect 18272 36272 18314 36508
rect 17994 36210 18314 36272
rect 18994 36828 19314 36890
rect 18994 36592 19036 36828
rect 19272 36592 19314 36828
rect 18994 36508 19314 36592
rect 18994 36272 19036 36508
rect 19272 36272 19314 36508
rect 18994 36210 19314 36272
rect 19994 36828 20314 36890
rect 19994 36592 20036 36828
rect 20272 36592 20314 36828
rect 19994 36508 20314 36592
rect 19994 36272 20036 36508
rect 20272 36272 20314 36508
rect 19994 36210 20314 36272
rect 20994 36828 21314 36890
rect 20994 36592 21036 36828
rect 21272 36592 21314 36828
rect 20994 36508 21314 36592
rect 20994 36272 21036 36508
rect 21272 36272 21314 36508
rect 20994 36210 21314 36272
rect 21994 36828 22314 36890
rect 21994 36592 22036 36828
rect 22272 36592 22314 36828
rect 21994 36508 22314 36592
rect 21994 36272 22036 36508
rect 22272 36272 22314 36508
rect 21994 36210 22314 36272
rect 22994 36828 23314 36890
rect 22994 36592 23036 36828
rect 23272 36592 23314 36828
rect 22994 36508 23314 36592
rect 22994 36272 23036 36508
rect 23272 36272 23314 36508
rect 22994 36210 23314 36272
rect 23994 36828 24314 36890
rect 23994 36592 24036 36828
rect 24272 36592 24314 36828
rect 23994 36508 24314 36592
rect 23994 36272 24036 36508
rect 24272 36272 24314 36508
rect 23994 36210 24314 36272
rect 24994 36828 25314 36890
rect 24994 36592 25036 36828
rect 25272 36592 25314 36828
rect 24994 36508 25314 36592
rect 24994 36272 25036 36508
rect 25272 36272 25314 36508
rect 24994 36210 25314 36272
rect 25994 36828 26314 36890
rect 25994 36592 26036 36828
rect 26272 36592 26314 36828
rect 25994 36508 26314 36592
rect 25994 36272 26036 36508
rect 26272 36272 26314 36508
rect 25994 36210 26314 36272
rect 26994 36828 27314 36890
rect 26994 36592 27036 36828
rect 27272 36592 27314 36828
rect 26994 36508 27314 36592
rect 26994 36272 27036 36508
rect 27272 36272 27314 36508
rect 26994 36210 27314 36272
rect 27994 36828 28314 36890
rect 27994 36592 28036 36828
rect 28272 36592 28314 36828
rect 27994 36508 28314 36592
rect 27994 36272 28036 36508
rect 28272 36272 28314 36508
rect 27994 36210 28314 36272
rect 28994 36828 29314 36890
rect 28994 36592 29036 36828
rect 29272 36592 29314 36828
rect 28994 36508 29314 36592
rect 28994 36272 29036 36508
rect 29272 36272 29314 36508
rect 28994 36210 29314 36272
rect 29994 36828 30314 36890
rect 29994 36592 30036 36828
rect 30272 36592 30314 36828
rect 29994 36508 30314 36592
rect 29994 36272 30036 36508
rect 30272 36272 30314 36508
rect 29994 36210 30314 36272
rect 30994 36828 31314 36890
rect 30994 36592 31036 36828
rect 31272 36592 31314 36828
rect 30994 36508 31314 36592
rect 30994 36272 31036 36508
rect 31272 36272 31314 36508
rect 30994 36210 31314 36272
rect 31994 36828 32314 36890
rect 31994 36592 32036 36828
rect 32272 36592 32314 36828
rect 31994 36508 32314 36592
rect 31994 36272 32036 36508
rect 32272 36272 32314 36508
rect 31994 36210 32314 36272
rect 32994 36828 33314 36890
rect 32994 36592 33036 36828
rect 33272 36592 33314 36828
rect 32994 36508 33314 36592
rect 32994 36272 33036 36508
rect 33272 36272 33314 36508
rect 32994 36210 33314 36272
rect 33994 36828 34314 36890
rect 33994 36592 34036 36828
rect 34272 36592 34314 36828
rect 33994 36508 34314 36592
rect 33994 36272 34036 36508
rect 34272 36272 34314 36508
rect 33994 36210 34314 36272
rect -74825 36168 -58825 36210
rect -74825 35932 -74783 36168
rect -74547 35932 -74443 36168
rect -74207 35932 -74103 36168
rect -73867 35932 -73783 36168
rect -73547 35932 -73443 36168
rect -73207 35932 -73103 36168
rect -72867 35932 -72783 36168
rect -72547 35932 -72443 36168
rect -72207 35932 -72103 36168
rect -71867 35932 -71783 36168
rect -71547 35932 -71443 36168
rect -71207 35932 -71103 36168
rect -70867 35932 -70783 36168
rect -70547 35932 -70443 36168
rect -70207 35932 -70103 36168
rect -69867 35932 -69783 36168
rect -69547 35932 -69443 36168
rect -69207 35932 -69103 36168
rect -68867 35932 -68783 36168
rect -68547 35932 -68443 36168
rect -68207 35932 -68103 36168
rect -67867 35932 -67783 36168
rect -67547 35932 -67443 36168
rect -67207 35932 -67103 36168
rect -66867 35932 -66783 36168
rect -66547 35932 -66443 36168
rect -66207 35932 -66103 36168
rect -65867 35932 -65783 36168
rect -65547 35932 -65443 36168
rect -65207 35932 -65103 36168
rect -64867 35932 -64783 36168
rect -64547 35932 -64443 36168
rect -64207 35932 -64103 36168
rect -63867 35932 -63783 36168
rect -63547 35932 -63443 36168
rect -63207 35932 -63103 36168
rect -62867 35932 -62783 36168
rect -62547 35932 -62443 36168
rect -62207 35932 -62103 36168
rect -61867 35932 -61783 36168
rect -61547 35932 -61443 36168
rect -61207 35932 -61103 36168
rect -60867 35932 -60783 36168
rect -60547 35932 -60443 36168
rect -60207 35932 -60103 36168
rect -59867 35932 -59783 36168
rect -59547 35932 -59443 36168
rect -59207 35932 -59103 36168
rect -58867 35932 -58825 36168
rect -74825 35890 -58825 35932
rect 9654 36168 34654 36210
rect 9654 35932 9696 36168
rect 9932 35932 10036 36168
rect 10272 35932 10376 36168
rect 10612 35932 10696 36168
rect 10932 35932 11036 36168
rect 11272 35932 11376 36168
rect 11612 35932 11696 36168
rect 11932 35932 12036 36168
rect 12272 35932 12376 36168
rect 12612 35932 12696 36168
rect 12932 35932 13036 36168
rect 13272 35932 13376 36168
rect 13612 35932 13696 36168
rect 13932 35932 14036 36168
rect 14272 35932 14376 36168
rect 14612 35932 14696 36168
rect 14932 35932 15036 36168
rect 15272 35932 15376 36168
rect 15612 35932 15696 36168
rect 15932 35932 16036 36168
rect 16272 35932 16376 36168
rect 16612 35932 16696 36168
rect 16932 35932 17036 36168
rect 17272 35932 17376 36168
rect 17612 35932 17696 36168
rect 17932 35932 18036 36168
rect 18272 35932 18376 36168
rect 18612 35932 18696 36168
rect 18932 35932 19036 36168
rect 19272 35932 19376 36168
rect 19612 35932 19696 36168
rect 19932 35932 20036 36168
rect 20272 35932 20376 36168
rect 20612 35932 20696 36168
rect 20932 35932 21036 36168
rect 21272 35932 21376 36168
rect 21612 35932 21696 36168
rect 21932 35932 22036 36168
rect 22272 35932 22376 36168
rect 22612 35932 22696 36168
rect 22932 35932 23036 36168
rect 23272 35932 23376 36168
rect 23612 35932 23696 36168
rect 23932 35932 24036 36168
rect 24272 35932 24376 36168
rect 24612 35932 24696 36168
rect 24932 35932 25036 36168
rect 25272 35932 25376 36168
rect 25612 35932 25696 36168
rect 25932 35932 26036 36168
rect 26272 35932 26376 36168
rect 26612 35932 26696 36168
rect 26932 35932 27036 36168
rect 27272 35932 27376 36168
rect 27612 35932 27696 36168
rect 27932 35932 28036 36168
rect 28272 35932 28376 36168
rect 28612 35932 28696 36168
rect 28932 35932 29036 36168
rect 29272 35932 29376 36168
rect 29612 35932 29696 36168
rect 29932 35932 30036 36168
rect 30272 35932 30376 36168
rect 30612 35932 30696 36168
rect 30932 35932 31036 36168
rect 31272 35932 31376 36168
rect 31612 35932 31696 36168
rect 31932 35932 32036 36168
rect 32272 35932 32376 36168
rect 32612 35932 32696 36168
rect 32932 35932 33036 36168
rect 33272 35932 33376 36168
rect 33612 35932 33696 36168
rect 33932 35932 34036 36168
rect 34272 35932 34376 36168
rect 34612 35932 34654 36168
rect 9654 35890 34654 35932
rect -74485 35828 -74165 35890
rect -74485 35592 -74443 35828
rect -74207 35592 -74165 35828
rect -74485 35508 -74165 35592
rect -74485 35272 -74443 35508
rect -74207 35272 -74165 35508
rect -74485 35210 -74165 35272
rect -73485 35828 -73165 35890
rect -73485 35592 -73443 35828
rect -73207 35592 -73165 35828
rect -73485 35508 -73165 35592
rect -73485 35272 -73443 35508
rect -73207 35272 -73165 35508
rect -73485 35210 -73165 35272
rect -72485 35828 -72165 35890
rect -72485 35592 -72443 35828
rect -72207 35592 -72165 35828
rect -72485 35508 -72165 35592
rect -72485 35272 -72443 35508
rect -72207 35272 -72165 35508
rect -72485 35210 -72165 35272
rect -71485 35828 -71165 35890
rect -71485 35592 -71443 35828
rect -71207 35592 -71165 35828
rect -71485 35508 -71165 35592
rect -71485 35272 -71443 35508
rect -71207 35272 -71165 35508
rect -71485 35210 -71165 35272
rect -70485 35828 -70165 35890
rect -70485 35592 -70443 35828
rect -70207 35592 -70165 35828
rect -70485 35508 -70165 35592
rect -70485 35272 -70443 35508
rect -70207 35272 -70165 35508
rect -70485 35210 -70165 35272
rect -69485 35828 -69165 35890
rect -69485 35592 -69443 35828
rect -69207 35592 -69165 35828
rect -69485 35508 -69165 35592
rect -69485 35272 -69443 35508
rect -69207 35272 -69165 35508
rect -69485 35210 -69165 35272
rect -68485 35828 -68165 35890
rect -68485 35592 -68443 35828
rect -68207 35592 -68165 35828
rect -68485 35508 -68165 35592
rect -68485 35272 -68443 35508
rect -68207 35272 -68165 35508
rect -68485 35210 -68165 35272
rect -67485 35828 -67165 35890
rect -67485 35592 -67443 35828
rect -67207 35592 -67165 35828
rect -67485 35508 -67165 35592
rect -67485 35272 -67443 35508
rect -67207 35272 -67165 35508
rect -67485 35210 -67165 35272
rect -66485 35828 -66165 35890
rect -66485 35592 -66443 35828
rect -66207 35592 -66165 35828
rect -66485 35508 -66165 35592
rect -66485 35272 -66443 35508
rect -66207 35272 -66165 35508
rect -66485 35210 -66165 35272
rect -65485 35828 -65165 35890
rect -65485 35592 -65443 35828
rect -65207 35592 -65165 35828
rect -65485 35508 -65165 35592
rect -65485 35272 -65443 35508
rect -65207 35272 -65165 35508
rect -65485 35210 -65165 35272
rect -64485 35828 -64165 35890
rect -64485 35592 -64443 35828
rect -64207 35592 -64165 35828
rect -64485 35508 -64165 35592
rect -64485 35272 -64443 35508
rect -64207 35272 -64165 35508
rect -64485 35210 -64165 35272
rect -63485 35828 -63165 35890
rect -63485 35592 -63443 35828
rect -63207 35592 -63165 35828
rect -63485 35508 -63165 35592
rect -63485 35272 -63443 35508
rect -63207 35272 -63165 35508
rect -63485 35210 -63165 35272
rect -62485 35828 -62165 35890
rect -62485 35592 -62443 35828
rect -62207 35592 -62165 35828
rect -62485 35508 -62165 35592
rect -62485 35272 -62443 35508
rect -62207 35272 -62165 35508
rect -62485 35210 -62165 35272
rect -61485 35828 -61165 35890
rect -61485 35592 -61443 35828
rect -61207 35592 -61165 35828
rect -61485 35508 -61165 35592
rect -61485 35272 -61443 35508
rect -61207 35272 -61165 35508
rect -61485 35210 -61165 35272
rect -60485 35828 -60165 35890
rect -60485 35592 -60443 35828
rect -60207 35592 -60165 35828
rect -60485 35508 -60165 35592
rect -60485 35272 -60443 35508
rect -60207 35272 -60165 35508
rect -60485 35210 -60165 35272
rect -59485 35828 -59165 35890
rect -59485 35592 -59443 35828
rect -59207 35592 -59165 35828
rect -59485 35508 -59165 35592
rect -59485 35272 -59443 35508
rect -59207 35272 -59165 35508
rect -59485 35210 -59165 35272
rect 9994 35828 10314 35890
rect 9994 35592 10036 35828
rect 10272 35592 10314 35828
rect 9994 35508 10314 35592
rect 9994 35272 10036 35508
rect 10272 35272 10314 35508
rect 9994 35210 10314 35272
rect 10994 35828 11314 35890
rect 10994 35592 11036 35828
rect 11272 35592 11314 35828
rect 10994 35508 11314 35592
rect 10994 35272 11036 35508
rect 11272 35272 11314 35508
rect 10994 35210 11314 35272
rect 11994 35828 12314 35890
rect 11994 35592 12036 35828
rect 12272 35592 12314 35828
rect 11994 35508 12314 35592
rect 11994 35272 12036 35508
rect 12272 35272 12314 35508
rect 11994 35210 12314 35272
rect 12994 35828 13314 35890
rect 12994 35592 13036 35828
rect 13272 35592 13314 35828
rect 12994 35508 13314 35592
rect 12994 35272 13036 35508
rect 13272 35272 13314 35508
rect 12994 35210 13314 35272
rect 13994 35828 14314 35890
rect 13994 35592 14036 35828
rect 14272 35592 14314 35828
rect 13994 35508 14314 35592
rect 13994 35272 14036 35508
rect 14272 35272 14314 35508
rect 13994 35210 14314 35272
rect 14994 35828 15314 35890
rect 14994 35592 15036 35828
rect 15272 35592 15314 35828
rect 14994 35508 15314 35592
rect 14994 35272 15036 35508
rect 15272 35272 15314 35508
rect 14994 35210 15314 35272
rect 15994 35828 16314 35890
rect 15994 35592 16036 35828
rect 16272 35592 16314 35828
rect 15994 35508 16314 35592
rect 15994 35272 16036 35508
rect 16272 35272 16314 35508
rect 15994 35210 16314 35272
rect 16994 35828 17314 35890
rect 16994 35592 17036 35828
rect 17272 35592 17314 35828
rect 16994 35508 17314 35592
rect 16994 35272 17036 35508
rect 17272 35272 17314 35508
rect 16994 35210 17314 35272
rect 17994 35828 18314 35890
rect 17994 35592 18036 35828
rect 18272 35592 18314 35828
rect 17994 35508 18314 35592
rect 17994 35272 18036 35508
rect 18272 35272 18314 35508
rect 17994 35210 18314 35272
rect 18994 35828 19314 35890
rect 18994 35592 19036 35828
rect 19272 35592 19314 35828
rect 18994 35508 19314 35592
rect 18994 35272 19036 35508
rect 19272 35272 19314 35508
rect 18994 35210 19314 35272
rect 19994 35828 20314 35890
rect 19994 35592 20036 35828
rect 20272 35592 20314 35828
rect 19994 35508 20314 35592
rect 19994 35272 20036 35508
rect 20272 35272 20314 35508
rect 19994 35210 20314 35272
rect 20994 35828 21314 35890
rect 20994 35592 21036 35828
rect 21272 35592 21314 35828
rect 20994 35508 21314 35592
rect 20994 35272 21036 35508
rect 21272 35272 21314 35508
rect 20994 35210 21314 35272
rect 21994 35828 22314 35890
rect 21994 35592 22036 35828
rect 22272 35592 22314 35828
rect 21994 35508 22314 35592
rect 21994 35272 22036 35508
rect 22272 35272 22314 35508
rect 21994 35210 22314 35272
rect 22994 35828 23314 35890
rect 22994 35592 23036 35828
rect 23272 35592 23314 35828
rect 22994 35508 23314 35592
rect 22994 35272 23036 35508
rect 23272 35272 23314 35508
rect 22994 35210 23314 35272
rect 23994 35828 24314 35890
rect 23994 35592 24036 35828
rect 24272 35592 24314 35828
rect 23994 35508 24314 35592
rect 23994 35272 24036 35508
rect 24272 35272 24314 35508
rect 23994 35210 24314 35272
rect 24994 35828 25314 35890
rect 24994 35592 25036 35828
rect 25272 35592 25314 35828
rect 24994 35508 25314 35592
rect 24994 35272 25036 35508
rect 25272 35272 25314 35508
rect 24994 35210 25314 35272
rect 25994 35828 26314 35890
rect 25994 35592 26036 35828
rect 26272 35592 26314 35828
rect 25994 35508 26314 35592
rect 25994 35272 26036 35508
rect 26272 35272 26314 35508
rect 25994 35210 26314 35272
rect 26994 35828 27314 35890
rect 26994 35592 27036 35828
rect 27272 35592 27314 35828
rect 26994 35508 27314 35592
rect 26994 35272 27036 35508
rect 27272 35272 27314 35508
rect 26994 35210 27314 35272
rect 27994 35828 28314 35890
rect 27994 35592 28036 35828
rect 28272 35592 28314 35828
rect 27994 35508 28314 35592
rect 27994 35272 28036 35508
rect 28272 35272 28314 35508
rect 27994 35210 28314 35272
rect 28994 35828 29314 35890
rect 28994 35592 29036 35828
rect 29272 35592 29314 35828
rect 28994 35508 29314 35592
rect 28994 35272 29036 35508
rect 29272 35272 29314 35508
rect 28994 35210 29314 35272
rect 29994 35828 30314 35890
rect 29994 35592 30036 35828
rect 30272 35592 30314 35828
rect 29994 35508 30314 35592
rect 29994 35272 30036 35508
rect 30272 35272 30314 35508
rect 29994 35210 30314 35272
rect 30994 35828 31314 35890
rect 30994 35592 31036 35828
rect 31272 35592 31314 35828
rect 30994 35508 31314 35592
rect 30994 35272 31036 35508
rect 31272 35272 31314 35508
rect 30994 35210 31314 35272
rect 31994 35828 32314 35890
rect 31994 35592 32036 35828
rect 32272 35592 32314 35828
rect 31994 35508 32314 35592
rect 31994 35272 32036 35508
rect 32272 35272 32314 35508
rect 31994 35210 32314 35272
rect 32994 35828 33314 35890
rect 32994 35592 33036 35828
rect 33272 35592 33314 35828
rect 32994 35508 33314 35592
rect 32994 35272 33036 35508
rect 33272 35272 33314 35508
rect 32994 35210 33314 35272
rect 33994 35828 34314 35890
rect 33994 35592 34036 35828
rect 34272 35592 34314 35828
rect 33994 35508 34314 35592
rect 33994 35272 34036 35508
rect 34272 35272 34314 35508
rect 33994 35210 34314 35272
rect -74825 35168 -58825 35210
rect -74825 34932 -74783 35168
rect -74547 34932 -74443 35168
rect -74207 34932 -74103 35168
rect -73867 34932 -73783 35168
rect -73547 34932 -73443 35168
rect -73207 34932 -73103 35168
rect -72867 34932 -72783 35168
rect -72547 34932 -72443 35168
rect -72207 34932 -72103 35168
rect -71867 34932 -71783 35168
rect -71547 34932 -71443 35168
rect -71207 34932 -71103 35168
rect -70867 34932 -70783 35168
rect -70547 34932 -70443 35168
rect -70207 34932 -70103 35168
rect -69867 34932 -69783 35168
rect -69547 34932 -69443 35168
rect -69207 34932 -69103 35168
rect -68867 34932 -68783 35168
rect -68547 34932 -68443 35168
rect -68207 34932 -68103 35168
rect -67867 34932 -67783 35168
rect -67547 34932 -67443 35168
rect -67207 34932 -67103 35168
rect -66867 34932 -66783 35168
rect -66547 34932 -66443 35168
rect -66207 34932 -66103 35168
rect -65867 34932 -65783 35168
rect -65547 34932 -65443 35168
rect -65207 34932 -65103 35168
rect -64867 34932 -64783 35168
rect -64547 34932 -64443 35168
rect -64207 34932 -64103 35168
rect -63867 34932 -63783 35168
rect -63547 34932 -63443 35168
rect -63207 34932 -63103 35168
rect -62867 34932 -62783 35168
rect -62547 34932 -62443 35168
rect -62207 34932 -62103 35168
rect -61867 34932 -61783 35168
rect -61547 34932 -61443 35168
rect -61207 34932 -61103 35168
rect -60867 34932 -60783 35168
rect -60547 34932 -60443 35168
rect -60207 34932 -60103 35168
rect -59867 34932 -59783 35168
rect -59547 34932 -59443 35168
rect -59207 34932 -59103 35168
rect -58867 34932 -58825 35168
rect -74825 34890 -58825 34932
rect 9654 35168 34654 35210
rect 9654 34932 9696 35168
rect 9932 34932 10036 35168
rect 10272 34932 10376 35168
rect 10612 34932 10696 35168
rect 10932 34932 11036 35168
rect 11272 34932 11376 35168
rect 11612 34932 11696 35168
rect 11932 34932 12036 35168
rect 12272 34932 12376 35168
rect 12612 34932 12696 35168
rect 12932 34932 13036 35168
rect 13272 34932 13376 35168
rect 13612 34932 13696 35168
rect 13932 34932 14036 35168
rect 14272 34932 14376 35168
rect 14612 34932 14696 35168
rect 14932 34932 15036 35168
rect 15272 34932 15376 35168
rect 15612 34932 15696 35168
rect 15932 34932 16036 35168
rect 16272 34932 16376 35168
rect 16612 34932 16696 35168
rect 16932 34932 17036 35168
rect 17272 34932 17376 35168
rect 17612 34932 17696 35168
rect 17932 34932 18036 35168
rect 18272 34932 18376 35168
rect 18612 34932 18696 35168
rect 18932 34932 19036 35168
rect 19272 34932 19376 35168
rect 19612 34932 19696 35168
rect 19932 34932 20036 35168
rect 20272 34932 20376 35168
rect 20612 34932 20696 35168
rect 20932 34932 21036 35168
rect 21272 34932 21376 35168
rect 21612 34932 21696 35168
rect 21932 34932 22036 35168
rect 22272 34932 22376 35168
rect 22612 34932 22696 35168
rect 22932 34932 23036 35168
rect 23272 34932 23376 35168
rect 23612 34932 23696 35168
rect 23932 34932 24036 35168
rect 24272 34932 24376 35168
rect 24612 34932 24696 35168
rect 24932 34932 25036 35168
rect 25272 34932 25376 35168
rect 25612 34932 25696 35168
rect 25932 34932 26036 35168
rect 26272 34932 26376 35168
rect 26612 34932 26696 35168
rect 26932 34932 27036 35168
rect 27272 34932 27376 35168
rect 27612 34932 27696 35168
rect 27932 34932 28036 35168
rect 28272 34932 28376 35168
rect 28612 34932 28696 35168
rect 28932 34932 29036 35168
rect 29272 34932 29376 35168
rect 29612 34932 29696 35168
rect 29932 34932 30036 35168
rect 30272 34932 30376 35168
rect 30612 34932 30696 35168
rect 30932 34932 31036 35168
rect 31272 34932 31376 35168
rect 31612 34932 31696 35168
rect 31932 34932 32036 35168
rect 32272 34932 32376 35168
rect 32612 34932 32696 35168
rect 32932 34932 33036 35168
rect 33272 34932 33376 35168
rect 33612 34932 33696 35168
rect 33932 34932 34036 35168
rect 34272 34932 34376 35168
rect 34612 34932 34654 35168
rect 9654 34890 34654 34932
rect -74485 34828 -74165 34890
rect -74485 34592 -74443 34828
rect -74207 34592 -74165 34828
rect -74485 34508 -74165 34592
rect -74485 34272 -74443 34508
rect -74207 34272 -74165 34508
rect -74485 34210 -74165 34272
rect -73485 34828 -73165 34890
rect -73485 34592 -73443 34828
rect -73207 34592 -73165 34828
rect -73485 34508 -73165 34592
rect -73485 34272 -73443 34508
rect -73207 34272 -73165 34508
rect -73485 34210 -73165 34272
rect -72485 34828 -72165 34890
rect -72485 34592 -72443 34828
rect -72207 34592 -72165 34828
rect -72485 34508 -72165 34592
rect -72485 34272 -72443 34508
rect -72207 34272 -72165 34508
rect -72485 34210 -72165 34272
rect -71485 34828 -71165 34890
rect -71485 34592 -71443 34828
rect -71207 34592 -71165 34828
rect -71485 34508 -71165 34592
rect -71485 34272 -71443 34508
rect -71207 34272 -71165 34508
rect -71485 34210 -71165 34272
rect -70485 34828 -70165 34890
rect -70485 34592 -70443 34828
rect -70207 34592 -70165 34828
rect -70485 34508 -70165 34592
rect -70485 34272 -70443 34508
rect -70207 34272 -70165 34508
rect -70485 34210 -70165 34272
rect -69485 34828 -69165 34890
rect -69485 34592 -69443 34828
rect -69207 34592 -69165 34828
rect -69485 34508 -69165 34592
rect -69485 34272 -69443 34508
rect -69207 34272 -69165 34508
rect -69485 34210 -69165 34272
rect -68485 34828 -68165 34890
rect -68485 34592 -68443 34828
rect -68207 34592 -68165 34828
rect -68485 34508 -68165 34592
rect -68485 34272 -68443 34508
rect -68207 34272 -68165 34508
rect -68485 34210 -68165 34272
rect -67485 34828 -67165 34890
rect -67485 34592 -67443 34828
rect -67207 34592 -67165 34828
rect -67485 34508 -67165 34592
rect -67485 34272 -67443 34508
rect -67207 34272 -67165 34508
rect -67485 34210 -67165 34272
rect -66485 34828 -66165 34890
rect -66485 34592 -66443 34828
rect -66207 34592 -66165 34828
rect -66485 34508 -66165 34592
rect -66485 34272 -66443 34508
rect -66207 34272 -66165 34508
rect -66485 34210 -66165 34272
rect -65485 34828 -65165 34890
rect -65485 34592 -65443 34828
rect -65207 34592 -65165 34828
rect -65485 34508 -65165 34592
rect -65485 34272 -65443 34508
rect -65207 34272 -65165 34508
rect -65485 34210 -65165 34272
rect -64485 34828 -64165 34890
rect -64485 34592 -64443 34828
rect -64207 34592 -64165 34828
rect -64485 34508 -64165 34592
rect -64485 34272 -64443 34508
rect -64207 34272 -64165 34508
rect -64485 34210 -64165 34272
rect -63485 34828 -63165 34890
rect -63485 34592 -63443 34828
rect -63207 34592 -63165 34828
rect -63485 34508 -63165 34592
rect -63485 34272 -63443 34508
rect -63207 34272 -63165 34508
rect -63485 34210 -63165 34272
rect -62485 34828 -62165 34890
rect -62485 34592 -62443 34828
rect -62207 34592 -62165 34828
rect -62485 34508 -62165 34592
rect -62485 34272 -62443 34508
rect -62207 34272 -62165 34508
rect -62485 34210 -62165 34272
rect -61485 34828 -61165 34890
rect -61485 34592 -61443 34828
rect -61207 34592 -61165 34828
rect -61485 34508 -61165 34592
rect -61485 34272 -61443 34508
rect -61207 34272 -61165 34508
rect -61485 34210 -61165 34272
rect -60485 34828 -60165 34890
rect -60485 34592 -60443 34828
rect -60207 34592 -60165 34828
rect -60485 34508 -60165 34592
rect -60485 34272 -60443 34508
rect -60207 34272 -60165 34508
rect -60485 34210 -60165 34272
rect -59485 34828 -59165 34890
rect -59485 34592 -59443 34828
rect -59207 34592 -59165 34828
rect -59485 34508 -59165 34592
rect -59485 34272 -59443 34508
rect -59207 34272 -59165 34508
rect -59485 34210 -59165 34272
rect 9994 34828 10314 34890
rect 9994 34592 10036 34828
rect 10272 34592 10314 34828
rect 9994 34508 10314 34592
rect 9994 34272 10036 34508
rect 10272 34272 10314 34508
rect 9994 34210 10314 34272
rect 10994 34828 11314 34890
rect 10994 34592 11036 34828
rect 11272 34592 11314 34828
rect 10994 34508 11314 34592
rect 10994 34272 11036 34508
rect 11272 34272 11314 34508
rect 10994 34210 11314 34272
rect 11994 34828 12314 34890
rect 11994 34592 12036 34828
rect 12272 34592 12314 34828
rect 11994 34508 12314 34592
rect 11994 34272 12036 34508
rect 12272 34272 12314 34508
rect 11994 34210 12314 34272
rect 12994 34828 13314 34890
rect 12994 34592 13036 34828
rect 13272 34592 13314 34828
rect 12994 34508 13314 34592
rect 12994 34272 13036 34508
rect 13272 34272 13314 34508
rect 12994 34210 13314 34272
rect 13994 34828 14314 34890
rect 13994 34592 14036 34828
rect 14272 34592 14314 34828
rect 13994 34508 14314 34592
rect 13994 34272 14036 34508
rect 14272 34272 14314 34508
rect 13994 34210 14314 34272
rect 14994 34828 15314 34890
rect 14994 34592 15036 34828
rect 15272 34592 15314 34828
rect 14994 34508 15314 34592
rect 14994 34272 15036 34508
rect 15272 34272 15314 34508
rect 14994 34210 15314 34272
rect 15994 34828 16314 34890
rect 15994 34592 16036 34828
rect 16272 34592 16314 34828
rect 15994 34508 16314 34592
rect 15994 34272 16036 34508
rect 16272 34272 16314 34508
rect 15994 34210 16314 34272
rect 16994 34828 17314 34890
rect 16994 34592 17036 34828
rect 17272 34592 17314 34828
rect 16994 34508 17314 34592
rect 16994 34272 17036 34508
rect 17272 34272 17314 34508
rect 16994 34210 17314 34272
rect 17994 34828 18314 34890
rect 17994 34592 18036 34828
rect 18272 34592 18314 34828
rect 17994 34508 18314 34592
rect 17994 34272 18036 34508
rect 18272 34272 18314 34508
rect 17994 34210 18314 34272
rect 18994 34828 19314 34890
rect 18994 34592 19036 34828
rect 19272 34592 19314 34828
rect 18994 34508 19314 34592
rect 18994 34272 19036 34508
rect 19272 34272 19314 34508
rect 18994 34210 19314 34272
rect 19994 34828 20314 34890
rect 19994 34592 20036 34828
rect 20272 34592 20314 34828
rect 19994 34508 20314 34592
rect 19994 34272 20036 34508
rect 20272 34272 20314 34508
rect 19994 34210 20314 34272
rect 20994 34828 21314 34890
rect 20994 34592 21036 34828
rect 21272 34592 21314 34828
rect 20994 34508 21314 34592
rect 20994 34272 21036 34508
rect 21272 34272 21314 34508
rect 20994 34210 21314 34272
rect 21994 34828 22314 34890
rect 21994 34592 22036 34828
rect 22272 34592 22314 34828
rect 21994 34508 22314 34592
rect 21994 34272 22036 34508
rect 22272 34272 22314 34508
rect 21994 34210 22314 34272
rect 22994 34828 23314 34890
rect 22994 34592 23036 34828
rect 23272 34592 23314 34828
rect 22994 34508 23314 34592
rect 22994 34272 23036 34508
rect 23272 34272 23314 34508
rect 22994 34210 23314 34272
rect 23994 34828 24314 34890
rect 23994 34592 24036 34828
rect 24272 34592 24314 34828
rect 23994 34508 24314 34592
rect 23994 34272 24036 34508
rect 24272 34272 24314 34508
rect 23994 34210 24314 34272
rect 24994 34828 25314 34890
rect 24994 34592 25036 34828
rect 25272 34592 25314 34828
rect 24994 34508 25314 34592
rect 24994 34272 25036 34508
rect 25272 34272 25314 34508
rect 24994 34210 25314 34272
rect 25994 34828 26314 34890
rect 25994 34592 26036 34828
rect 26272 34592 26314 34828
rect 25994 34508 26314 34592
rect 25994 34272 26036 34508
rect 26272 34272 26314 34508
rect 25994 34210 26314 34272
rect 26994 34828 27314 34890
rect 26994 34592 27036 34828
rect 27272 34592 27314 34828
rect 26994 34508 27314 34592
rect 26994 34272 27036 34508
rect 27272 34272 27314 34508
rect 26994 34210 27314 34272
rect 27994 34828 28314 34890
rect 27994 34592 28036 34828
rect 28272 34592 28314 34828
rect 27994 34508 28314 34592
rect 27994 34272 28036 34508
rect 28272 34272 28314 34508
rect 27994 34210 28314 34272
rect 28994 34828 29314 34890
rect 28994 34592 29036 34828
rect 29272 34592 29314 34828
rect 28994 34508 29314 34592
rect 28994 34272 29036 34508
rect 29272 34272 29314 34508
rect 28994 34210 29314 34272
rect 29994 34828 30314 34890
rect 29994 34592 30036 34828
rect 30272 34592 30314 34828
rect 29994 34508 30314 34592
rect 29994 34272 30036 34508
rect 30272 34272 30314 34508
rect 29994 34210 30314 34272
rect 30994 34828 31314 34890
rect 30994 34592 31036 34828
rect 31272 34592 31314 34828
rect 30994 34508 31314 34592
rect 30994 34272 31036 34508
rect 31272 34272 31314 34508
rect 30994 34210 31314 34272
rect 31994 34828 32314 34890
rect 31994 34592 32036 34828
rect 32272 34592 32314 34828
rect 31994 34508 32314 34592
rect 31994 34272 32036 34508
rect 32272 34272 32314 34508
rect 31994 34210 32314 34272
rect 32994 34828 33314 34890
rect 32994 34592 33036 34828
rect 33272 34592 33314 34828
rect 32994 34508 33314 34592
rect 32994 34272 33036 34508
rect 33272 34272 33314 34508
rect 32994 34210 33314 34272
rect 33994 34828 34314 34890
rect 33994 34592 34036 34828
rect 34272 34592 34314 34828
rect 33994 34508 34314 34592
rect 33994 34272 34036 34508
rect 34272 34272 34314 34508
rect 33994 34210 34314 34272
rect -74825 34168 -58825 34210
rect -74825 33932 -74783 34168
rect -74547 33932 -74443 34168
rect -74207 33932 -74103 34168
rect -73867 33932 -73783 34168
rect -73547 33932 -73443 34168
rect -73207 33932 -73103 34168
rect -72867 33932 -72783 34168
rect -72547 33932 -72443 34168
rect -72207 33932 -72103 34168
rect -71867 33932 -71783 34168
rect -71547 33932 -71443 34168
rect -71207 33932 -71103 34168
rect -70867 33932 -70783 34168
rect -70547 33932 -70443 34168
rect -70207 33932 -70103 34168
rect -69867 33932 -69783 34168
rect -69547 33932 -69443 34168
rect -69207 33932 -69103 34168
rect -68867 33932 -68783 34168
rect -68547 33932 -68443 34168
rect -68207 33932 -68103 34168
rect -67867 33932 -67783 34168
rect -67547 33932 -67443 34168
rect -67207 33932 -67103 34168
rect -66867 33932 -66783 34168
rect -66547 33932 -66443 34168
rect -66207 33932 -66103 34168
rect -65867 33932 -65783 34168
rect -65547 33932 -65443 34168
rect -65207 33932 -65103 34168
rect -64867 33932 -64783 34168
rect -64547 33932 -64443 34168
rect -64207 33932 -64103 34168
rect -63867 33932 -63783 34168
rect -63547 33932 -63443 34168
rect -63207 33932 -63103 34168
rect -62867 33932 -62783 34168
rect -62547 33932 -62443 34168
rect -62207 33932 -62103 34168
rect -61867 33932 -61783 34168
rect -61547 33932 -61443 34168
rect -61207 33932 -61103 34168
rect -60867 33932 -60783 34168
rect -60547 33932 -60443 34168
rect -60207 33932 -60103 34168
rect -59867 33932 -59783 34168
rect -59547 33932 -59443 34168
rect -59207 33932 -59103 34168
rect -58867 33932 -58825 34168
rect -74825 33890 -58825 33932
rect 9654 34168 34654 34210
rect 9654 33932 9696 34168
rect 9932 33932 10036 34168
rect 10272 33932 10376 34168
rect 10612 33932 10696 34168
rect 10932 33932 11036 34168
rect 11272 33932 11376 34168
rect 11612 33932 11696 34168
rect 11932 33932 12036 34168
rect 12272 33932 12376 34168
rect 12612 33932 12696 34168
rect 12932 33932 13036 34168
rect 13272 33932 13376 34168
rect 13612 33932 13696 34168
rect 13932 33932 14036 34168
rect 14272 33932 14376 34168
rect 14612 33932 14696 34168
rect 14932 33932 15036 34168
rect 15272 33932 15376 34168
rect 15612 33932 15696 34168
rect 15932 33932 16036 34168
rect 16272 33932 16376 34168
rect 16612 33932 16696 34168
rect 16932 33932 17036 34168
rect 17272 33932 17376 34168
rect 17612 33932 17696 34168
rect 17932 33932 18036 34168
rect 18272 33932 18376 34168
rect 18612 33932 18696 34168
rect 18932 33932 19036 34168
rect 19272 33932 19376 34168
rect 19612 33932 19696 34168
rect 19932 33932 20036 34168
rect 20272 33932 20376 34168
rect 20612 33932 20696 34168
rect 20932 33932 21036 34168
rect 21272 33932 21376 34168
rect 21612 33932 21696 34168
rect 21932 33932 22036 34168
rect 22272 33932 22376 34168
rect 22612 33932 22696 34168
rect 22932 33932 23036 34168
rect 23272 33932 23376 34168
rect 23612 33932 23696 34168
rect 23932 33932 24036 34168
rect 24272 33932 24376 34168
rect 24612 33932 24696 34168
rect 24932 33932 25036 34168
rect 25272 33932 25376 34168
rect 25612 33932 25696 34168
rect 25932 33932 26036 34168
rect 26272 33932 26376 34168
rect 26612 33932 26696 34168
rect 26932 33932 27036 34168
rect 27272 33932 27376 34168
rect 27612 33932 27696 34168
rect 27932 33932 28036 34168
rect 28272 33932 28376 34168
rect 28612 33932 28696 34168
rect 28932 33932 29036 34168
rect 29272 33932 29376 34168
rect 29612 33932 29696 34168
rect 29932 33932 30036 34168
rect 30272 33932 30376 34168
rect 30612 33932 30696 34168
rect 30932 33932 31036 34168
rect 31272 33932 31376 34168
rect 31612 33932 31696 34168
rect 31932 33932 32036 34168
rect 32272 33932 32376 34168
rect 32612 33932 32696 34168
rect 32932 33932 33036 34168
rect 33272 33932 33376 34168
rect 33612 33932 33696 34168
rect 33932 33932 34036 34168
rect 34272 33932 34376 34168
rect 34612 33932 34654 34168
rect 9654 33890 34654 33932
rect -74485 33828 -74165 33890
rect -74485 33592 -74443 33828
rect -74207 33592 -74165 33828
rect -74485 33508 -74165 33592
rect -74485 33272 -74443 33508
rect -74207 33272 -74165 33508
rect -74485 33210 -74165 33272
rect -73485 33828 -73165 33890
rect -73485 33592 -73443 33828
rect -73207 33592 -73165 33828
rect -73485 33508 -73165 33592
rect -73485 33272 -73443 33508
rect -73207 33272 -73165 33508
rect -73485 33210 -73165 33272
rect -72485 33828 -72165 33890
rect -72485 33592 -72443 33828
rect -72207 33592 -72165 33828
rect -72485 33508 -72165 33592
rect -72485 33272 -72443 33508
rect -72207 33272 -72165 33508
rect -72485 33210 -72165 33272
rect -71485 33828 -71165 33890
rect -71485 33592 -71443 33828
rect -71207 33592 -71165 33828
rect -71485 33508 -71165 33592
rect -71485 33272 -71443 33508
rect -71207 33272 -71165 33508
rect -71485 33210 -71165 33272
rect -70485 33828 -70165 33890
rect -70485 33592 -70443 33828
rect -70207 33592 -70165 33828
rect -70485 33508 -70165 33592
rect -70485 33272 -70443 33508
rect -70207 33272 -70165 33508
rect -70485 33210 -70165 33272
rect -69485 33828 -69165 33890
rect -69485 33592 -69443 33828
rect -69207 33592 -69165 33828
rect -69485 33508 -69165 33592
rect -69485 33272 -69443 33508
rect -69207 33272 -69165 33508
rect -69485 33210 -69165 33272
rect -68485 33828 -68165 33890
rect -68485 33592 -68443 33828
rect -68207 33592 -68165 33828
rect -68485 33508 -68165 33592
rect -68485 33272 -68443 33508
rect -68207 33272 -68165 33508
rect -68485 33210 -68165 33272
rect -67485 33828 -67165 33890
rect -67485 33592 -67443 33828
rect -67207 33592 -67165 33828
rect -67485 33508 -67165 33592
rect -67485 33272 -67443 33508
rect -67207 33272 -67165 33508
rect -67485 33210 -67165 33272
rect -66485 33828 -66165 33890
rect -66485 33592 -66443 33828
rect -66207 33592 -66165 33828
rect -66485 33508 -66165 33592
rect -66485 33272 -66443 33508
rect -66207 33272 -66165 33508
rect -66485 33210 -66165 33272
rect -65485 33828 -65165 33890
rect -65485 33592 -65443 33828
rect -65207 33592 -65165 33828
rect -65485 33508 -65165 33592
rect -65485 33272 -65443 33508
rect -65207 33272 -65165 33508
rect -65485 33210 -65165 33272
rect -64485 33828 -64165 33890
rect -64485 33592 -64443 33828
rect -64207 33592 -64165 33828
rect -64485 33508 -64165 33592
rect -64485 33272 -64443 33508
rect -64207 33272 -64165 33508
rect -64485 33210 -64165 33272
rect -63485 33828 -63165 33890
rect -63485 33592 -63443 33828
rect -63207 33592 -63165 33828
rect -63485 33508 -63165 33592
rect -63485 33272 -63443 33508
rect -63207 33272 -63165 33508
rect -63485 33210 -63165 33272
rect -62485 33828 -62165 33890
rect -62485 33592 -62443 33828
rect -62207 33592 -62165 33828
rect -62485 33508 -62165 33592
rect -62485 33272 -62443 33508
rect -62207 33272 -62165 33508
rect -62485 33210 -62165 33272
rect -61485 33828 -61165 33890
rect -61485 33592 -61443 33828
rect -61207 33592 -61165 33828
rect -61485 33508 -61165 33592
rect -61485 33272 -61443 33508
rect -61207 33272 -61165 33508
rect -61485 33210 -61165 33272
rect -60485 33828 -60165 33890
rect -60485 33592 -60443 33828
rect -60207 33592 -60165 33828
rect -60485 33508 -60165 33592
rect -60485 33272 -60443 33508
rect -60207 33272 -60165 33508
rect -60485 33210 -60165 33272
rect -59485 33828 -59165 33890
rect -59485 33592 -59443 33828
rect -59207 33592 -59165 33828
rect -59485 33508 -59165 33592
rect -59485 33272 -59443 33508
rect -59207 33272 -59165 33508
rect -59485 33210 -59165 33272
rect 9994 33828 10314 33890
rect 9994 33592 10036 33828
rect 10272 33592 10314 33828
rect 9994 33508 10314 33592
rect 9994 33272 10036 33508
rect 10272 33272 10314 33508
rect 9994 33210 10314 33272
rect 10994 33828 11314 33890
rect 10994 33592 11036 33828
rect 11272 33592 11314 33828
rect 10994 33508 11314 33592
rect 10994 33272 11036 33508
rect 11272 33272 11314 33508
rect 10994 33210 11314 33272
rect 11994 33828 12314 33890
rect 11994 33592 12036 33828
rect 12272 33592 12314 33828
rect 11994 33508 12314 33592
rect 11994 33272 12036 33508
rect 12272 33272 12314 33508
rect 11994 33210 12314 33272
rect 12994 33828 13314 33890
rect 12994 33592 13036 33828
rect 13272 33592 13314 33828
rect 12994 33508 13314 33592
rect 12994 33272 13036 33508
rect 13272 33272 13314 33508
rect 12994 33210 13314 33272
rect 13994 33828 14314 33890
rect 13994 33592 14036 33828
rect 14272 33592 14314 33828
rect 13994 33508 14314 33592
rect 13994 33272 14036 33508
rect 14272 33272 14314 33508
rect 13994 33210 14314 33272
rect 14994 33828 15314 33890
rect 14994 33592 15036 33828
rect 15272 33592 15314 33828
rect 14994 33508 15314 33592
rect 14994 33272 15036 33508
rect 15272 33272 15314 33508
rect 14994 33210 15314 33272
rect 15994 33828 16314 33890
rect 15994 33592 16036 33828
rect 16272 33592 16314 33828
rect 15994 33508 16314 33592
rect 15994 33272 16036 33508
rect 16272 33272 16314 33508
rect 15994 33210 16314 33272
rect 16994 33828 17314 33890
rect 16994 33592 17036 33828
rect 17272 33592 17314 33828
rect 16994 33508 17314 33592
rect 16994 33272 17036 33508
rect 17272 33272 17314 33508
rect 16994 33210 17314 33272
rect 17994 33828 18314 33890
rect 17994 33592 18036 33828
rect 18272 33592 18314 33828
rect 17994 33508 18314 33592
rect 17994 33272 18036 33508
rect 18272 33272 18314 33508
rect 17994 33210 18314 33272
rect 18994 33828 19314 33890
rect 18994 33592 19036 33828
rect 19272 33592 19314 33828
rect 18994 33508 19314 33592
rect 18994 33272 19036 33508
rect 19272 33272 19314 33508
rect 18994 33210 19314 33272
rect 19994 33828 20314 33890
rect 19994 33592 20036 33828
rect 20272 33592 20314 33828
rect 19994 33508 20314 33592
rect 19994 33272 20036 33508
rect 20272 33272 20314 33508
rect 19994 33210 20314 33272
rect 20994 33828 21314 33890
rect 20994 33592 21036 33828
rect 21272 33592 21314 33828
rect 20994 33508 21314 33592
rect 20994 33272 21036 33508
rect 21272 33272 21314 33508
rect 20994 33210 21314 33272
rect 21994 33828 22314 33890
rect 21994 33592 22036 33828
rect 22272 33592 22314 33828
rect 21994 33508 22314 33592
rect 21994 33272 22036 33508
rect 22272 33272 22314 33508
rect 21994 33210 22314 33272
rect 22994 33828 23314 33890
rect 22994 33592 23036 33828
rect 23272 33592 23314 33828
rect 22994 33508 23314 33592
rect 22994 33272 23036 33508
rect 23272 33272 23314 33508
rect 22994 33210 23314 33272
rect 23994 33828 24314 33890
rect 23994 33592 24036 33828
rect 24272 33592 24314 33828
rect 23994 33508 24314 33592
rect 23994 33272 24036 33508
rect 24272 33272 24314 33508
rect 23994 33210 24314 33272
rect 24994 33828 25314 33890
rect 24994 33592 25036 33828
rect 25272 33592 25314 33828
rect 24994 33508 25314 33592
rect 24994 33272 25036 33508
rect 25272 33272 25314 33508
rect 24994 33210 25314 33272
rect 25994 33828 26314 33890
rect 25994 33592 26036 33828
rect 26272 33592 26314 33828
rect 25994 33508 26314 33592
rect 25994 33272 26036 33508
rect 26272 33272 26314 33508
rect 25994 33210 26314 33272
rect 26994 33828 27314 33890
rect 26994 33592 27036 33828
rect 27272 33592 27314 33828
rect 26994 33508 27314 33592
rect 26994 33272 27036 33508
rect 27272 33272 27314 33508
rect 26994 33210 27314 33272
rect 27994 33828 28314 33890
rect 27994 33592 28036 33828
rect 28272 33592 28314 33828
rect 27994 33508 28314 33592
rect 27994 33272 28036 33508
rect 28272 33272 28314 33508
rect 27994 33210 28314 33272
rect 28994 33828 29314 33890
rect 28994 33592 29036 33828
rect 29272 33592 29314 33828
rect 28994 33508 29314 33592
rect 28994 33272 29036 33508
rect 29272 33272 29314 33508
rect 28994 33210 29314 33272
rect 29994 33828 30314 33890
rect 29994 33592 30036 33828
rect 30272 33592 30314 33828
rect 29994 33508 30314 33592
rect 29994 33272 30036 33508
rect 30272 33272 30314 33508
rect 29994 33210 30314 33272
rect 30994 33828 31314 33890
rect 30994 33592 31036 33828
rect 31272 33592 31314 33828
rect 30994 33508 31314 33592
rect 30994 33272 31036 33508
rect 31272 33272 31314 33508
rect 30994 33210 31314 33272
rect 31994 33828 32314 33890
rect 31994 33592 32036 33828
rect 32272 33592 32314 33828
rect 31994 33508 32314 33592
rect 31994 33272 32036 33508
rect 32272 33272 32314 33508
rect 31994 33210 32314 33272
rect 32994 33828 33314 33890
rect 32994 33592 33036 33828
rect 33272 33592 33314 33828
rect 32994 33508 33314 33592
rect 32994 33272 33036 33508
rect 33272 33272 33314 33508
rect 32994 33210 33314 33272
rect 33994 33828 34314 33890
rect 33994 33592 34036 33828
rect 34272 33592 34314 33828
rect 33994 33508 34314 33592
rect 33994 33272 34036 33508
rect 34272 33272 34314 33508
rect 33994 33210 34314 33272
rect -74825 33168 -58825 33210
rect -74825 32932 -74783 33168
rect -74547 32932 -74443 33168
rect -74207 32932 -74103 33168
rect -73867 32932 -73783 33168
rect -73547 32932 -73443 33168
rect -73207 32932 -73103 33168
rect -72867 32932 -72783 33168
rect -72547 32932 -72443 33168
rect -72207 32932 -72103 33168
rect -71867 32932 -71783 33168
rect -71547 32932 -71443 33168
rect -71207 32932 -71103 33168
rect -70867 32932 -70783 33168
rect -70547 32932 -70443 33168
rect -70207 32932 -70103 33168
rect -69867 32932 -69783 33168
rect -69547 32932 -69443 33168
rect -69207 32932 -69103 33168
rect -68867 32932 -68783 33168
rect -68547 32932 -68443 33168
rect -68207 32932 -68103 33168
rect -67867 32932 -67783 33168
rect -67547 32932 -67443 33168
rect -67207 32932 -67103 33168
rect -66867 32932 -66783 33168
rect -66547 32932 -66443 33168
rect -66207 32932 -66103 33168
rect -65867 32932 -65783 33168
rect -65547 32932 -65443 33168
rect -65207 32932 -65103 33168
rect -64867 32932 -64783 33168
rect -64547 32932 -64443 33168
rect -64207 32932 -64103 33168
rect -63867 32932 -63783 33168
rect -63547 32932 -63443 33168
rect -63207 32932 -63103 33168
rect -62867 32932 -62783 33168
rect -62547 32932 -62443 33168
rect -62207 32932 -62103 33168
rect -61867 32932 -61783 33168
rect -61547 32932 -61443 33168
rect -61207 32932 -61103 33168
rect -60867 32932 -60783 33168
rect -60547 32932 -60443 33168
rect -60207 32932 -60103 33168
rect -59867 32932 -59783 33168
rect -59547 32932 -59443 33168
rect -59207 32932 -59103 33168
rect -58867 32932 -58825 33168
rect -74825 32890 -58825 32932
rect 9654 33168 34654 33210
rect 9654 32932 9696 33168
rect 9932 32932 10036 33168
rect 10272 32932 10376 33168
rect 10612 32932 10696 33168
rect 10932 32932 11036 33168
rect 11272 32932 11376 33168
rect 11612 32932 11696 33168
rect 11932 32932 12036 33168
rect 12272 32932 12376 33168
rect 12612 32932 12696 33168
rect 12932 32932 13036 33168
rect 13272 32932 13376 33168
rect 13612 32932 13696 33168
rect 13932 32932 14036 33168
rect 14272 32932 14376 33168
rect 14612 32932 14696 33168
rect 14932 32932 15036 33168
rect 15272 32932 15376 33168
rect 15612 32932 15696 33168
rect 15932 32932 16036 33168
rect 16272 32932 16376 33168
rect 16612 32932 16696 33168
rect 16932 32932 17036 33168
rect 17272 32932 17376 33168
rect 17612 32932 17696 33168
rect 17932 32932 18036 33168
rect 18272 32932 18376 33168
rect 18612 32932 18696 33168
rect 18932 32932 19036 33168
rect 19272 32932 19376 33168
rect 19612 32932 19696 33168
rect 19932 32932 20036 33168
rect 20272 32932 20376 33168
rect 20612 32932 20696 33168
rect 20932 32932 21036 33168
rect 21272 32932 21376 33168
rect 21612 32932 21696 33168
rect 21932 32932 22036 33168
rect 22272 32932 22376 33168
rect 22612 32932 22696 33168
rect 22932 32932 23036 33168
rect 23272 32932 23376 33168
rect 23612 32932 23696 33168
rect 23932 32932 24036 33168
rect 24272 32932 24376 33168
rect 24612 32932 24696 33168
rect 24932 32932 25036 33168
rect 25272 32932 25376 33168
rect 25612 32932 25696 33168
rect 25932 32932 26036 33168
rect 26272 32932 26376 33168
rect 26612 32932 26696 33168
rect 26932 32932 27036 33168
rect 27272 32932 27376 33168
rect 27612 32932 27696 33168
rect 27932 32932 28036 33168
rect 28272 32932 28376 33168
rect 28612 32932 28696 33168
rect 28932 32932 29036 33168
rect 29272 32932 29376 33168
rect 29612 32932 29696 33168
rect 29932 32932 30036 33168
rect 30272 32932 30376 33168
rect 30612 32932 30696 33168
rect 30932 32932 31036 33168
rect 31272 32932 31376 33168
rect 31612 32932 31696 33168
rect 31932 32932 32036 33168
rect 32272 32932 32376 33168
rect 32612 32932 32696 33168
rect 32932 32932 33036 33168
rect 33272 32932 33376 33168
rect 33612 32932 33696 33168
rect 33932 32932 34036 33168
rect 34272 32932 34376 33168
rect 34612 32932 34654 33168
rect 9654 32890 34654 32932
rect -74485 32828 -74165 32890
rect -74485 32592 -74443 32828
rect -74207 32592 -74165 32828
rect -74485 32508 -74165 32592
rect -74485 32272 -74443 32508
rect -74207 32272 -74165 32508
rect -74485 32210 -74165 32272
rect -73485 32828 -73165 32890
rect -73485 32592 -73443 32828
rect -73207 32592 -73165 32828
rect -73485 32508 -73165 32592
rect -73485 32272 -73443 32508
rect -73207 32272 -73165 32508
rect -73485 32210 -73165 32272
rect -72485 32828 -72165 32890
rect -72485 32592 -72443 32828
rect -72207 32592 -72165 32828
rect -72485 32508 -72165 32592
rect -72485 32272 -72443 32508
rect -72207 32272 -72165 32508
rect -72485 32210 -72165 32272
rect -71485 32828 -71165 32890
rect -71485 32592 -71443 32828
rect -71207 32592 -71165 32828
rect -71485 32508 -71165 32592
rect -71485 32272 -71443 32508
rect -71207 32272 -71165 32508
rect -71485 32210 -71165 32272
rect -70485 32828 -70165 32890
rect -70485 32592 -70443 32828
rect -70207 32592 -70165 32828
rect -70485 32508 -70165 32592
rect -70485 32272 -70443 32508
rect -70207 32272 -70165 32508
rect -70485 32210 -70165 32272
rect -69485 32828 -69165 32890
rect -69485 32592 -69443 32828
rect -69207 32592 -69165 32828
rect -69485 32508 -69165 32592
rect -69485 32272 -69443 32508
rect -69207 32272 -69165 32508
rect -69485 32210 -69165 32272
rect -68485 32828 -68165 32890
rect -68485 32592 -68443 32828
rect -68207 32592 -68165 32828
rect -68485 32508 -68165 32592
rect -68485 32272 -68443 32508
rect -68207 32272 -68165 32508
rect -68485 32210 -68165 32272
rect -67485 32828 -67165 32890
rect -67485 32592 -67443 32828
rect -67207 32592 -67165 32828
rect -67485 32508 -67165 32592
rect -67485 32272 -67443 32508
rect -67207 32272 -67165 32508
rect -67485 32210 -67165 32272
rect -66485 32828 -66165 32890
rect -66485 32592 -66443 32828
rect -66207 32592 -66165 32828
rect -66485 32508 -66165 32592
rect -66485 32272 -66443 32508
rect -66207 32272 -66165 32508
rect -66485 32210 -66165 32272
rect -65485 32828 -65165 32890
rect -65485 32592 -65443 32828
rect -65207 32592 -65165 32828
rect -65485 32508 -65165 32592
rect -65485 32272 -65443 32508
rect -65207 32272 -65165 32508
rect -65485 32210 -65165 32272
rect -64485 32828 -64165 32890
rect -64485 32592 -64443 32828
rect -64207 32592 -64165 32828
rect -64485 32508 -64165 32592
rect -64485 32272 -64443 32508
rect -64207 32272 -64165 32508
rect -64485 32210 -64165 32272
rect -63485 32828 -63165 32890
rect -63485 32592 -63443 32828
rect -63207 32592 -63165 32828
rect -63485 32508 -63165 32592
rect -63485 32272 -63443 32508
rect -63207 32272 -63165 32508
rect -63485 32210 -63165 32272
rect -62485 32828 -62165 32890
rect -62485 32592 -62443 32828
rect -62207 32592 -62165 32828
rect -62485 32508 -62165 32592
rect -62485 32272 -62443 32508
rect -62207 32272 -62165 32508
rect -62485 32210 -62165 32272
rect -61485 32828 -61165 32890
rect -61485 32592 -61443 32828
rect -61207 32592 -61165 32828
rect -61485 32508 -61165 32592
rect -61485 32272 -61443 32508
rect -61207 32272 -61165 32508
rect -61485 32210 -61165 32272
rect -60485 32828 -60165 32890
rect -60485 32592 -60443 32828
rect -60207 32592 -60165 32828
rect -60485 32508 -60165 32592
rect -60485 32272 -60443 32508
rect -60207 32272 -60165 32508
rect -60485 32210 -60165 32272
rect -59485 32828 -59165 32890
rect -59485 32592 -59443 32828
rect -59207 32592 -59165 32828
rect -59485 32508 -59165 32592
rect -59485 32272 -59443 32508
rect -59207 32272 -59165 32508
rect -59485 32210 -59165 32272
rect 9994 32828 10314 32890
rect 9994 32592 10036 32828
rect 10272 32592 10314 32828
rect 9994 32508 10314 32592
rect 9994 32272 10036 32508
rect 10272 32272 10314 32508
rect 9994 32210 10314 32272
rect 10994 32828 11314 32890
rect 10994 32592 11036 32828
rect 11272 32592 11314 32828
rect 10994 32508 11314 32592
rect 10994 32272 11036 32508
rect 11272 32272 11314 32508
rect 10994 32210 11314 32272
rect 11994 32828 12314 32890
rect 11994 32592 12036 32828
rect 12272 32592 12314 32828
rect 11994 32508 12314 32592
rect 11994 32272 12036 32508
rect 12272 32272 12314 32508
rect 11994 32210 12314 32272
rect 12994 32828 13314 32890
rect 12994 32592 13036 32828
rect 13272 32592 13314 32828
rect 12994 32508 13314 32592
rect 12994 32272 13036 32508
rect 13272 32272 13314 32508
rect 12994 32210 13314 32272
rect 13994 32828 14314 32890
rect 13994 32592 14036 32828
rect 14272 32592 14314 32828
rect 13994 32508 14314 32592
rect 13994 32272 14036 32508
rect 14272 32272 14314 32508
rect 13994 32210 14314 32272
rect 14994 32828 15314 32890
rect 14994 32592 15036 32828
rect 15272 32592 15314 32828
rect 14994 32508 15314 32592
rect 14994 32272 15036 32508
rect 15272 32272 15314 32508
rect 14994 32210 15314 32272
rect 15994 32828 16314 32890
rect 15994 32592 16036 32828
rect 16272 32592 16314 32828
rect 15994 32508 16314 32592
rect 15994 32272 16036 32508
rect 16272 32272 16314 32508
rect 15994 32210 16314 32272
rect 16994 32828 17314 32890
rect 16994 32592 17036 32828
rect 17272 32592 17314 32828
rect 16994 32508 17314 32592
rect 16994 32272 17036 32508
rect 17272 32272 17314 32508
rect 16994 32210 17314 32272
rect 17994 32828 18314 32890
rect 17994 32592 18036 32828
rect 18272 32592 18314 32828
rect 17994 32508 18314 32592
rect 17994 32272 18036 32508
rect 18272 32272 18314 32508
rect 17994 32210 18314 32272
rect 18994 32828 19314 32890
rect 18994 32592 19036 32828
rect 19272 32592 19314 32828
rect 18994 32508 19314 32592
rect 18994 32272 19036 32508
rect 19272 32272 19314 32508
rect 18994 32210 19314 32272
rect 19994 32828 20314 32890
rect 19994 32592 20036 32828
rect 20272 32592 20314 32828
rect 19994 32508 20314 32592
rect 19994 32272 20036 32508
rect 20272 32272 20314 32508
rect 19994 32210 20314 32272
rect 20994 32828 21314 32890
rect 20994 32592 21036 32828
rect 21272 32592 21314 32828
rect 20994 32508 21314 32592
rect 20994 32272 21036 32508
rect 21272 32272 21314 32508
rect 20994 32210 21314 32272
rect 21994 32828 22314 32890
rect 21994 32592 22036 32828
rect 22272 32592 22314 32828
rect 21994 32508 22314 32592
rect 21994 32272 22036 32508
rect 22272 32272 22314 32508
rect 21994 32210 22314 32272
rect 22994 32828 23314 32890
rect 22994 32592 23036 32828
rect 23272 32592 23314 32828
rect 22994 32508 23314 32592
rect 22994 32272 23036 32508
rect 23272 32272 23314 32508
rect 22994 32210 23314 32272
rect 23994 32828 24314 32890
rect 23994 32592 24036 32828
rect 24272 32592 24314 32828
rect 23994 32508 24314 32592
rect 23994 32272 24036 32508
rect 24272 32272 24314 32508
rect 23994 32210 24314 32272
rect 24994 32828 25314 32890
rect 24994 32592 25036 32828
rect 25272 32592 25314 32828
rect 24994 32508 25314 32592
rect 24994 32272 25036 32508
rect 25272 32272 25314 32508
rect 24994 32210 25314 32272
rect 25994 32828 26314 32890
rect 25994 32592 26036 32828
rect 26272 32592 26314 32828
rect 25994 32508 26314 32592
rect 25994 32272 26036 32508
rect 26272 32272 26314 32508
rect 25994 32210 26314 32272
rect 26994 32828 27314 32890
rect 26994 32592 27036 32828
rect 27272 32592 27314 32828
rect 26994 32508 27314 32592
rect 26994 32272 27036 32508
rect 27272 32272 27314 32508
rect 26994 32210 27314 32272
rect 27994 32828 28314 32890
rect 27994 32592 28036 32828
rect 28272 32592 28314 32828
rect 27994 32508 28314 32592
rect 27994 32272 28036 32508
rect 28272 32272 28314 32508
rect 27994 32210 28314 32272
rect 28994 32828 29314 32890
rect 28994 32592 29036 32828
rect 29272 32592 29314 32828
rect 28994 32508 29314 32592
rect 28994 32272 29036 32508
rect 29272 32272 29314 32508
rect 28994 32210 29314 32272
rect 29994 32828 30314 32890
rect 29994 32592 30036 32828
rect 30272 32592 30314 32828
rect 29994 32508 30314 32592
rect 29994 32272 30036 32508
rect 30272 32272 30314 32508
rect 29994 32210 30314 32272
rect 30994 32828 31314 32890
rect 30994 32592 31036 32828
rect 31272 32592 31314 32828
rect 30994 32508 31314 32592
rect 30994 32272 31036 32508
rect 31272 32272 31314 32508
rect 30994 32210 31314 32272
rect 31994 32828 32314 32890
rect 31994 32592 32036 32828
rect 32272 32592 32314 32828
rect 31994 32508 32314 32592
rect 31994 32272 32036 32508
rect 32272 32272 32314 32508
rect 31994 32210 32314 32272
rect 32994 32828 33314 32890
rect 32994 32592 33036 32828
rect 33272 32592 33314 32828
rect 32994 32508 33314 32592
rect 32994 32272 33036 32508
rect 33272 32272 33314 32508
rect 32994 32210 33314 32272
rect 33994 32828 34314 32890
rect 33994 32592 34036 32828
rect 34272 32592 34314 32828
rect 33994 32508 34314 32592
rect 33994 32272 34036 32508
rect 34272 32272 34314 32508
rect 33994 32210 34314 32272
rect -74825 32168 -58825 32210
rect -74825 31932 -74783 32168
rect -74547 31932 -74443 32168
rect -74207 31932 -74103 32168
rect -73867 31932 -73783 32168
rect -73547 31932 -73443 32168
rect -73207 31932 -73103 32168
rect -72867 31932 -72783 32168
rect -72547 31932 -72443 32168
rect -72207 31932 -72103 32168
rect -71867 31932 -71783 32168
rect -71547 31932 -71443 32168
rect -71207 31932 -71103 32168
rect -70867 31932 -70783 32168
rect -70547 31932 -70443 32168
rect -70207 31932 -70103 32168
rect -69867 31932 -69783 32168
rect -69547 31932 -69443 32168
rect -69207 31932 -69103 32168
rect -68867 31932 -68783 32168
rect -68547 31932 -68443 32168
rect -68207 31932 -68103 32168
rect -67867 31932 -67783 32168
rect -67547 31932 -67443 32168
rect -67207 31932 -67103 32168
rect -66867 31932 -66783 32168
rect -66547 31932 -66443 32168
rect -66207 31932 -66103 32168
rect -65867 31932 -65783 32168
rect -65547 31932 -65443 32168
rect -65207 31932 -65103 32168
rect -64867 31932 -64783 32168
rect -64547 31932 -64443 32168
rect -64207 31932 -64103 32168
rect -63867 31932 -63783 32168
rect -63547 31932 -63443 32168
rect -63207 31932 -63103 32168
rect -62867 31932 -62783 32168
rect -62547 31932 -62443 32168
rect -62207 31932 -62103 32168
rect -61867 31932 -61783 32168
rect -61547 31932 -61443 32168
rect -61207 31932 -61103 32168
rect -60867 31932 -60783 32168
rect -60547 31932 -60443 32168
rect -60207 31932 -60103 32168
rect -59867 31932 -59783 32168
rect -59547 31932 -59443 32168
rect -59207 31932 -59103 32168
rect -58867 31932 -58825 32168
rect -74825 31890 -58825 31932
rect 9654 32168 34654 32210
rect 9654 31932 9696 32168
rect 9932 31932 10036 32168
rect 10272 31932 10376 32168
rect 10612 31932 10696 32168
rect 10932 31932 11036 32168
rect 11272 31932 11376 32168
rect 11612 31932 11696 32168
rect 11932 31932 12036 32168
rect 12272 31932 12376 32168
rect 12612 31932 12696 32168
rect 12932 31932 13036 32168
rect 13272 31932 13376 32168
rect 13612 31932 13696 32168
rect 13932 31932 14036 32168
rect 14272 31932 14376 32168
rect 14612 31932 14696 32168
rect 14932 31932 15036 32168
rect 15272 31932 15376 32168
rect 15612 31932 15696 32168
rect 15932 31932 16036 32168
rect 16272 31932 16376 32168
rect 16612 31932 16696 32168
rect 16932 31932 17036 32168
rect 17272 31932 17376 32168
rect 17612 31932 17696 32168
rect 17932 31932 18036 32168
rect 18272 31932 18376 32168
rect 18612 31932 18696 32168
rect 18932 31932 19036 32168
rect 19272 31932 19376 32168
rect 19612 31932 19696 32168
rect 19932 31932 20036 32168
rect 20272 31932 20376 32168
rect 20612 31932 20696 32168
rect 20932 31932 21036 32168
rect 21272 31932 21376 32168
rect 21612 31932 21696 32168
rect 21932 31932 22036 32168
rect 22272 31932 22376 32168
rect 22612 31932 22696 32168
rect 22932 31932 23036 32168
rect 23272 31932 23376 32168
rect 23612 31932 23696 32168
rect 23932 31932 24036 32168
rect 24272 31932 24376 32168
rect 24612 31932 24696 32168
rect 24932 31932 25036 32168
rect 25272 31932 25376 32168
rect 25612 31932 25696 32168
rect 25932 31932 26036 32168
rect 26272 31932 26376 32168
rect 26612 31932 26696 32168
rect 26932 31932 27036 32168
rect 27272 31932 27376 32168
rect 27612 31932 27696 32168
rect 27932 31932 28036 32168
rect 28272 31932 28376 32168
rect 28612 31932 28696 32168
rect 28932 31932 29036 32168
rect 29272 31932 29376 32168
rect 29612 31932 29696 32168
rect 29932 31932 30036 32168
rect 30272 31932 30376 32168
rect 30612 31932 30696 32168
rect 30932 31932 31036 32168
rect 31272 31932 31376 32168
rect 31612 31932 31696 32168
rect 31932 31932 32036 32168
rect 32272 31932 32376 32168
rect 32612 31932 32696 32168
rect 32932 31932 33036 32168
rect 33272 31932 33376 32168
rect 33612 31932 33696 32168
rect 33932 31932 34036 32168
rect 34272 31932 34376 32168
rect 34612 31932 34654 32168
rect 9654 31890 34654 31932
rect -74485 31828 -74165 31890
rect -74485 31592 -74443 31828
rect -74207 31592 -74165 31828
rect -74485 31508 -74165 31592
rect -74485 31272 -74443 31508
rect -74207 31272 -74165 31508
rect -74485 31210 -74165 31272
rect -73485 31828 -73165 31890
rect -73485 31592 -73443 31828
rect -73207 31592 -73165 31828
rect -73485 31508 -73165 31592
rect -73485 31272 -73443 31508
rect -73207 31272 -73165 31508
rect -73485 31210 -73165 31272
rect -72485 31828 -72165 31890
rect -72485 31592 -72443 31828
rect -72207 31592 -72165 31828
rect -72485 31508 -72165 31592
rect -72485 31272 -72443 31508
rect -72207 31272 -72165 31508
rect -72485 31210 -72165 31272
rect -71485 31828 -71165 31890
rect -71485 31592 -71443 31828
rect -71207 31592 -71165 31828
rect -71485 31508 -71165 31592
rect -71485 31272 -71443 31508
rect -71207 31272 -71165 31508
rect -71485 31210 -71165 31272
rect -70485 31828 -70165 31890
rect -70485 31592 -70443 31828
rect -70207 31592 -70165 31828
rect -70485 31508 -70165 31592
rect -70485 31272 -70443 31508
rect -70207 31272 -70165 31508
rect -70485 31210 -70165 31272
rect -69485 31828 -69165 31890
rect -69485 31592 -69443 31828
rect -69207 31592 -69165 31828
rect -69485 31508 -69165 31592
rect -69485 31272 -69443 31508
rect -69207 31272 -69165 31508
rect -69485 31210 -69165 31272
rect -68485 31828 -68165 31890
rect -68485 31592 -68443 31828
rect -68207 31592 -68165 31828
rect -68485 31508 -68165 31592
rect -68485 31272 -68443 31508
rect -68207 31272 -68165 31508
rect -68485 31210 -68165 31272
rect -67485 31828 -67165 31890
rect -67485 31592 -67443 31828
rect -67207 31592 -67165 31828
rect -67485 31508 -67165 31592
rect -67485 31272 -67443 31508
rect -67207 31272 -67165 31508
rect -67485 31210 -67165 31272
rect -66485 31828 -66165 31890
rect -66485 31592 -66443 31828
rect -66207 31592 -66165 31828
rect -66485 31508 -66165 31592
rect -66485 31272 -66443 31508
rect -66207 31272 -66165 31508
rect -66485 31210 -66165 31272
rect -65485 31828 -65165 31890
rect -65485 31592 -65443 31828
rect -65207 31592 -65165 31828
rect -65485 31508 -65165 31592
rect -65485 31272 -65443 31508
rect -65207 31272 -65165 31508
rect -65485 31210 -65165 31272
rect -64485 31828 -64165 31890
rect -64485 31592 -64443 31828
rect -64207 31592 -64165 31828
rect -64485 31508 -64165 31592
rect -64485 31272 -64443 31508
rect -64207 31272 -64165 31508
rect -64485 31210 -64165 31272
rect -63485 31828 -63165 31890
rect -63485 31592 -63443 31828
rect -63207 31592 -63165 31828
rect -63485 31508 -63165 31592
rect -63485 31272 -63443 31508
rect -63207 31272 -63165 31508
rect -63485 31210 -63165 31272
rect -62485 31828 -62165 31890
rect -62485 31592 -62443 31828
rect -62207 31592 -62165 31828
rect -62485 31508 -62165 31592
rect -62485 31272 -62443 31508
rect -62207 31272 -62165 31508
rect -62485 31210 -62165 31272
rect -61485 31828 -61165 31890
rect -61485 31592 -61443 31828
rect -61207 31592 -61165 31828
rect -61485 31508 -61165 31592
rect -61485 31272 -61443 31508
rect -61207 31272 -61165 31508
rect -61485 31210 -61165 31272
rect -60485 31828 -60165 31890
rect -60485 31592 -60443 31828
rect -60207 31592 -60165 31828
rect -60485 31508 -60165 31592
rect -60485 31272 -60443 31508
rect -60207 31272 -60165 31508
rect -60485 31210 -60165 31272
rect -59485 31828 -59165 31890
rect -59485 31592 -59443 31828
rect -59207 31592 -59165 31828
rect -59485 31508 -59165 31592
rect -59485 31272 -59443 31508
rect -59207 31272 -59165 31508
rect -59485 31210 -59165 31272
rect 9994 31828 10314 31890
rect 9994 31592 10036 31828
rect 10272 31592 10314 31828
rect 9994 31508 10314 31592
rect 9994 31272 10036 31508
rect 10272 31272 10314 31508
rect 9994 31210 10314 31272
rect 10994 31828 11314 31890
rect 10994 31592 11036 31828
rect 11272 31592 11314 31828
rect 10994 31508 11314 31592
rect 10994 31272 11036 31508
rect 11272 31272 11314 31508
rect 10994 31210 11314 31272
rect 11994 31828 12314 31890
rect 11994 31592 12036 31828
rect 12272 31592 12314 31828
rect 11994 31508 12314 31592
rect 11994 31272 12036 31508
rect 12272 31272 12314 31508
rect 11994 31210 12314 31272
rect 12994 31828 13314 31890
rect 12994 31592 13036 31828
rect 13272 31592 13314 31828
rect 12994 31508 13314 31592
rect 12994 31272 13036 31508
rect 13272 31272 13314 31508
rect 12994 31210 13314 31272
rect 13994 31828 14314 31890
rect 13994 31592 14036 31828
rect 14272 31592 14314 31828
rect 13994 31508 14314 31592
rect 13994 31272 14036 31508
rect 14272 31272 14314 31508
rect 13994 31210 14314 31272
rect 14994 31828 15314 31890
rect 14994 31592 15036 31828
rect 15272 31592 15314 31828
rect 14994 31508 15314 31592
rect 14994 31272 15036 31508
rect 15272 31272 15314 31508
rect 14994 31210 15314 31272
rect 15994 31828 16314 31890
rect 15994 31592 16036 31828
rect 16272 31592 16314 31828
rect 15994 31508 16314 31592
rect 15994 31272 16036 31508
rect 16272 31272 16314 31508
rect 15994 31210 16314 31272
rect 16994 31828 17314 31890
rect 16994 31592 17036 31828
rect 17272 31592 17314 31828
rect 16994 31508 17314 31592
rect 16994 31272 17036 31508
rect 17272 31272 17314 31508
rect 16994 31210 17314 31272
rect 17994 31828 18314 31890
rect 17994 31592 18036 31828
rect 18272 31592 18314 31828
rect 17994 31508 18314 31592
rect 17994 31272 18036 31508
rect 18272 31272 18314 31508
rect 17994 31210 18314 31272
rect 18994 31828 19314 31890
rect 18994 31592 19036 31828
rect 19272 31592 19314 31828
rect 18994 31508 19314 31592
rect 18994 31272 19036 31508
rect 19272 31272 19314 31508
rect 18994 31210 19314 31272
rect 19994 31828 20314 31890
rect 19994 31592 20036 31828
rect 20272 31592 20314 31828
rect 19994 31508 20314 31592
rect 19994 31272 20036 31508
rect 20272 31272 20314 31508
rect 19994 31210 20314 31272
rect 20994 31828 21314 31890
rect 20994 31592 21036 31828
rect 21272 31592 21314 31828
rect 20994 31508 21314 31592
rect 20994 31272 21036 31508
rect 21272 31272 21314 31508
rect 20994 31210 21314 31272
rect 21994 31828 22314 31890
rect 21994 31592 22036 31828
rect 22272 31592 22314 31828
rect 21994 31508 22314 31592
rect 21994 31272 22036 31508
rect 22272 31272 22314 31508
rect 21994 31210 22314 31272
rect 22994 31828 23314 31890
rect 22994 31592 23036 31828
rect 23272 31592 23314 31828
rect 22994 31508 23314 31592
rect 22994 31272 23036 31508
rect 23272 31272 23314 31508
rect 22994 31210 23314 31272
rect 23994 31828 24314 31890
rect 23994 31592 24036 31828
rect 24272 31592 24314 31828
rect 23994 31508 24314 31592
rect 23994 31272 24036 31508
rect 24272 31272 24314 31508
rect 23994 31210 24314 31272
rect 24994 31828 25314 31890
rect 24994 31592 25036 31828
rect 25272 31592 25314 31828
rect 24994 31508 25314 31592
rect 24994 31272 25036 31508
rect 25272 31272 25314 31508
rect 24994 31210 25314 31272
rect 25994 31828 26314 31890
rect 25994 31592 26036 31828
rect 26272 31592 26314 31828
rect 25994 31508 26314 31592
rect 25994 31272 26036 31508
rect 26272 31272 26314 31508
rect 25994 31210 26314 31272
rect 26994 31828 27314 31890
rect 26994 31592 27036 31828
rect 27272 31592 27314 31828
rect 26994 31508 27314 31592
rect 26994 31272 27036 31508
rect 27272 31272 27314 31508
rect 26994 31210 27314 31272
rect 27994 31828 28314 31890
rect 27994 31592 28036 31828
rect 28272 31592 28314 31828
rect 27994 31508 28314 31592
rect 27994 31272 28036 31508
rect 28272 31272 28314 31508
rect 27994 31210 28314 31272
rect 28994 31828 29314 31890
rect 28994 31592 29036 31828
rect 29272 31592 29314 31828
rect 28994 31508 29314 31592
rect 28994 31272 29036 31508
rect 29272 31272 29314 31508
rect 28994 31210 29314 31272
rect 29994 31828 30314 31890
rect 29994 31592 30036 31828
rect 30272 31592 30314 31828
rect 29994 31508 30314 31592
rect 29994 31272 30036 31508
rect 30272 31272 30314 31508
rect 29994 31210 30314 31272
rect 30994 31828 31314 31890
rect 30994 31592 31036 31828
rect 31272 31592 31314 31828
rect 30994 31508 31314 31592
rect 30994 31272 31036 31508
rect 31272 31272 31314 31508
rect 30994 31210 31314 31272
rect 31994 31828 32314 31890
rect 31994 31592 32036 31828
rect 32272 31592 32314 31828
rect 31994 31508 32314 31592
rect 31994 31272 32036 31508
rect 32272 31272 32314 31508
rect 31994 31210 32314 31272
rect 32994 31828 33314 31890
rect 32994 31592 33036 31828
rect 33272 31592 33314 31828
rect 32994 31508 33314 31592
rect 32994 31272 33036 31508
rect 33272 31272 33314 31508
rect 32994 31210 33314 31272
rect 33994 31828 34314 31890
rect 33994 31592 34036 31828
rect 34272 31592 34314 31828
rect 33994 31508 34314 31592
rect 33994 31272 34036 31508
rect 34272 31272 34314 31508
rect 33994 31210 34314 31272
rect -74825 31168 -58825 31210
rect -74825 30932 -74783 31168
rect -74547 30932 -74443 31168
rect -74207 30932 -74103 31168
rect -73867 30932 -73783 31168
rect -73547 30932 -73443 31168
rect -73207 30932 -73103 31168
rect -72867 30932 -72783 31168
rect -72547 30932 -72443 31168
rect -72207 30932 -72103 31168
rect -71867 30932 -71783 31168
rect -71547 30932 -71443 31168
rect -71207 30932 -71103 31168
rect -70867 30932 -70783 31168
rect -70547 30932 -70443 31168
rect -70207 30932 -70103 31168
rect -69867 30932 -69783 31168
rect -69547 30932 -69443 31168
rect -69207 30932 -69103 31168
rect -68867 30932 -68783 31168
rect -68547 30932 -68443 31168
rect -68207 30932 -68103 31168
rect -67867 30932 -67783 31168
rect -67547 30932 -67443 31168
rect -67207 30932 -67103 31168
rect -66867 30932 -66783 31168
rect -66547 30932 -66443 31168
rect -66207 30932 -66103 31168
rect -65867 30932 -65783 31168
rect -65547 30932 -65443 31168
rect -65207 30932 -65103 31168
rect -64867 30932 -64783 31168
rect -64547 30932 -64443 31168
rect -64207 30932 -64103 31168
rect -63867 30932 -63783 31168
rect -63547 30932 -63443 31168
rect -63207 30932 -63103 31168
rect -62867 30932 -62783 31168
rect -62547 30932 -62443 31168
rect -62207 30932 -62103 31168
rect -61867 30932 -61783 31168
rect -61547 30932 -61443 31168
rect -61207 30932 -61103 31168
rect -60867 30932 -60783 31168
rect -60547 30932 -60443 31168
rect -60207 30932 -60103 31168
rect -59867 30932 -59783 31168
rect -59547 30932 -59443 31168
rect -59207 30932 -59103 31168
rect -58867 30932 -58825 31168
rect -74825 30890 -58825 30932
rect 9654 31168 34654 31210
rect 9654 30932 9696 31168
rect 9932 30932 10036 31168
rect 10272 30932 10376 31168
rect 10612 30932 10696 31168
rect 10932 30932 11036 31168
rect 11272 30932 11376 31168
rect 11612 30932 11696 31168
rect 11932 30932 12036 31168
rect 12272 30932 12376 31168
rect 12612 30932 12696 31168
rect 12932 30932 13036 31168
rect 13272 30932 13376 31168
rect 13612 30932 13696 31168
rect 13932 30932 14036 31168
rect 14272 30932 14376 31168
rect 14612 30932 14696 31168
rect 14932 30932 15036 31168
rect 15272 30932 15376 31168
rect 15612 30932 15696 31168
rect 15932 30932 16036 31168
rect 16272 30932 16376 31168
rect 16612 30932 16696 31168
rect 16932 30932 17036 31168
rect 17272 30932 17376 31168
rect 17612 30932 17696 31168
rect 17932 30932 18036 31168
rect 18272 30932 18376 31168
rect 18612 30932 18696 31168
rect 18932 30932 19036 31168
rect 19272 30932 19376 31168
rect 19612 30932 19696 31168
rect 19932 30932 20036 31168
rect 20272 30932 20376 31168
rect 20612 30932 20696 31168
rect 20932 30932 21036 31168
rect 21272 30932 21376 31168
rect 21612 30932 21696 31168
rect 21932 30932 22036 31168
rect 22272 30932 22376 31168
rect 22612 30932 22696 31168
rect 22932 30932 23036 31168
rect 23272 30932 23376 31168
rect 23612 30932 23696 31168
rect 23932 30932 24036 31168
rect 24272 30932 24376 31168
rect 24612 30932 24696 31168
rect 24932 30932 25036 31168
rect 25272 30932 25376 31168
rect 25612 30932 25696 31168
rect 25932 30932 26036 31168
rect 26272 30932 26376 31168
rect 26612 30932 26696 31168
rect 26932 30932 27036 31168
rect 27272 30932 27376 31168
rect 27612 30932 27696 31168
rect 27932 30932 28036 31168
rect 28272 30932 28376 31168
rect 28612 30932 28696 31168
rect 28932 30932 29036 31168
rect 29272 30932 29376 31168
rect 29612 30932 29696 31168
rect 29932 30932 30036 31168
rect 30272 30932 30376 31168
rect 30612 30932 30696 31168
rect 30932 30932 31036 31168
rect 31272 30932 31376 31168
rect 31612 30932 31696 31168
rect 31932 30932 32036 31168
rect 32272 30932 32376 31168
rect 32612 30932 32696 31168
rect 32932 30932 33036 31168
rect 33272 30932 33376 31168
rect 33612 30932 33696 31168
rect 33932 30932 34036 31168
rect 34272 30932 34376 31168
rect 34612 30932 34654 31168
rect 9654 30890 34654 30932
rect -74485 30828 -74165 30890
rect -74485 30592 -74443 30828
rect -74207 30592 -74165 30828
rect -74485 30508 -74165 30592
rect -74485 30272 -74443 30508
rect -74207 30272 -74165 30508
rect -74485 30210 -74165 30272
rect -73485 30828 -73165 30890
rect -73485 30592 -73443 30828
rect -73207 30592 -73165 30828
rect -73485 30508 -73165 30592
rect -73485 30272 -73443 30508
rect -73207 30272 -73165 30508
rect -73485 30210 -73165 30272
rect -72485 30828 -72165 30890
rect -72485 30592 -72443 30828
rect -72207 30592 -72165 30828
rect -72485 30508 -72165 30592
rect -72485 30272 -72443 30508
rect -72207 30272 -72165 30508
rect -72485 30210 -72165 30272
rect -71485 30828 -71165 30890
rect -71485 30592 -71443 30828
rect -71207 30592 -71165 30828
rect -71485 30508 -71165 30592
rect -71485 30272 -71443 30508
rect -71207 30272 -71165 30508
rect -71485 30210 -71165 30272
rect -70485 30828 -70165 30890
rect -70485 30592 -70443 30828
rect -70207 30592 -70165 30828
rect -70485 30508 -70165 30592
rect -70485 30272 -70443 30508
rect -70207 30272 -70165 30508
rect -70485 30210 -70165 30272
rect -69485 30828 -69165 30890
rect -69485 30592 -69443 30828
rect -69207 30592 -69165 30828
rect -69485 30508 -69165 30592
rect -69485 30272 -69443 30508
rect -69207 30272 -69165 30508
rect -69485 30210 -69165 30272
rect -68485 30828 -68165 30890
rect -68485 30592 -68443 30828
rect -68207 30592 -68165 30828
rect -68485 30508 -68165 30592
rect -68485 30272 -68443 30508
rect -68207 30272 -68165 30508
rect -68485 30210 -68165 30272
rect -67485 30828 -67165 30890
rect -67485 30592 -67443 30828
rect -67207 30592 -67165 30828
rect -67485 30508 -67165 30592
rect -67485 30272 -67443 30508
rect -67207 30272 -67165 30508
rect -67485 30210 -67165 30272
rect -66485 30828 -66165 30890
rect -66485 30592 -66443 30828
rect -66207 30592 -66165 30828
rect -66485 30508 -66165 30592
rect -66485 30272 -66443 30508
rect -66207 30272 -66165 30508
rect -66485 30210 -66165 30272
rect -65485 30828 -65165 30890
rect -65485 30592 -65443 30828
rect -65207 30592 -65165 30828
rect -65485 30508 -65165 30592
rect -65485 30272 -65443 30508
rect -65207 30272 -65165 30508
rect -65485 30210 -65165 30272
rect -64485 30828 -64165 30890
rect -64485 30592 -64443 30828
rect -64207 30592 -64165 30828
rect -64485 30508 -64165 30592
rect -64485 30272 -64443 30508
rect -64207 30272 -64165 30508
rect -64485 30210 -64165 30272
rect -63485 30828 -63165 30890
rect -63485 30592 -63443 30828
rect -63207 30592 -63165 30828
rect -63485 30508 -63165 30592
rect -63485 30272 -63443 30508
rect -63207 30272 -63165 30508
rect -63485 30210 -63165 30272
rect -62485 30828 -62165 30890
rect -62485 30592 -62443 30828
rect -62207 30592 -62165 30828
rect -62485 30508 -62165 30592
rect -62485 30272 -62443 30508
rect -62207 30272 -62165 30508
rect -62485 30210 -62165 30272
rect -61485 30828 -61165 30890
rect -61485 30592 -61443 30828
rect -61207 30592 -61165 30828
rect -61485 30508 -61165 30592
rect -61485 30272 -61443 30508
rect -61207 30272 -61165 30508
rect -61485 30210 -61165 30272
rect -60485 30828 -60165 30890
rect -60485 30592 -60443 30828
rect -60207 30592 -60165 30828
rect -60485 30508 -60165 30592
rect -60485 30272 -60443 30508
rect -60207 30272 -60165 30508
rect -60485 30210 -60165 30272
rect -59485 30828 -59165 30890
rect -59485 30592 -59443 30828
rect -59207 30592 -59165 30828
rect -59485 30508 -59165 30592
rect -59485 30272 -59443 30508
rect -59207 30272 -59165 30508
rect -59485 30210 -59165 30272
rect 9994 30828 10314 30890
rect 9994 30592 10036 30828
rect 10272 30592 10314 30828
rect 9994 30508 10314 30592
rect 9994 30272 10036 30508
rect 10272 30272 10314 30508
rect 9994 30210 10314 30272
rect 10994 30828 11314 30890
rect 10994 30592 11036 30828
rect 11272 30592 11314 30828
rect 10994 30508 11314 30592
rect 10994 30272 11036 30508
rect 11272 30272 11314 30508
rect 10994 30210 11314 30272
rect 11994 30828 12314 30890
rect 11994 30592 12036 30828
rect 12272 30592 12314 30828
rect 11994 30508 12314 30592
rect 11994 30272 12036 30508
rect 12272 30272 12314 30508
rect 11994 30210 12314 30272
rect 12994 30828 13314 30890
rect 12994 30592 13036 30828
rect 13272 30592 13314 30828
rect 12994 30508 13314 30592
rect 12994 30272 13036 30508
rect 13272 30272 13314 30508
rect 12994 30210 13314 30272
rect 13994 30828 14314 30890
rect 13994 30592 14036 30828
rect 14272 30592 14314 30828
rect 13994 30508 14314 30592
rect 13994 30272 14036 30508
rect 14272 30272 14314 30508
rect 13994 30210 14314 30272
rect 14994 30828 15314 30890
rect 14994 30592 15036 30828
rect 15272 30592 15314 30828
rect 14994 30508 15314 30592
rect 14994 30272 15036 30508
rect 15272 30272 15314 30508
rect 14994 30210 15314 30272
rect 15994 30828 16314 30890
rect 15994 30592 16036 30828
rect 16272 30592 16314 30828
rect 15994 30508 16314 30592
rect 15994 30272 16036 30508
rect 16272 30272 16314 30508
rect 15994 30210 16314 30272
rect 16994 30828 17314 30890
rect 16994 30592 17036 30828
rect 17272 30592 17314 30828
rect 16994 30508 17314 30592
rect 16994 30272 17036 30508
rect 17272 30272 17314 30508
rect 16994 30210 17314 30272
rect 17994 30828 18314 30890
rect 17994 30592 18036 30828
rect 18272 30592 18314 30828
rect 17994 30508 18314 30592
rect 17994 30272 18036 30508
rect 18272 30272 18314 30508
rect 17994 30210 18314 30272
rect 18994 30828 19314 30890
rect 18994 30592 19036 30828
rect 19272 30592 19314 30828
rect 18994 30508 19314 30592
rect 18994 30272 19036 30508
rect 19272 30272 19314 30508
rect 18994 30210 19314 30272
rect 19994 30828 20314 30890
rect 19994 30592 20036 30828
rect 20272 30592 20314 30828
rect 19994 30508 20314 30592
rect 19994 30272 20036 30508
rect 20272 30272 20314 30508
rect 19994 30210 20314 30272
rect 20994 30828 21314 30890
rect 20994 30592 21036 30828
rect 21272 30592 21314 30828
rect 20994 30508 21314 30592
rect 20994 30272 21036 30508
rect 21272 30272 21314 30508
rect 20994 30210 21314 30272
rect 21994 30828 22314 30890
rect 21994 30592 22036 30828
rect 22272 30592 22314 30828
rect 21994 30508 22314 30592
rect 21994 30272 22036 30508
rect 22272 30272 22314 30508
rect 21994 30210 22314 30272
rect 22994 30828 23314 30890
rect 22994 30592 23036 30828
rect 23272 30592 23314 30828
rect 22994 30508 23314 30592
rect 22994 30272 23036 30508
rect 23272 30272 23314 30508
rect 22994 30210 23314 30272
rect 23994 30828 24314 30890
rect 23994 30592 24036 30828
rect 24272 30592 24314 30828
rect 23994 30508 24314 30592
rect 23994 30272 24036 30508
rect 24272 30272 24314 30508
rect 23994 30210 24314 30272
rect 24994 30828 25314 30890
rect 24994 30592 25036 30828
rect 25272 30592 25314 30828
rect 24994 30508 25314 30592
rect 24994 30272 25036 30508
rect 25272 30272 25314 30508
rect 24994 30210 25314 30272
rect 25994 30828 26314 30890
rect 25994 30592 26036 30828
rect 26272 30592 26314 30828
rect 25994 30508 26314 30592
rect 25994 30272 26036 30508
rect 26272 30272 26314 30508
rect 25994 30210 26314 30272
rect 26994 30828 27314 30890
rect 26994 30592 27036 30828
rect 27272 30592 27314 30828
rect 26994 30508 27314 30592
rect 26994 30272 27036 30508
rect 27272 30272 27314 30508
rect 26994 30210 27314 30272
rect 27994 30828 28314 30890
rect 27994 30592 28036 30828
rect 28272 30592 28314 30828
rect 27994 30508 28314 30592
rect 27994 30272 28036 30508
rect 28272 30272 28314 30508
rect 27994 30210 28314 30272
rect 28994 30828 29314 30890
rect 28994 30592 29036 30828
rect 29272 30592 29314 30828
rect 28994 30508 29314 30592
rect 28994 30272 29036 30508
rect 29272 30272 29314 30508
rect 28994 30210 29314 30272
rect 29994 30828 30314 30890
rect 29994 30592 30036 30828
rect 30272 30592 30314 30828
rect 29994 30508 30314 30592
rect 29994 30272 30036 30508
rect 30272 30272 30314 30508
rect 29994 30210 30314 30272
rect 30994 30828 31314 30890
rect 30994 30592 31036 30828
rect 31272 30592 31314 30828
rect 30994 30508 31314 30592
rect 30994 30272 31036 30508
rect 31272 30272 31314 30508
rect 30994 30210 31314 30272
rect 31994 30828 32314 30890
rect 31994 30592 32036 30828
rect 32272 30592 32314 30828
rect 31994 30508 32314 30592
rect 31994 30272 32036 30508
rect 32272 30272 32314 30508
rect 31994 30210 32314 30272
rect 32994 30828 33314 30890
rect 32994 30592 33036 30828
rect 33272 30592 33314 30828
rect 32994 30508 33314 30592
rect 32994 30272 33036 30508
rect 33272 30272 33314 30508
rect 32994 30210 33314 30272
rect 33994 30828 34314 30890
rect 33994 30592 34036 30828
rect 34272 30592 34314 30828
rect 33994 30508 34314 30592
rect 33994 30272 34036 30508
rect 34272 30272 34314 30508
rect 33994 30210 34314 30272
rect -74825 30168 -58825 30210
rect -74825 29932 -74783 30168
rect -74547 29932 -74443 30168
rect -74207 29932 -74103 30168
rect -73867 29932 -73783 30168
rect -73547 29932 -73443 30168
rect -73207 29932 -73103 30168
rect -72867 29932 -72783 30168
rect -72547 29932 -72443 30168
rect -72207 29932 -72103 30168
rect -71867 29932 -71783 30168
rect -71547 29932 -71443 30168
rect -71207 29932 -71103 30168
rect -70867 29932 -70783 30168
rect -70547 29932 -70443 30168
rect -70207 29932 -70103 30168
rect -69867 29932 -69783 30168
rect -69547 29932 -69443 30168
rect -69207 29932 -69103 30168
rect -68867 29932 -68783 30168
rect -68547 29932 -68443 30168
rect -68207 29932 -68103 30168
rect -67867 29932 -67783 30168
rect -67547 29932 -67443 30168
rect -67207 29932 -67103 30168
rect -66867 29932 -66783 30168
rect -66547 29932 -66443 30168
rect -66207 29932 -66103 30168
rect -65867 29932 -65783 30168
rect -65547 29932 -65443 30168
rect -65207 29932 -65103 30168
rect -64867 29932 -64783 30168
rect -64547 29932 -64443 30168
rect -64207 29932 -64103 30168
rect -63867 29932 -63783 30168
rect -63547 29932 -63443 30168
rect -63207 29932 -63103 30168
rect -62867 29932 -62783 30168
rect -62547 29932 -62443 30168
rect -62207 29932 -62103 30168
rect -61867 29932 -61783 30168
rect -61547 29932 -61443 30168
rect -61207 29932 -61103 30168
rect -60867 29932 -60783 30168
rect -60547 29932 -60443 30168
rect -60207 29932 -60103 30168
rect -59867 29932 -59783 30168
rect -59547 29932 -59443 30168
rect -59207 29932 -59103 30168
rect -58867 29932 -58825 30168
rect -74825 29890 -58825 29932
rect 9654 30168 34654 30210
rect 9654 29932 9696 30168
rect 9932 29932 10036 30168
rect 10272 29932 10376 30168
rect 10612 29932 10696 30168
rect 10932 29932 11036 30168
rect 11272 29932 11376 30168
rect 11612 29932 11696 30168
rect 11932 29932 12036 30168
rect 12272 29932 12376 30168
rect 12612 29932 12696 30168
rect 12932 29932 13036 30168
rect 13272 29932 13376 30168
rect 13612 29932 13696 30168
rect 13932 29932 14036 30168
rect 14272 29932 14376 30168
rect 14612 29932 14696 30168
rect 14932 29932 15036 30168
rect 15272 29932 15376 30168
rect 15612 29932 15696 30168
rect 15932 29932 16036 30168
rect 16272 29932 16376 30168
rect 16612 29932 16696 30168
rect 16932 29932 17036 30168
rect 17272 29932 17376 30168
rect 17612 29932 17696 30168
rect 17932 29932 18036 30168
rect 18272 29932 18376 30168
rect 18612 29932 18696 30168
rect 18932 29932 19036 30168
rect 19272 29932 19376 30168
rect 19612 29932 19696 30168
rect 19932 29932 20036 30168
rect 20272 29932 20376 30168
rect 20612 29932 20696 30168
rect 20932 29932 21036 30168
rect 21272 29932 21376 30168
rect 21612 29932 21696 30168
rect 21932 29932 22036 30168
rect 22272 29932 22376 30168
rect 22612 29932 22696 30168
rect 22932 29932 23036 30168
rect 23272 29932 23376 30168
rect 23612 29932 23696 30168
rect 23932 29932 24036 30168
rect 24272 29932 24376 30168
rect 24612 29932 24696 30168
rect 24932 29932 25036 30168
rect 25272 29932 25376 30168
rect 25612 29932 25696 30168
rect 25932 29932 26036 30168
rect 26272 29932 26376 30168
rect 26612 29932 26696 30168
rect 26932 29932 27036 30168
rect 27272 29932 27376 30168
rect 27612 29932 27696 30168
rect 27932 29932 28036 30168
rect 28272 29932 28376 30168
rect 28612 29932 28696 30168
rect 28932 29932 29036 30168
rect 29272 29932 29376 30168
rect 29612 29932 29696 30168
rect 29932 29932 30036 30168
rect 30272 29932 30376 30168
rect 30612 29932 30696 30168
rect 30932 29932 31036 30168
rect 31272 29932 31376 30168
rect 31612 29932 31696 30168
rect 31932 29932 32036 30168
rect 32272 29932 32376 30168
rect 32612 29932 32696 30168
rect 32932 29932 33036 30168
rect 33272 29932 33376 30168
rect 33612 29932 33696 30168
rect 33932 29932 34036 30168
rect 34272 29932 34376 30168
rect 34612 29932 34654 30168
rect 9654 29890 34654 29932
rect -74485 29828 -74165 29890
rect -74485 29592 -74443 29828
rect -74207 29592 -74165 29828
rect -74485 29508 -74165 29592
rect -74485 29272 -74443 29508
rect -74207 29272 -74165 29508
rect -74485 29210 -74165 29272
rect -73485 29828 -73165 29890
rect -73485 29592 -73443 29828
rect -73207 29592 -73165 29828
rect -73485 29508 -73165 29592
rect -73485 29272 -73443 29508
rect -73207 29272 -73165 29508
rect -73485 29210 -73165 29272
rect -72485 29828 -72165 29890
rect -72485 29592 -72443 29828
rect -72207 29592 -72165 29828
rect -72485 29508 -72165 29592
rect -72485 29272 -72443 29508
rect -72207 29272 -72165 29508
rect -72485 29210 -72165 29272
rect -71485 29828 -71165 29890
rect -71485 29592 -71443 29828
rect -71207 29592 -71165 29828
rect -71485 29508 -71165 29592
rect -71485 29272 -71443 29508
rect -71207 29272 -71165 29508
rect -71485 29210 -71165 29272
rect -70485 29828 -70165 29890
rect -70485 29592 -70443 29828
rect -70207 29592 -70165 29828
rect -70485 29508 -70165 29592
rect -70485 29272 -70443 29508
rect -70207 29272 -70165 29508
rect -70485 29210 -70165 29272
rect -69485 29828 -69165 29890
rect -69485 29592 -69443 29828
rect -69207 29592 -69165 29828
rect -69485 29508 -69165 29592
rect -69485 29272 -69443 29508
rect -69207 29272 -69165 29508
rect -69485 29210 -69165 29272
rect -68485 29828 -68165 29890
rect -68485 29592 -68443 29828
rect -68207 29592 -68165 29828
rect -68485 29508 -68165 29592
rect -68485 29272 -68443 29508
rect -68207 29272 -68165 29508
rect -68485 29210 -68165 29272
rect -67485 29828 -67165 29890
rect -67485 29592 -67443 29828
rect -67207 29592 -67165 29828
rect -67485 29508 -67165 29592
rect -67485 29272 -67443 29508
rect -67207 29272 -67165 29508
rect -67485 29210 -67165 29272
rect -66485 29828 -66165 29890
rect -66485 29592 -66443 29828
rect -66207 29592 -66165 29828
rect -66485 29508 -66165 29592
rect -66485 29272 -66443 29508
rect -66207 29272 -66165 29508
rect -66485 29210 -66165 29272
rect -65485 29828 -65165 29890
rect -65485 29592 -65443 29828
rect -65207 29592 -65165 29828
rect -65485 29508 -65165 29592
rect -65485 29272 -65443 29508
rect -65207 29272 -65165 29508
rect -65485 29210 -65165 29272
rect -64485 29828 -64165 29890
rect -64485 29592 -64443 29828
rect -64207 29592 -64165 29828
rect -64485 29508 -64165 29592
rect -64485 29272 -64443 29508
rect -64207 29272 -64165 29508
rect -64485 29210 -64165 29272
rect -63485 29828 -63165 29890
rect -63485 29592 -63443 29828
rect -63207 29592 -63165 29828
rect -63485 29508 -63165 29592
rect -63485 29272 -63443 29508
rect -63207 29272 -63165 29508
rect -63485 29210 -63165 29272
rect -62485 29828 -62165 29890
rect -62485 29592 -62443 29828
rect -62207 29592 -62165 29828
rect -62485 29508 -62165 29592
rect -62485 29272 -62443 29508
rect -62207 29272 -62165 29508
rect -62485 29210 -62165 29272
rect -61485 29828 -61165 29890
rect -61485 29592 -61443 29828
rect -61207 29592 -61165 29828
rect -61485 29508 -61165 29592
rect -61485 29272 -61443 29508
rect -61207 29272 -61165 29508
rect -61485 29210 -61165 29272
rect -60485 29828 -60165 29890
rect -60485 29592 -60443 29828
rect -60207 29592 -60165 29828
rect -60485 29508 -60165 29592
rect -60485 29272 -60443 29508
rect -60207 29272 -60165 29508
rect -60485 29210 -60165 29272
rect -59485 29828 -59165 29890
rect -59485 29592 -59443 29828
rect -59207 29592 -59165 29828
rect -59485 29508 -59165 29592
rect -59485 29272 -59443 29508
rect -59207 29272 -59165 29508
rect -59485 29210 -59165 29272
rect 9994 29828 10314 29890
rect 9994 29592 10036 29828
rect 10272 29592 10314 29828
rect 9994 29508 10314 29592
rect 9994 29272 10036 29508
rect 10272 29272 10314 29508
rect 9994 29210 10314 29272
rect 10994 29828 11314 29890
rect 10994 29592 11036 29828
rect 11272 29592 11314 29828
rect 10994 29508 11314 29592
rect 10994 29272 11036 29508
rect 11272 29272 11314 29508
rect 10994 29210 11314 29272
rect 11994 29828 12314 29890
rect 11994 29592 12036 29828
rect 12272 29592 12314 29828
rect 11994 29508 12314 29592
rect 11994 29272 12036 29508
rect 12272 29272 12314 29508
rect 11994 29210 12314 29272
rect 12994 29828 13314 29890
rect 12994 29592 13036 29828
rect 13272 29592 13314 29828
rect 12994 29508 13314 29592
rect 12994 29272 13036 29508
rect 13272 29272 13314 29508
rect 12994 29210 13314 29272
rect 13994 29828 14314 29890
rect 13994 29592 14036 29828
rect 14272 29592 14314 29828
rect 13994 29508 14314 29592
rect 13994 29272 14036 29508
rect 14272 29272 14314 29508
rect 13994 29210 14314 29272
rect 14994 29828 15314 29890
rect 14994 29592 15036 29828
rect 15272 29592 15314 29828
rect 14994 29508 15314 29592
rect 14994 29272 15036 29508
rect 15272 29272 15314 29508
rect 14994 29210 15314 29272
rect 15994 29828 16314 29890
rect 15994 29592 16036 29828
rect 16272 29592 16314 29828
rect 15994 29508 16314 29592
rect 15994 29272 16036 29508
rect 16272 29272 16314 29508
rect 15994 29210 16314 29272
rect 16994 29828 17314 29890
rect 16994 29592 17036 29828
rect 17272 29592 17314 29828
rect 16994 29508 17314 29592
rect 16994 29272 17036 29508
rect 17272 29272 17314 29508
rect 16994 29210 17314 29272
rect 17994 29828 18314 29890
rect 17994 29592 18036 29828
rect 18272 29592 18314 29828
rect 17994 29508 18314 29592
rect 17994 29272 18036 29508
rect 18272 29272 18314 29508
rect 17994 29210 18314 29272
rect 18994 29828 19314 29890
rect 18994 29592 19036 29828
rect 19272 29592 19314 29828
rect 18994 29508 19314 29592
rect 18994 29272 19036 29508
rect 19272 29272 19314 29508
rect 18994 29210 19314 29272
rect 19994 29828 20314 29890
rect 19994 29592 20036 29828
rect 20272 29592 20314 29828
rect 19994 29508 20314 29592
rect 19994 29272 20036 29508
rect 20272 29272 20314 29508
rect 19994 29210 20314 29272
rect 20994 29828 21314 29890
rect 20994 29592 21036 29828
rect 21272 29592 21314 29828
rect 20994 29508 21314 29592
rect 20994 29272 21036 29508
rect 21272 29272 21314 29508
rect 20994 29210 21314 29272
rect 21994 29828 22314 29890
rect 21994 29592 22036 29828
rect 22272 29592 22314 29828
rect 21994 29508 22314 29592
rect 21994 29272 22036 29508
rect 22272 29272 22314 29508
rect 21994 29210 22314 29272
rect 22994 29828 23314 29890
rect 22994 29592 23036 29828
rect 23272 29592 23314 29828
rect 22994 29508 23314 29592
rect 22994 29272 23036 29508
rect 23272 29272 23314 29508
rect 22994 29210 23314 29272
rect 23994 29828 24314 29890
rect 23994 29592 24036 29828
rect 24272 29592 24314 29828
rect 23994 29508 24314 29592
rect 23994 29272 24036 29508
rect 24272 29272 24314 29508
rect 23994 29210 24314 29272
rect 24994 29828 25314 29890
rect 24994 29592 25036 29828
rect 25272 29592 25314 29828
rect 24994 29508 25314 29592
rect 24994 29272 25036 29508
rect 25272 29272 25314 29508
rect 24994 29210 25314 29272
rect 25994 29828 26314 29890
rect 25994 29592 26036 29828
rect 26272 29592 26314 29828
rect 25994 29508 26314 29592
rect 25994 29272 26036 29508
rect 26272 29272 26314 29508
rect 25994 29210 26314 29272
rect 26994 29828 27314 29890
rect 26994 29592 27036 29828
rect 27272 29592 27314 29828
rect 26994 29508 27314 29592
rect 26994 29272 27036 29508
rect 27272 29272 27314 29508
rect 26994 29210 27314 29272
rect 27994 29828 28314 29890
rect 27994 29592 28036 29828
rect 28272 29592 28314 29828
rect 27994 29508 28314 29592
rect 27994 29272 28036 29508
rect 28272 29272 28314 29508
rect 27994 29210 28314 29272
rect 28994 29828 29314 29890
rect 28994 29592 29036 29828
rect 29272 29592 29314 29828
rect 28994 29508 29314 29592
rect 28994 29272 29036 29508
rect 29272 29272 29314 29508
rect 28994 29210 29314 29272
rect 29994 29828 30314 29890
rect 29994 29592 30036 29828
rect 30272 29592 30314 29828
rect 29994 29508 30314 29592
rect 29994 29272 30036 29508
rect 30272 29272 30314 29508
rect 29994 29210 30314 29272
rect 30994 29828 31314 29890
rect 30994 29592 31036 29828
rect 31272 29592 31314 29828
rect 30994 29508 31314 29592
rect 30994 29272 31036 29508
rect 31272 29272 31314 29508
rect 30994 29210 31314 29272
rect 31994 29828 32314 29890
rect 31994 29592 32036 29828
rect 32272 29592 32314 29828
rect 31994 29508 32314 29592
rect 31994 29272 32036 29508
rect 32272 29272 32314 29508
rect 31994 29210 32314 29272
rect 32994 29828 33314 29890
rect 32994 29592 33036 29828
rect 33272 29592 33314 29828
rect 32994 29508 33314 29592
rect 32994 29272 33036 29508
rect 33272 29272 33314 29508
rect 32994 29210 33314 29272
rect 33994 29828 34314 29890
rect 33994 29592 34036 29828
rect 34272 29592 34314 29828
rect 33994 29508 34314 29592
rect 33994 29272 34036 29508
rect 34272 29272 34314 29508
rect 33994 29210 34314 29272
rect -74825 29168 -58825 29210
rect -74825 28932 -74783 29168
rect -74547 28932 -74443 29168
rect -74207 28932 -74103 29168
rect -73867 28932 -73783 29168
rect -73547 28932 -73443 29168
rect -73207 28932 -73103 29168
rect -72867 28932 -72783 29168
rect -72547 28932 -72443 29168
rect -72207 28932 -72103 29168
rect -71867 28932 -71783 29168
rect -71547 28932 -71443 29168
rect -71207 28932 -71103 29168
rect -70867 28932 -70783 29168
rect -70547 28932 -70443 29168
rect -70207 28932 -70103 29168
rect -69867 28932 -69783 29168
rect -69547 28932 -69443 29168
rect -69207 28932 -69103 29168
rect -68867 28932 -68783 29168
rect -68547 28932 -68443 29168
rect -68207 28932 -68103 29168
rect -67867 28932 -67783 29168
rect -67547 28932 -67443 29168
rect -67207 28932 -67103 29168
rect -66867 28932 -66783 29168
rect -66547 28932 -66443 29168
rect -66207 28932 -66103 29168
rect -65867 28932 -65783 29168
rect -65547 28932 -65443 29168
rect -65207 28932 -65103 29168
rect -64867 28932 -64783 29168
rect -64547 28932 -64443 29168
rect -64207 28932 -64103 29168
rect -63867 28932 -63783 29168
rect -63547 28932 -63443 29168
rect -63207 28932 -63103 29168
rect -62867 28932 -62783 29168
rect -62547 28932 -62443 29168
rect -62207 28932 -62103 29168
rect -61867 28932 -61783 29168
rect -61547 28932 -61443 29168
rect -61207 28932 -61103 29168
rect -60867 28932 -60783 29168
rect -60547 28932 -60443 29168
rect -60207 28932 -60103 29168
rect -59867 28932 -59783 29168
rect -59547 28932 -59443 29168
rect -59207 28932 -59103 29168
rect -58867 28932 -58825 29168
rect -74825 28890 -58825 28932
rect 9654 29168 34654 29210
rect 9654 28932 9696 29168
rect 9932 28932 10036 29168
rect 10272 28932 10376 29168
rect 10612 28932 10696 29168
rect 10932 28932 11036 29168
rect 11272 28932 11376 29168
rect 11612 28932 11696 29168
rect 11932 28932 12036 29168
rect 12272 28932 12376 29168
rect 12612 28932 12696 29168
rect 12932 28932 13036 29168
rect 13272 28932 13376 29168
rect 13612 28932 13696 29168
rect 13932 28932 14036 29168
rect 14272 28932 14376 29168
rect 14612 28932 14696 29168
rect 14932 28932 15036 29168
rect 15272 28932 15376 29168
rect 15612 28932 15696 29168
rect 15932 28932 16036 29168
rect 16272 28932 16376 29168
rect 16612 28932 16696 29168
rect 16932 28932 17036 29168
rect 17272 28932 17376 29168
rect 17612 28932 17696 29168
rect 17932 28932 18036 29168
rect 18272 28932 18376 29168
rect 18612 28932 18696 29168
rect 18932 28932 19036 29168
rect 19272 28932 19376 29168
rect 19612 28932 19696 29168
rect 19932 28932 20036 29168
rect 20272 28932 20376 29168
rect 20612 28932 20696 29168
rect 20932 28932 21036 29168
rect 21272 28932 21376 29168
rect 21612 28932 21696 29168
rect 21932 28932 22036 29168
rect 22272 28932 22376 29168
rect 22612 28932 22696 29168
rect 22932 28932 23036 29168
rect 23272 28932 23376 29168
rect 23612 28932 23696 29168
rect 23932 28932 24036 29168
rect 24272 28932 24376 29168
rect 24612 28932 24696 29168
rect 24932 28932 25036 29168
rect 25272 28932 25376 29168
rect 25612 28932 25696 29168
rect 25932 28932 26036 29168
rect 26272 28932 26376 29168
rect 26612 28932 26696 29168
rect 26932 28932 27036 29168
rect 27272 28932 27376 29168
rect 27612 28932 27696 29168
rect 27932 28932 28036 29168
rect 28272 28932 28376 29168
rect 28612 28932 28696 29168
rect 28932 28932 29036 29168
rect 29272 28932 29376 29168
rect 29612 28932 29696 29168
rect 29932 28932 30036 29168
rect 30272 28932 30376 29168
rect 30612 28932 30696 29168
rect 30932 28932 31036 29168
rect 31272 28932 31376 29168
rect 31612 28932 31696 29168
rect 31932 28932 32036 29168
rect 32272 28932 32376 29168
rect 32612 28932 32696 29168
rect 32932 28932 33036 29168
rect 33272 28932 33376 29168
rect 33612 28932 33696 29168
rect 33932 28932 34036 29168
rect 34272 28932 34376 29168
rect 34612 28932 34654 29168
rect 9654 28890 34654 28932
rect -74485 28828 -74165 28890
rect -74485 28592 -74443 28828
rect -74207 28592 -74165 28828
rect -74485 28550 -74165 28592
rect -73485 28828 -73165 28890
rect -73485 28592 -73443 28828
rect -73207 28592 -73165 28828
rect -73485 28550 -73165 28592
rect -72485 28828 -72165 28890
rect -72485 28592 -72443 28828
rect -72207 28592 -72165 28828
rect -72485 28550 -72165 28592
rect -71485 28828 -71165 28890
rect -71485 28592 -71443 28828
rect -71207 28592 -71165 28828
rect -71485 28550 -71165 28592
rect -70485 28828 -70165 28890
rect -70485 28592 -70443 28828
rect -70207 28592 -70165 28828
rect -70485 28550 -70165 28592
rect -69485 28828 -69165 28890
rect -69485 28592 -69443 28828
rect -69207 28592 -69165 28828
rect -69485 28550 -69165 28592
rect -68485 28828 -68165 28890
rect -68485 28592 -68443 28828
rect -68207 28592 -68165 28828
rect -68485 28550 -68165 28592
rect -67485 28828 -67165 28890
rect -67485 28592 -67443 28828
rect -67207 28592 -67165 28828
rect -67485 28550 -67165 28592
rect -66485 28828 -66165 28890
rect -66485 28592 -66443 28828
rect -66207 28592 -66165 28828
rect -66485 28550 -66165 28592
rect -65485 28828 -65165 28890
rect -65485 28592 -65443 28828
rect -65207 28592 -65165 28828
rect -65485 28550 -65165 28592
rect -64485 28828 -64165 28890
rect -64485 28592 -64443 28828
rect -64207 28592 -64165 28828
rect -64485 28550 -64165 28592
rect -63485 28828 -63165 28890
rect -63485 28592 -63443 28828
rect -63207 28592 -63165 28828
rect -63485 28550 -63165 28592
rect -62485 28828 -62165 28890
rect -62485 28592 -62443 28828
rect -62207 28592 -62165 28828
rect -62485 28550 -62165 28592
rect -61485 28828 -61165 28890
rect -61485 28592 -61443 28828
rect -61207 28592 -61165 28828
rect -61485 28550 -61165 28592
rect -60485 28828 -60165 28890
rect -60485 28592 -60443 28828
rect -60207 28592 -60165 28828
rect -60485 28550 -60165 28592
rect -59485 28828 -59165 28890
rect -59485 28592 -59443 28828
rect -59207 28592 -59165 28828
rect -59485 28550 -59165 28592
rect 9994 28828 10314 28890
rect 9994 28592 10036 28828
rect 10272 28592 10314 28828
rect 9994 28550 10314 28592
rect 10994 28828 11314 28890
rect 10994 28592 11036 28828
rect 11272 28592 11314 28828
rect 10994 28550 11314 28592
rect 11994 28828 12314 28890
rect 11994 28592 12036 28828
rect 12272 28592 12314 28828
rect 11994 28550 12314 28592
rect 12994 28828 13314 28890
rect 12994 28592 13036 28828
rect 13272 28592 13314 28828
rect 12994 28550 13314 28592
rect 13994 28828 14314 28890
rect 13994 28592 14036 28828
rect 14272 28592 14314 28828
rect 13994 28550 14314 28592
rect 14994 28828 15314 28890
rect 14994 28592 15036 28828
rect 15272 28592 15314 28828
rect 14994 28550 15314 28592
rect 15994 28828 16314 28890
rect 15994 28592 16036 28828
rect 16272 28592 16314 28828
rect 15994 28550 16314 28592
rect 16994 28828 17314 28890
rect 16994 28592 17036 28828
rect 17272 28592 17314 28828
rect 16994 28550 17314 28592
rect 17994 28828 18314 28890
rect 17994 28592 18036 28828
rect 18272 28592 18314 28828
rect 17994 28550 18314 28592
rect 18994 28828 19314 28890
rect 18994 28592 19036 28828
rect 19272 28592 19314 28828
rect 18994 28550 19314 28592
rect 19994 28828 20314 28890
rect 19994 28592 20036 28828
rect 20272 28592 20314 28828
rect 19994 28550 20314 28592
rect 20994 28828 21314 28890
rect 20994 28592 21036 28828
rect 21272 28592 21314 28828
rect 20994 28550 21314 28592
rect 21994 28828 22314 28890
rect 21994 28592 22036 28828
rect 22272 28592 22314 28828
rect 21994 28550 22314 28592
rect 22994 28828 23314 28890
rect 22994 28592 23036 28828
rect 23272 28592 23314 28828
rect 22994 28550 23314 28592
rect 23994 28828 24314 28890
rect 23994 28592 24036 28828
rect 24272 28592 24314 28828
rect 23994 28550 24314 28592
rect 24994 28828 25314 28890
rect 24994 28592 25036 28828
rect 25272 28592 25314 28828
rect 24994 28550 25314 28592
rect 25994 28828 26314 28890
rect 25994 28592 26036 28828
rect 26272 28592 26314 28828
rect 25994 28550 26314 28592
rect 26994 28828 27314 28890
rect 26994 28592 27036 28828
rect 27272 28592 27314 28828
rect 26994 28550 27314 28592
rect 27994 28828 28314 28890
rect 27994 28592 28036 28828
rect 28272 28592 28314 28828
rect 27994 28550 28314 28592
rect 28994 28828 29314 28890
rect 28994 28592 29036 28828
rect 29272 28592 29314 28828
rect 28994 28550 29314 28592
rect 29994 28828 30314 28890
rect 29994 28592 30036 28828
rect 30272 28592 30314 28828
rect 29994 28550 30314 28592
rect 30994 28828 31314 28890
rect 30994 28592 31036 28828
rect 31272 28592 31314 28828
rect 30994 28550 31314 28592
rect 31994 28828 32314 28890
rect 31994 28592 32036 28828
rect 32272 28592 32314 28828
rect 31994 28550 32314 28592
rect 32994 28828 33314 28890
rect 32994 28592 33036 28828
rect 33272 28592 33314 28828
rect 32994 28550 33314 28592
rect 33994 28828 34314 28890
rect 33994 28592 34036 28828
rect 34272 28592 34314 28828
rect 33994 28550 34314 28592
rect -72825 25918 -60825 26000
rect -72825 16082 -72708 25918
rect -60952 21850 -60825 25918
rect 20275 25918 32275 26000
tri -60825 21850 -58825 23850 sw
tri 18275 21850 20275 23850 se
rect 20275 21850 20392 25918
rect -60952 16082 -58825 21850
rect -72825 16030 -58825 16082
tri -58825 16030 -53005 21850 sw
tri 12455 16030 18275 21850 se
rect 18275 16082 20392 21850
rect 32148 16082 32275 25918
rect 18275 16030 32275 16082
rect -72825 16000 -53005 16030
tri -53005 16000 -52975 16030 sw
tri 12425 16000 12455 16030 se
rect 12455 16000 32275 16030
tri -60975 15850 -60825 16000 ne
rect -60825 15850 -52975 16000
tri -52975 15850 -52825 16000 sw
tri 12275 15850 12425 16000 se
rect 12425 15850 20275 16000
tri 20275 15850 20425 16000 nw
tri -60825 13850 -58825 15850 ne
rect -58825 13850 -52825 15850
tri -52825 13850 -50825 15850 sw
tri 10275 13850 12275 15850 se
rect 12275 13850 18275 15850
tri 18275 13850 20275 15850 nw
tri -58825 13820 -58795 13850 ne
rect -58795 13820 15306 13850
tri -58795 10881 -55856 13820 ne
rect -55856 13688 15306 13820
rect -55856 10881 -42308 13688
tri -55856 10436 -55411 10881 ne
rect -55411 10436 -42308 10881
tri -55411 10435 -55410 10436 ne
rect -55410 10435 -42308 10436
tri -55410 10308 -55283 10435 ne
rect -55283 10308 -42308 10435
tri -55283 10307 -55282 10308 ne
rect -55282 10307 -42308 10308
tri -55282 9972 -54947 10307 ne
rect -54947 9972 -42308 10307
tri -54947 9971 -54946 9972 ne
rect -54946 9971 -42308 9972
tri -54946 9959 -54934 9971 ne
rect -54934 9959 -42308 9971
tri -54934 9958 -54933 9959 ne
rect -54933 9958 -42308 9959
tri -54933 9949 -54924 9958 ne
rect -54924 9949 -42308 9958
tri -54924 9948 -54923 9949 ne
rect -54923 9948 -42308 9949
tri -54923 9947 -54922 9948 ne
rect -54922 9947 -42308 9948
tri -54922 8153 -53128 9947 ne
rect -53128 8153 -42308 9947
tri -53128 8150 -53125 8153 ne
rect -53125 8150 -42308 8153
tri -53125 7880 -52855 8150 ne
rect -52855 8012 -42308 8150
rect -40792 10881 -24233 13688
rect -40792 10436 -34520 10881
tri -34520 10436 -34075 10881 nw
tri -29024 10436 -28579 10881 ne
rect -28579 10436 -24233 10881
rect -40792 10435 -34521 10436
tri -34521 10435 -34520 10436 nw
tri -28579 10435 -28578 10436 ne
rect -28578 10435 -24233 10436
rect -40792 10308 -34648 10435
tri -34648 10308 -34521 10435 nw
tri -28578 10308 -28451 10435 ne
rect -28451 10308 -24233 10435
rect -40792 10307 -34649 10308
tri -34649 10307 -34648 10308 nw
tri -28451 10307 -28450 10308 ne
rect -28450 10307 -24233 10308
rect -40792 9972 -34984 10307
tri -34984 9972 -34649 10307 nw
tri -28450 9972 -28115 10307 ne
rect -28115 9972 -24233 10307
rect -40792 9971 -34985 9972
tri -34985 9971 -34984 9972 nw
tri -28115 9971 -28114 9972 ne
rect -28114 9971 -24233 9972
rect -40792 9959 -34997 9971
tri -34997 9959 -34985 9971 nw
tri -28114 9959 -28102 9971 ne
rect -28102 9959 -24233 9971
rect -40792 9958 -34998 9959
tri -34998 9958 -34997 9959 nw
tri -28102 9958 -28101 9959 ne
rect -28101 9958 -24233 9959
rect -40792 9949 -35007 9958
tri -35007 9949 -34998 9958 nw
tri -28101 9949 -28092 9958 ne
rect -28092 9949 -24233 9958
rect -40792 9948 -35008 9949
tri -35008 9948 -35007 9949 nw
tri -28092 9948 -28091 9949 ne
rect -28091 9948 -24233 9949
rect -40792 9947 -35009 9948
tri -35009 9947 -35008 9948 nw
tri -28091 9947 -28090 9948 ne
rect -28090 9947 -24233 9948
rect -40792 8389 -36567 9947
tri -36567 8389 -35009 9947 nw
tri -28090 9716 -27859 9947 ne
rect -27859 9716 -24233 9947
rect -27858 9715 -24233 9716
tri -27858 9233 -27376 9715 ne
rect -27376 9233 -24233 9715
rect -27375 9232 -24233 9233
tri -27375 8390 -26533 9232 ne
rect -26533 8390 -24233 9232
rect -26532 8389 -24233 8390
rect -40792 8331 -36625 8389
tri -36625 8331 -36567 8389 nw
tri -26532 8331 -26474 8389 ne
rect -26474 8331 -24233 8389
rect -40792 8330 -36626 8331
tri -36626 8330 -36625 8331 nw
rect -26473 8330 -24233 8331
rect -40792 8310 -36646 8330
tri -36646 8310 -36626 8330 nw
tri -26473 8310 -26453 8330 ne
rect -26453 8310 -24233 8330
rect -40792 8309 -36647 8310
tri -36647 8309 -36646 8310 nw
rect -26452 8309 -24233 8310
rect -40792 8299 -36657 8309
tri -36657 8299 -36647 8309 nw
tri -26452 8299 -26442 8309 ne
rect -26442 8299 -24233 8309
rect -40792 8298 -36658 8299
tri -36658 8298 -36657 8299 nw
rect -26441 8298 -24233 8299
rect -40792 8294 -36662 8298
tri -36662 8294 -36658 8298 nw
tri -26441 8294 -26437 8298 ne
rect -26437 8294 -24233 8298
rect -40792 8293 -36663 8294
tri -36663 8293 -36662 8294 nw
rect -26436 8293 -24233 8294
rect -40792 8292 -36664 8293
tri -36664 8292 -36663 8293 nw
tri -26436 8292 -26435 8293 ne
rect -26435 8292 -24233 8293
rect -40792 8291 -36665 8292
tri -36665 8291 -36664 8292 nw
rect -26434 8291 -24233 8292
rect -40792 8290 -36666 8291
tri -36666 8290 -36665 8291 nw
tri -26434 8290 -26433 8291 ne
rect -26433 8290 -24233 8291
rect -40792 8289 -36667 8290
tri -36667 8289 -36666 8290 nw
rect -26432 8289 -24233 8290
rect -40792 8172 -36784 8289
tri -36784 8172 -36667 8289 nw
tri -26431 8172 -26314 8289 ne
rect -26314 8172 -24233 8289
rect -40792 8153 -36803 8172
tri -36803 8153 -36784 8172 nw
tri -32971 8153 -32952 8172 se
rect -32952 8153 -32665 8172
rect -40792 8150 -36806 8153
tri -36806 8150 -36803 8153 nw
tri -32974 8150 -32971 8153 se
rect -32971 8150 -32665 8153
rect -40792 8012 -36955 8150
rect -52855 8001 -36955 8012
tri -36955 8001 -36806 8150 nw
tri -33123 8001 -32974 8150 se
rect -32974 8001 -32665 8150
rect -52855 7880 -37076 8001
tri -37076 7880 -36955 8001 nw
tri -33125 7999 -33123 8001 se
rect -33123 7999 -32665 8001
tri -33126 7998 -33125 7999 se
rect -33125 7998 -32665 7999
tri -33127 7997 -33126 7998 se
rect -33126 7997 -32665 7998
tri -33129 7995 -33127 7997 se
rect -33127 7995 -32665 7997
tri -33130 7994 -33129 7995 se
rect -33129 7994 -32665 7995
tri -33133 7991 -33130 7994 se
rect -33130 7991 -32665 7994
tri -33134 7990 -33133 7991 se
rect -33133 7990 -32665 7991
tri -33148 7976 -33134 7990 se
rect -33134 7976 -32665 7990
tri -33149 7975 -33148 7976 se
rect -33148 7975 -32665 7976
tri -33244 7880 -33149 7975 se
rect -33149 7880 -32665 7975
tri -52855 7850 -52825 7880 ne
rect -52825 7850 -37106 7880
tri -37106 7850 -37076 7880 nw
tri -33274 7850 -33244 7880 se
rect -33244 7850 -32665 7880
tri -33955 7169 -33274 7850 se
rect -33274 7478 -32665 7850
rect -30434 8153 -30147 8172
tri -30147 8153 -30128 8172 sw
tri -26314 8153 -26295 8172 ne
rect -26295 8153 -24233 8172
rect -30434 8150 -30128 8153
tri -30128 8150 -30125 8153 sw
tri -26295 8150 -26292 8153 ne
rect -26292 8150 -24233 8153
rect -30434 8001 -30125 8150
tri -30125 8001 -29976 8150 sw
tri -26292 8001 -26143 8150 ne
rect -26143 8012 -24233 8150
rect -16317 10881 242 13688
rect -16317 10436 -11971 10881
tri -11971 10436 -11526 10881 nw
tri -6475 10436 -6030 10881 ne
rect -6030 10436 242 10881
rect -16317 10435 -11972 10436
tri -6030 10435 -6029 10436 ne
rect -6029 10435 242 10436
rect -16317 10308 -12099 10435
tri -12099 10308 -11972 10435 nw
tri -6029 10308 -5902 10435 ne
rect -5902 10308 242 10435
rect -16317 10307 -12100 10308
rect -16317 9972 -12435 10307
tri -12435 9972 -12100 10307 nw
tri -5902 9972 -5566 10308 ne
rect -5566 9972 242 10308
rect -16317 9971 -12436 9972
rect -16317 9959 -12448 9971
tri -12448 9959 -12436 9971 nw
tri -5566 9959 -5553 9972 ne
rect -5553 9959 242 9972
rect -16317 9958 -12449 9959
rect -16317 9949 -12458 9958
tri -12458 9949 -12449 9958 nw
tri -5553 9949 -5543 9959 ne
rect -5543 9949 242 9959
rect -16317 9948 -12459 9949
tri -5543 9948 -5542 9949 ne
rect -5542 9948 242 9949
rect -16317 9947 -12460 9948
tri -5542 9947 -5541 9948 ne
rect -5541 9947 242 9948
rect -16317 8172 -14236 9947
tri -14236 8172 -12461 9947 nw
tri -5541 8172 -3766 9947 ne
rect -3766 8172 242 9947
rect -16317 8152 -14255 8172
tri -14255 8153 -14236 8172 nw
tri -10421 8153 -10402 8172 se
rect -10402 8153 -10115 8172
tri -10422 8152 -10421 8153 se
rect -10421 8152 -10115 8153
rect -16317 8151 -14256 8152
tri -10423 8151 -10422 8152 se
rect -10422 8151 -10115 8152
rect -16317 8150 -14257 8151
tri -10424 8150 -10423 8151 se
rect -10423 8150 -10115 8151
rect -16317 8012 -14527 8150
rect -30434 7999 -29976 8001
tri -29976 7999 -29974 8001 sw
rect -26143 8000 -14527 8012
rect -26142 7999 -14527 8000
rect -30434 7998 -29974 7999
tri -29974 7998 -29973 7999 sw
tri -26142 7998 -26141 7999 ne
rect -26141 7998 -14527 7999
rect -30434 7997 -29973 7998
tri -29973 7997 -29972 7998 sw
rect -26140 7997 -14527 7998
rect -30434 7995 -29972 7997
tri -29972 7995 -29970 7997 sw
tri -26140 7995 -26138 7997 ne
rect -26138 7995 -14527 7997
rect -30434 7994 -29970 7995
tri -29970 7994 -29969 7995 sw
rect -26137 7994 -14527 7995
rect -30434 7991 -29969 7994
tri -29969 7991 -29966 7994 sw
tri -26137 7991 -26134 7994 ne
rect -26134 7991 -14527 7994
rect -30434 7990 -29966 7991
tri -29966 7990 -29965 7991 sw
rect -26133 7990 -14527 7991
rect -30434 7976 -29965 7990
tri -29965 7976 -29951 7990 sw
tri -26133 7976 -26119 7990 ne
rect -26119 7976 -14527 7990
rect -30434 7975 -29951 7976
tri -29951 7975 -29950 7976 sw
rect -26118 7975 -14527 7976
rect -30434 7880 -29950 7975
tri -29950 7880 -29855 7975 sw
tri -26118 7880 -26023 7975 ne
rect -26023 7880 -14527 7975
tri -14527 7880 -14257 8150 nw
tri -10694 7880 -10424 8150 se
rect -10424 7880 -10115 8150
rect -30434 7850 -29855 7880
tri -29855 7850 -29825 7880 sw
tri -26023 7850 -25993 7880 ne
rect -25993 7850 -14557 7880
tri -14557 7850 -14527 7880 nw
tri -10724 7850 -10694 7880 se
rect -10694 7850 -10115 7880
rect -30434 7478 -29825 7850
rect -33274 7191 -32952 7478
tri -32952 7191 -32665 7478 nw
tri -30434 7191 -30147 7478 ne
rect -30147 7191 -29825 7478
tri -29825 7191 -29166 7850 sw
tri -11383 7191 -10724 7850 se
rect -10724 7478 -10115 7850
rect -7884 8150 -7597 8172
tri -7597 8150 -7575 8172 sw
tri -3766 8150 -3744 8172 ne
rect -3744 8150 242 8172
rect -7884 7880 -7575 8150
tri -7575 7880 -7305 8150 sw
tri -3744 7880 -3474 8150 ne
rect -3474 8012 242 8150
rect 1758 10881 15306 13688
tri 15306 10881 18275 13850 nw
rect 1758 10436 14861 10881
tri 14861 10436 15306 10881 nw
rect 1758 10308 14733 10436
tri 14733 10308 14861 10436 nw
rect 1758 9972 14397 10308
tri 14397 9972 14733 10308 nw
rect 1758 9959 14384 9972
tri 14384 9959 14397 9972 nw
rect 1758 9949 14374 9959
tri 14374 9949 14384 9959 nw
rect 1758 9948 14373 9949
tri 14373 9948 14374 9949 nw
rect 1758 9947 14372 9948
tri 14372 9947 14373 9948 nw
rect 1758 8172 12597 9947
tri 12597 8172 14372 9947 nw
rect 1758 8012 12305 8172
rect -3474 7880 12305 8012
tri 12305 7880 12597 8172 nw
rect -7884 7478 -7305 7880
rect -10724 7191 -10402 7478
tri -10402 7191 -10115 7478 nw
tri -7884 7191 -7597 7478 ne
rect -7597 7191 -7305 7478
tri -7305 7191 -6616 7880 sw
tri -3474 7850 -3444 7880 ne
rect -3444 7850 12275 7880
tri 12275 7850 12305 7880 nw
rect -33274 7169 -32974 7191
tri -32974 7169 -32952 7191 nw
tri -30147 7169 -30125 7191 ne
rect -30125 7169 -29166 7191
tri -29166 7169 -29144 7191 sw
tri -11405 7169 -11383 7191 se
rect -11383 7169 -10424 7191
tri -10424 7169 -10402 7191 nw
tri -7597 7169 -7575 7191 ne
rect -7575 7169 -6616 7191
tri -6616 7169 -6594 7191 sw
tri -34936 6188 -33955 7169 se
rect -33955 6210 -33933 7169
tri -33933 6210 -32974 7169 nw
tri -30125 6210 -29166 7169 ne
rect -29166 6210 -29144 7169
tri -29144 6210 -28185 7169 sw
tri -12364 6210 -11405 7169 se
rect -11405 6210 -11383 7169
tri -11383 6210 -10424 7169 nw
tri -7575 6210 -6616 7169 ne
rect -6616 6210 -6594 7169
tri -6594 6210 -5635 7169 sw
tri -33955 6188 -33933 6210 nw
tri -29166 6188 -29144 6210 ne
rect -29144 6188 -28185 6210
tri -28185 6188 -28163 6210 sw
tri -72825 2600 -70825 4600 se
rect -70825 2895 -62825 4600
tri -62825 2895 -61120 4600 sw
rect -34936 3381 -34243 6188
tri -34243 5900 -33955 6188 nw
tri -29144 5900 -28856 6188 ne
tri -34243 3381 -33955 3669 sw
tri -29144 3381 -28856 3669 se
rect -28856 3381 -28163 6188
tri -34936 2895 -34450 3381 ne
rect -34450 2895 -33955 3381
tri -33955 2895 -33469 3381 sw
tri -29630 2895 -29144 3381 se
rect -29144 2895 -28649 3381
tri -28649 2895 -28163 3381 nw
tri -12386 6188 -12364 6210 se
rect -12364 6188 -11405 6210
tri -11405 6188 -11383 6210 nw
tri -6616 6188 -6594 6210 ne
rect -6594 6188 -5635 6210
tri -5635 6188 -5613 6210 sw
rect -12386 3381 -11693 6188
tri -11693 5900 -11405 6188 nw
tri -6594 5900 -6306 6188 ne
tri -11693 3381 -11405 3669 sw
tri -6594 3381 -6306 3669 se
rect -6306 3381 -5613 6188
tri -12386 2895 -11900 3381 ne
rect -11900 2895 -11405 3381
tri -11405 2895 -10919 3381 sw
tri -7080 2895 -6594 3381 se
rect -6594 2895 -6099 3381
tri -6099 2895 -5613 3381 nw
tri 20571 2896 22275 4600 se
rect 22275 2896 30275 4600
tri 30275 2896 31979 4600 sw
tri 20570 2895 20571 2896 se
rect 20571 2895 31979 2896
rect -70825 2600 -61120 2895
tri -61120 2600 -60825 2895 sw
rect -72825 2350 -60825 2600
rect -34450 2894 -33469 2895
tri -33469 2894 -33468 2895 sw
tri -29631 2894 -29630 2895 se
rect -29630 2894 -28650 2895
tri -28650 2894 -28649 2895 nw
rect -11900 2894 -10919 2895
tri -10919 2894 -10918 2895 sw
tri -7081 2894 -7080 2895 se
rect -7080 2894 -6100 2895
tri -6100 2894 -6099 2895 nw
tri 20569 2894 20570 2895 se
rect 20570 2894 31979 2895
rect -34450 2600 -33468 2894
tri -33468 2600 -33174 2894 sw
tri -29925 2600 -29631 2894 se
rect -29631 2600 -28650 2894
rect -34450 2350 -33174 2600
tri -33174 2350 -32924 2600 sw
tri -30175 2350 -29925 2600 se
rect -29925 2350 -28650 2600
rect -11900 2350 -10918 2894
rect -72825 2276 -32924 2350
tri -32924 2276 -32850 2350 sw
rect -72825 2198 -32850 2276
rect -72825 -2198 -42308 2198
rect -40792 50 -32850 2198
rect -40792 -2198 -35250 50
rect -72825 -2350 -35250 -2198
tri -35250 -2350 -32850 50 nw
tri -30250 2275 -30175 2350 se
rect -30175 2276 -10918 2350
tri -10918 2276 -10300 2894 sw
rect -30175 2275 -10300 2276
rect -30250 50 -10300 2275
tri -30250 -2350 -27850 50 ne
rect -27850 -2350 -12700 50
tri -12700 -2350 -10300 50 nw
tri -7700 2275 -7081 2894 se
rect -7081 2350 -6100 2894
tri 20275 2600 20569 2894 se
rect 20569 2600 31979 2894
tri 31979 2600 32275 2896 sw
rect 20275 2350 32275 2600
rect -7081 2275 32275 2350
rect -7700 2198 32275 2275
rect -7700 50 242 2198
tri -7700 -2350 -5300 50 ne
rect -5300 -2198 242 50
rect 1758 -2198 32275 2198
rect -5300 -2350 32275 -2198
rect -72825 -2600 -60825 -2350
tri -72825 -4600 -70825 -2600 ne
rect -70825 -4600 -62825 -2600
tri -62825 -4600 -60825 -2600 nw
tri -52855 -7880 -52825 -7850 se
rect -52825 -7880 -28125 -7850
tri -58795 -13820 -52855 -7880 se
rect -52855 -8012 -28125 -7880
rect -52855 -13688 -42308 -8012
rect -40792 -8017 -28125 -8012
rect -40792 -13688 -29423 -8017
rect -52855 -13693 -29423 -13688
rect -28227 -13693 -28125 -8017
rect -52855 -13820 -28125 -13693
tri -58805 -13830 -58795 -13820 se
rect -58795 -13830 -28125 -13820
tri -58814 -13839 -58805 -13830 se
rect -58805 -13839 -28125 -13830
tri -58825 -13850 -58814 -13839 se
rect -58814 -13850 -28125 -13839
tri -60975 -16000 -58825 -13850 se
rect -58825 -16000 -52975 -13850
tri -52975 -16000 -50825 -13850 nw
rect -72825 -16030 -53005 -16000
tri -53005 -16030 -52975 -16000 nw
rect -72825 -16082 -58825 -16030
rect -72825 -25918 -72708 -16082
rect -60952 -21850 -58825 -16082
tri -58825 -21850 -53005 -16030 nw
rect -60952 -22550 -59525 -21850
tri -59525 -22550 -58825 -21850 nw
rect -60952 -25918 -60825 -22550
tri -60825 -23850 -59525 -22550 nw
tri -35425 -23850 -34125 -22550 se
rect -34125 -23850 -28125 -13850
tri -36125 -24550 -35425 -23850 se
rect -35425 -24550 -28125 -23850
rect -72825 -26000 -60825 -25918
tri -37545 -25970 -36125 -24550 se
rect -36125 -25970 -29545 -24550
tri -29545 -25970 -28125 -24550 nw
tri -37575 -26000 -37545 -25970 se
rect -37545 -26000 -29575 -25970
tri -29575 -26000 -29545 -25970 nw
tri -40125 -28550 -37575 -26000 se
rect -37575 -28550 -32125 -26000
tri -32125 -28550 -29575 -26000 nw
rect -74485 -28592 -74165 -28550
rect -74485 -28828 -74443 -28592
rect -74207 -28828 -74165 -28592
rect -74485 -28890 -74165 -28828
rect -73485 -28592 -73165 -28550
rect -73485 -28828 -73443 -28592
rect -73207 -28828 -73165 -28592
rect -73485 -28890 -73165 -28828
rect -72485 -28592 -72165 -28550
rect -72485 -28828 -72443 -28592
rect -72207 -28828 -72165 -28592
rect -72485 -28890 -72165 -28828
rect -71485 -28592 -71165 -28550
rect -71485 -28828 -71443 -28592
rect -71207 -28828 -71165 -28592
rect -71485 -28890 -71165 -28828
rect -70485 -28592 -70165 -28550
rect -70485 -28828 -70443 -28592
rect -70207 -28828 -70165 -28592
rect -70485 -28890 -70165 -28828
rect -69485 -28592 -69165 -28550
rect -69485 -28828 -69443 -28592
rect -69207 -28828 -69165 -28592
rect -69485 -28890 -69165 -28828
rect -68485 -28592 -68165 -28550
rect -68485 -28828 -68443 -28592
rect -68207 -28828 -68165 -28592
rect -68485 -28890 -68165 -28828
rect -67485 -28592 -67165 -28550
rect -67485 -28828 -67443 -28592
rect -67207 -28828 -67165 -28592
rect -67485 -28890 -67165 -28828
rect -66485 -28592 -66165 -28550
rect -66485 -28828 -66443 -28592
rect -66207 -28828 -66165 -28592
rect -66485 -28890 -66165 -28828
rect -65485 -28592 -65165 -28550
rect -65485 -28828 -65443 -28592
rect -65207 -28828 -65165 -28592
rect -65485 -28890 -65165 -28828
rect -64485 -28592 -64165 -28550
rect -64485 -28828 -64443 -28592
rect -64207 -28828 -64165 -28592
rect -64485 -28890 -64165 -28828
rect -63485 -28592 -63165 -28550
rect -63485 -28828 -63443 -28592
rect -63207 -28828 -63165 -28592
rect -63485 -28890 -63165 -28828
rect -62485 -28592 -62165 -28550
rect -62485 -28828 -62443 -28592
rect -62207 -28828 -62165 -28592
rect -62485 -28890 -62165 -28828
rect -61485 -28592 -61165 -28550
rect -61485 -28828 -61443 -28592
rect -61207 -28828 -61165 -28592
rect -61485 -28890 -61165 -28828
rect -60485 -28592 -60165 -28550
rect -60485 -28828 -60443 -28592
rect -60207 -28828 -60165 -28592
rect -60485 -28890 -60165 -28828
rect -59485 -28592 -59165 -28550
rect -59485 -28828 -59443 -28592
rect -59207 -28828 -59165 -28592
rect -59485 -28890 -59165 -28828
rect -58485 -28592 -58165 -28550
rect -58485 -28828 -58443 -28592
rect -58207 -28828 -58165 -28592
rect -58485 -28890 -58165 -28828
rect -57485 -28592 -57165 -28550
rect -57485 -28828 -57443 -28592
rect -57207 -28828 -57165 -28592
rect -57485 -28890 -57165 -28828
rect -56485 -28592 -56165 -28550
rect -56485 -28828 -56443 -28592
rect -56207 -28828 -56165 -28592
rect -56485 -28890 -56165 -28828
rect -55485 -28592 -55165 -28550
rect -55485 -28828 -55443 -28592
rect -55207 -28828 -55165 -28592
rect -55485 -28890 -55165 -28828
rect -54485 -28592 -54165 -28550
rect -54485 -28828 -54443 -28592
rect -54207 -28828 -54165 -28592
rect -54485 -28890 -54165 -28828
rect -53485 -28592 -53165 -28550
rect -53485 -28828 -53443 -28592
rect -53207 -28828 -53165 -28592
rect -53485 -28890 -53165 -28828
rect -52485 -28592 -52165 -28550
rect -52485 -28828 -52443 -28592
rect -52207 -28828 -52165 -28592
rect -52485 -28890 -52165 -28828
rect -51485 -28592 -51165 -28550
rect -51485 -28828 -51443 -28592
rect -51207 -28828 -51165 -28592
rect -51485 -28890 -51165 -28828
rect -50485 -28592 -50165 -28550
rect -50485 -28828 -50443 -28592
rect -50207 -28828 -50165 -28592
rect -50485 -28890 -50165 -28828
rect -49485 -28592 -49165 -28550
rect -49485 -28828 -49443 -28592
rect -49207 -28828 -49165 -28592
rect -49485 -28890 -49165 -28828
tri -40465 -28890 -40125 -28550 se
rect -40125 -28890 -32465 -28550
tri -32465 -28890 -32125 -28550 nw
rect -74825 -28932 -48825 -28890
rect -74825 -29168 -74783 -28932
rect -74547 -29168 -74443 -28932
rect -74207 -29168 -74103 -28932
rect -73867 -29168 -73783 -28932
rect -73547 -29168 -73443 -28932
rect -73207 -29168 -73103 -28932
rect -72867 -29168 -72783 -28932
rect -72547 -29168 -72443 -28932
rect -72207 -29168 -72103 -28932
rect -71867 -29168 -71783 -28932
rect -71547 -29168 -71443 -28932
rect -71207 -29168 -71103 -28932
rect -70867 -29168 -70783 -28932
rect -70547 -29168 -70443 -28932
rect -70207 -29168 -70103 -28932
rect -69867 -29168 -69783 -28932
rect -69547 -29168 -69443 -28932
rect -69207 -29168 -69103 -28932
rect -68867 -29168 -68783 -28932
rect -68547 -29168 -68443 -28932
rect -68207 -29168 -68103 -28932
rect -67867 -29168 -67783 -28932
rect -67547 -29168 -67443 -28932
rect -67207 -29168 -67103 -28932
rect -66867 -29168 -66783 -28932
rect -66547 -29168 -66443 -28932
rect -66207 -29168 -66103 -28932
rect -65867 -29168 -65783 -28932
rect -65547 -29168 -65443 -28932
rect -65207 -29168 -65103 -28932
rect -64867 -29168 -64783 -28932
rect -64547 -29168 -64443 -28932
rect -64207 -29168 -64103 -28932
rect -63867 -29168 -63783 -28932
rect -63547 -29168 -63443 -28932
rect -63207 -29168 -63103 -28932
rect -62867 -29168 -62783 -28932
rect -62547 -29168 -62443 -28932
rect -62207 -29168 -62103 -28932
rect -61867 -29168 -61783 -28932
rect -61547 -29168 -61443 -28932
rect -61207 -29168 -61103 -28932
rect -60867 -29168 -60783 -28932
rect -60547 -29168 -60443 -28932
rect -60207 -29168 -60103 -28932
rect -59867 -29168 -59783 -28932
rect -59547 -29168 -59443 -28932
rect -59207 -29168 -59103 -28932
rect -58867 -29168 -58783 -28932
rect -58547 -29168 -58443 -28932
rect -58207 -29168 -58103 -28932
rect -57867 -29168 -57783 -28932
rect -57547 -29168 -57443 -28932
rect -57207 -29168 -57103 -28932
rect -56867 -29168 -56783 -28932
rect -56547 -29168 -56443 -28932
rect -56207 -29168 -56103 -28932
rect -55867 -29168 -55783 -28932
rect -55547 -29168 -55443 -28932
rect -55207 -29168 -55103 -28932
rect -54867 -29168 -54783 -28932
rect -54547 -29168 -54443 -28932
rect -54207 -29168 -54103 -28932
rect -53867 -29168 -53783 -28932
rect -53547 -29168 -53443 -28932
rect -53207 -29168 -53103 -28932
rect -52867 -29168 -52783 -28932
rect -52547 -29168 -52443 -28932
rect -52207 -29168 -52103 -28932
rect -51867 -29168 -51783 -28932
rect -51547 -29168 -51443 -28932
rect -51207 -29168 -51103 -28932
rect -50867 -29168 -50783 -28932
rect -50547 -29168 -50443 -28932
rect -50207 -29168 -50103 -28932
rect -49867 -29168 -49783 -28932
rect -49547 -29168 -49443 -28932
rect -49207 -29168 -49103 -28932
rect -48867 -29168 -48825 -28932
rect -74825 -29210 -48825 -29168
tri -40785 -29210 -40465 -28890 se
rect -40465 -29210 -32785 -28890
tri -32785 -29210 -32465 -28890 nw
rect -74485 -29272 -74165 -29210
rect -74485 -29508 -74443 -29272
rect -74207 -29508 -74165 -29272
rect -74485 -29592 -74165 -29508
rect -74485 -29828 -74443 -29592
rect -74207 -29828 -74165 -29592
rect -74485 -29890 -74165 -29828
rect -73485 -29272 -73165 -29210
rect -73485 -29508 -73443 -29272
rect -73207 -29508 -73165 -29272
rect -73485 -29592 -73165 -29508
rect -73485 -29828 -73443 -29592
rect -73207 -29828 -73165 -29592
rect -73485 -29890 -73165 -29828
rect -72485 -29272 -72165 -29210
rect -72485 -29508 -72443 -29272
rect -72207 -29508 -72165 -29272
rect -72485 -29592 -72165 -29508
rect -72485 -29828 -72443 -29592
rect -72207 -29828 -72165 -29592
rect -72485 -29890 -72165 -29828
rect -71485 -29272 -71165 -29210
rect -71485 -29508 -71443 -29272
rect -71207 -29508 -71165 -29272
rect -71485 -29592 -71165 -29508
rect -71485 -29828 -71443 -29592
rect -71207 -29828 -71165 -29592
rect -71485 -29890 -71165 -29828
rect -70485 -29272 -70165 -29210
rect -70485 -29508 -70443 -29272
rect -70207 -29508 -70165 -29272
rect -70485 -29592 -70165 -29508
rect -70485 -29828 -70443 -29592
rect -70207 -29828 -70165 -29592
rect -70485 -29890 -70165 -29828
rect -69485 -29272 -69165 -29210
rect -69485 -29508 -69443 -29272
rect -69207 -29508 -69165 -29272
rect -69485 -29592 -69165 -29508
rect -69485 -29828 -69443 -29592
rect -69207 -29828 -69165 -29592
rect -69485 -29890 -69165 -29828
rect -68485 -29272 -68165 -29210
rect -68485 -29508 -68443 -29272
rect -68207 -29508 -68165 -29272
rect -68485 -29592 -68165 -29508
rect -68485 -29828 -68443 -29592
rect -68207 -29828 -68165 -29592
rect -68485 -29890 -68165 -29828
rect -67485 -29272 -67165 -29210
rect -67485 -29508 -67443 -29272
rect -67207 -29508 -67165 -29272
rect -67485 -29592 -67165 -29508
rect -67485 -29828 -67443 -29592
rect -67207 -29828 -67165 -29592
rect -67485 -29890 -67165 -29828
rect -66485 -29272 -66165 -29210
rect -66485 -29508 -66443 -29272
rect -66207 -29508 -66165 -29272
rect -66485 -29592 -66165 -29508
rect -66485 -29828 -66443 -29592
rect -66207 -29828 -66165 -29592
rect -66485 -29890 -66165 -29828
rect -65485 -29272 -65165 -29210
rect -65485 -29508 -65443 -29272
rect -65207 -29508 -65165 -29272
rect -65485 -29592 -65165 -29508
rect -65485 -29828 -65443 -29592
rect -65207 -29828 -65165 -29592
rect -65485 -29890 -65165 -29828
rect -64485 -29272 -64165 -29210
rect -64485 -29508 -64443 -29272
rect -64207 -29508 -64165 -29272
rect -64485 -29592 -64165 -29508
rect -64485 -29828 -64443 -29592
rect -64207 -29828 -64165 -29592
rect -64485 -29890 -64165 -29828
rect -63485 -29272 -63165 -29210
rect -63485 -29508 -63443 -29272
rect -63207 -29508 -63165 -29272
rect -63485 -29592 -63165 -29508
rect -63485 -29828 -63443 -29592
rect -63207 -29828 -63165 -29592
rect -63485 -29890 -63165 -29828
rect -62485 -29272 -62165 -29210
rect -62485 -29508 -62443 -29272
rect -62207 -29508 -62165 -29272
rect -62485 -29592 -62165 -29508
rect -62485 -29828 -62443 -29592
rect -62207 -29828 -62165 -29592
rect -62485 -29890 -62165 -29828
rect -61485 -29272 -61165 -29210
rect -61485 -29508 -61443 -29272
rect -61207 -29508 -61165 -29272
rect -61485 -29592 -61165 -29508
rect -61485 -29828 -61443 -29592
rect -61207 -29828 -61165 -29592
rect -61485 -29890 -61165 -29828
rect -60485 -29272 -60165 -29210
rect -60485 -29508 -60443 -29272
rect -60207 -29508 -60165 -29272
rect -60485 -29592 -60165 -29508
rect -60485 -29828 -60443 -29592
rect -60207 -29828 -60165 -29592
rect -60485 -29890 -60165 -29828
rect -59485 -29272 -59165 -29210
rect -59485 -29508 -59443 -29272
rect -59207 -29508 -59165 -29272
rect -59485 -29592 -59165 -29508
rect -59485 -29828 -59443 -29592
rect -59207 -29828 -59165 -29592
rect -59485 -29890 -59165 -29828
rect -58485 -29272 -58165 -29210
rect -58485 -29508 -58443 -29272
rect -58207 -29508 -58165 -29272
rect -58485 -29592 -58165 -29508
rect -58485 -29828 -58443 -29592
rect -58207 -29828 -58165 -29592
rect -58485 -29890 -58165 -29828
rect -57485 -29272 -57165 -29210
rect -57485 -29508 -57443 -29272
rect -57207 -29508 -57165 -29272
rect -57485 -29592 -57165 -29508
rect -57485 -29828 -57443 -29592
rect -57207 -29828 -57165 -29592
rect -57485 -29890 -57165 -29828
rect -56485 -29272 -56165 -29210
rect -56485 -29508 -56443 -29272
rect -56207 -29508 -56165 -29272
rect -56485 -29592 -56165 -29508
rect -56485 -29828 -56443 -29592
rect -56207 -29828 -56165 -29592
rect -56485 -29890 -56165 -29828
rect -55485 -29272 -55165 -29210
rect -55485 -29508 -55443 -29272
rect -55207 -29508 -55165 -29272
rect -55485 -29592 -55165 -29508
rect -55485 -29828 -55443 -29592
rect -55207 -29828 -55165 -29592
rect -55485 -29890 -55165 -29828
rect -54485 -29272 -54165 -29210
rect -54485 -29508 -54443 -29272
rect -54207 -29508 -54165 -29272
rect -54485 -29592 -54165 -29508
rect -54485 -29828 -54443 -29592
rect -54207 -29828 -54165 -29592
rect -54485 -29890 -54165 -29828
rect -53485 -29272 -53165 -29210
rect -53485 -29508 -53443 -29272
rect -53207 -29508 -53165 -29272
rect -53485 -29592 -53165 -29508
rect -53485 -29828 -53443 -29592
rect -53207 -29828 -53165 -29592
rect -53485 -29890 -53165 -29828
rect -52485 -29272 -52165 -29210
rect -52485 -29508 -52443 -29272
rect -52207 -29508 -52165 -29272
rect -52485 -29592 -52165 -29508
rect -52485 -29828 -52443 -29592
rect -52207 -29828 -52165 -29592
rect -52485 -29890 -52165 -29828
rect -51485 -29272 -51165 -29210
rect -51485 -29508 -51443 -29272
rect -51207 -29508 -51165 -29272
rect -51485 -29592 -51165 -29508
rect -51485 -29828 -51443 -29592
rect -51207 -29828 -51165 -29592
rect -51485 -29890 -51165 -29828
rect -50485 -29272 -50165 -29210
rect -50485 -29508 -50443 -29272
rect -50207 -29508 -50165 -29272
rect -50485 -29592 -50165 -29508
rect -50485 -29828 -50443 -29592
rect -50207 -29828 -50165 -29592
rect -50485 -29890 -50165 -29828
rect -49485 -29272 -49165 -29210
rect -49485 -29508 -49443 -29272
rect -49207 -29508 -49165 -29272
rect -49485 -29592 -49165 -29508
rect -49485 -29828 -49443 -29592
rect -49207 -29828 -49165 -29592
rect -49485 -29890 -49165 -29828
tri -41465 -29890 -40785 -29210 se
rect -40785 -29890 -33465 -29210
tri -33465 -29890 -32785 -29210 nw
rect -74825 -29932 -48825 -29890
rect -74825 -30168 -74783 -29932
rect -74547 -30168 -74443 -29932
rect -74207 -30168 -74103 -29932
rect -73867 -30168 -73783 -29932
rect -73547 -30168 -73443 -29932
rect -73207 -30168 -73103 -29932
rect -72867 -30168 -72783 -29932
rect -72547 -30168 -72443 -29932
rect -72207 -30168 -72103 -29932
rect -71867 -30168 -71783 -29932
rect -71547 -30168 -71443 -29932
rect -71207 -30168 -71103 -29932
rect -70867 -30168 -70783 -29932
rect -70547 -30168 -70443 -29932
rect -70207 -30168 -70103 -29932
rect -69867 -30168 -69783 -29932
rect -69547 -30168 -69443 -29932
rect -69207 -30168 -69103 -29932
rect -68867 -30168 -68783 -29932
rect -68547 -30168 -68443 -29932
rect -68207 -30168 -68103 -29932
rect -67867 -30168 -67783 -29932
rect -67547 -30168 -67443 -29932
rect -67207 -30168 -67103 -29932
rect -66867 -30168 -66783 -29932
rect -66547 -30168 -66443 -29932
rect -66207 -30168 -66103 -29932
rect -65867 -30168 -65783 -29932
rect -65547 -30168 -65443 -29932
rect -65207 -30168 -65103 -29932
rect -64867 -30168 -64783 -29932
rect -64547 -30168 -64443 -29932
rect -64207 -30168 -64103 -29932
rect -63867 -30168 -63783 -29932
rect -63547 -30168 -63443 -29932
rect -63207 -30168 -63103 -29932
rect -62867 -30168 -62783 -29932
rect -62547 -30168 -62443 -29932
rect -62207 -30168 -62103 -29932
rect -61867 -30168 -61783 -29932
rect -61547 -30168 -61443 -29932
rect -61207 -30168 -61103 -29932
rect -60867 -30168 -60783 -29932
rect -60547 -30168 -60443 -29932
rect -60207 -30168 -60103 -29932
rect -59867 -30168 -59783 -29932
rect -59547 -30168 -59443 -29932
rect -59207 -30168 -59103 -29932
rect -58867 -30168 -58783 -29932
rect -58547 -30168 -58443 -29932
rect -58207 -30168 -58103 -29932
rect -57867 -30168 -57783 -29932
rect -57547 -30168 -57443 -29932
rect -57207 -30168 -57103 -29932
rect -56867 -30168 -56783 -29932
rect -56547 -30168 -56443 -29932
rect -56207 -30168 -56103 -29932
rect -55867 -30168 -55783 -29932
rect -55547 -30168 -55443 -29932
rect -55207 -30168 -55103 -29932
rect -54867 -30168 -54783 -29932
rect -54547 -30168 -54443 -29932
rect -54207 -30168 -54103 -29932
rect -53867 -30168 -53783 -29932
rect -53547 -30168 -53443 -29932
rect -53207 -30168 -53103 -29932
rect -52867 -30168 -52783 -29932
rect -52547 -30168 -52443 -29932
rect -52207 -30168 -52103 -29932
rect -51867 -30168 -51783 -29932
rect -51547 -30168 -51443 -29932
rect -51207 -30168 -51103 -29932
rect -50867 -30168 -50783 -29932
rect -50547 -30168 -50443 -29932
rect -50207 -30168 -50103 -29932
rect -49867 -30168 -49783 -29932
rect -49547 -30168 -49443 -29932
rect -49207 -30168 -49103 -29932
rect -48867 -30168 -48825 -29932
rect -74825 -30210 -48825 -30168
tri -41785 -30210 -41465 -29890 se
rect -41465 -30210 -33785 -29890
tri -33785 -30210 -33465 -29890 nw
rect -74485 -30272 -74165 -30210
rect -74485 -30508 -74443 -30272
rect -74207 -30508 -74165 -30272
rect -74485 -30592 -74165 -30508
rect -74485 -30828 -74443 -30592
rect -74207 -30828 -74165 -30592
rect -74485 -30890 -74165 -30828
rect -73485 -30272 -73165 -30210
rect -73485 -30508 -73443 -30272
rect -73207 -30508 -73165 -30272
rect -73485 -30592 -73165 -30508
rect -73485 -30828 -73443 -30592
rect -73207 -30828 -73165 -30592
rect -73485 -30890 -73165 -30828
rect -72485 -30272 -72165 -30210
rect -72485 -30508 -72443 -30272
rect -72207 -30508 -72165 -30272
rect -72485 -30592 -72165 -30508
rect -72485 -30828 -72443 -30592
rect -72207 -30828 -72165 -30592
rect -72485 -30890 -72165 -30828
rect -71485 -30272 -71165 -30210
rect -71485 -30508 -71443 -30272
rect -71207 -30508 -71165 -30272
rect -71485 -30592 -71165 -30508
rect -71485 -30828 -71443 -30592
rect -71207 -30828 -71165 -30592
rect -71485 -30890 -71165 -30828
rect -70485 -30272 -70165 -30210
rect -70485 -30508 -70443 -30272
rect -70207 -30508 -70165 -30272
rect -70485 -30592 -70165 -30508
rect -70485 -30828 -70443 -30592
rect -70207 -30828 -70165 -30592
rect -70485 -30890 -70165 -30828
rect -69485 -30272 -69165 -30210
rect -69485 -30508 -69443 -30272
rect -69207 -30508 -69165 -30272
rect -69485 -30592 -69165 -30508
rect -69485 -30828 -69443 -30592
rect -69207 -30828 -69165 -30592
rect -69485 -30890 -69165 -30828
rect -68485 -30272 -68165 -30210
rect -68485 -30508 -68443 -30272
rect -68207 -30508 -68165 -30272
rect -68485 -30592 -68165 -30508
rect -68485 -30828 -68443 -30592
rect -68207 -30828 -68165 -30592
rect -68485 -30890 -68165 -30828
rect -67485 -30272 -67165 -30210
rect -67485 -30508 -67443 -30272
rect -67207 -30508 -67165 -30272
rect -67485 -30592 -67165 -30508
rect -67485 -30828 -67443 -30592
rect -67207 -30828 -67165 -30592
rect -67485 -30890 -67165 -30828
rect -66485 -30272 -66165 -30210
rect -66485 -30508 -66443 -30272
rect -66207 -30508 -66165 -30272
rect -66485 -30592 -66165 -30508
rect -66485 -30828 -66443 -30592
rect -66207 -30828 -66165 -30592
rect -66485 -30890 -66165 -30828
rect -65485 -30272 -65165 -30210
rect -65485 -30508 -65443 -30272
rect -65207 -30508 -65165 -30272
rect -65485 -30592 -65165 -30508
rect -65485 -30828 -65443 -30592
rect -65207 -30828 -65165 -30592
rect -65485 -30890 -65165 -30828
rect -64485 -30272 -64165 -30210
rect -64485 -30508 -64443 -30272
rect -64207 -30508 -64165 -30272
rect -64485 -30592 -64165 -30508
rect -64485 -30828 -64443 -30592
rect -64207 -30828 -64165 -30592
rect -64485 -30890 -64165 -30828
rect -63485 -30272 -63165 -30210
rect -63485 -30508 -63443 -30272
rect -63207 -30508 -63165 -30272
rect -63485 -30592 -63165 -30508
rect -63485 -30828 -63443 -30592
rect -63207 -30828 -63165 -30592
rect -63485 -30890 -63165 -30828
rect -62485 -30272 -62165 -30210
rect -62485 -30508 -62443 -30272
rect -62207 -30508 -62165 -30272
rect -62485 -30592 -62165 -30508
rect -62485 -30828 -62443 -30592
rect -62207 -30828 -62165 -30592
rect -62485 -30890 -62165 -30828
rect -61485 -30272 -61165 -30210
rect -61485 -30508 -61443 -30272
rect -61207 -30508 -61165 -30272
rect -61485 -30592 -61165 -30508
rect -61485 -30828 -61443 -30592
rect -61207 -30828 -61165 -30592
rect -61485 -30890 -61165 -30828
rect -60485 -30272 -60165 -30210
rect -60485 -30508 -60443 -30272
rect -60207 -30508 -60165 -30272
rect -60485 -30592 -60165 -30508
rect -60485 -30828 -60443 -30592
rect -60207 -30828 -60165 -30592
rect -60485 -30890 -60165 -30828
rect -59485 -30272 -59165 -30210
rect -59485 -30508 -59443 -30272
rect -59207 -30508 -59165 -30272
rect -59485 -30592 -59165 -30508
rect -59485 -30828 -59443 -30592
rect -59207 -30828 -59165 -30592
rect -59485 -30890 -59165 -30828
rect -58485 -30272 -58165 -30210
rect -58485 -30508 -58443 -30272
rect -58207 -30508 -58165 -30272
rect -58485 -30592 -58165 -30508
rect -58485 -30828 -58443 -30592
rect -58207 -30828 -58165 -30592
rect -58485 -30890 -58165 -30828
rect -57485 -30272 -57165 -30210
rect -57485 -30508 -57443 -30272
rect -57207 -30508 -57165 -30272
rect -57485 -30592 -57165 -30508
rect -57485 -30828 -57443 -30592
rect -57207 -30828 -57165 -30592
rect -57485 -30890 -57165 -30828
rect -56485 -30272 -56165 -30210
rect -56485 -30508 -56443 -30272
rect -56207 -30508 -56165 -30272
rect -56485 -30592 -56165 -30508
rect -56485 -30828 -56443 -30592
rect -56207 -30828 -56165 -30592
rect -56485 -30890 -56165 -30828
rect -55485 -30272 -55165 -30210
rect -55485 -30508 -55443 -30272
rect -55207 -30508 -55165 -30272
rect -55485 -30592 -55165 -30508
rect -55485 -30828 -55443 -30592
rect -55207 -30828 -55165 -30592
rect -55485 -30890 -55165 -30828
rect -54485 -30272 -54165 -30210
rect -54485 -30508 -54443 -30272
rect -54207 -30508 -54165 -30272
rect -54485 -30592 -54165 -30508
rect -54485 -30828 -54443 -30592
rect -54207 -30828 -54165 -30592
rect -54485 -30890 -54165 -30828
rect -53485 -30272 -53165 -30210
rect -53485 -30508 -53443 -30272
rect -53207 -30508 -53165 -30272
rect -53485 -30592 -53165 -30508
rect -53485 -30828 -53443 -30592
rect -53207 -30828 -53165 -30592
rect -53485 -30890 -53165 -30828
rect -52485 -30272 -52165 -30210
rect -52485 -30508 -52443 -30272
rect -52207 -30508 -52165 -30272
rect -52485 -30592 -52165 -30508
rect -52485 -30828 -52443 -30592
rect -52207 -30828 -52165 -30592
rect -52485 -30890 -52165 -30828
rect -51485 -30272 -51165 -30210
rect -51485 -30508 -51443 -30272
rect -51207 -30508 -51165 -30272
rect -51485 -30592 -51165 -30508
rect -51485 -30828 -51443 -30592
rect -51207 -30828 -51165 -30592
rect -51485 -30890 -51165 -30828
rect -50485 -30272 -50165 -30210
rect -50485 -30508 -50443 -30272
rect -50207 -30508 -50165 -30272
rect -50485 -30592 -50165 -30508
rect -50485 -30828 -50443 -30592
rect -50207 -30828 -50165 -30592
rect -50485 -30890 -50165 -30828
rect -49485 -30272 -49165 -30210
rect -49485 -30508 -49443 -30272
rect -49207 -30508 -49165 -30272
rect -49485 -30592 -49165 -30508
rect -49485 -30828 -49443 -30592
rect -49207 -30828 -49165 -30592
rect -49485 -30890 -49165 -30828
tri -42465 -30890 -41785 -30210 se
rect -41785 -30890 -34465 -30210
tri -34465 -30890 -33785 -30210 nw
rect -74825 -30932 -48825 -30890
rect -74825 -31168 -74783 -30932
rect -74547 -31168 -74443 -30932
rect -74207 -31168 -74103 -30932
rect -73867 -31168 -73783 -30932
rect -73547 -31168 -73443 -30932
rect -73207 -31168 -73103 -30932
rect -72867 -31168 -72783 -30932
rect -72547 -31168 -72443 -30932
rect -72207 -31168 -72103 -30932
rect -71867 -31168 -71783 -30932
rect -71547 -31168 -71443 -30932
rect -71207 -31168 -71103 -30932
rect -70867 -31168 -70783 -30932
rect -70547 -31168 -70443 -30932
rect -70207 -31168 -70103 -30932
rect -69867 -31168 -69783 -30932
rect -69547 -31168 -69443 -30932
rect -69207 -31168 -69103 -30932
rect -68867 -31168 -68783 -30932
rect -68547 -31168 -68443 -30932
rect -68207 -31168 -68103 -30932
rect -67867 -31168 -67783 -30932
rect -67547 -31168 -67443 -30932
rect -67207 -31168 -67103 -30932
rect -66867 -31168 -66783 -30932
rect -66547 -31168 -66443 -30932
rect -66207 -31168 -66103 -30932
rect -65867 -31168 -65783 -30932
rect -65547 -31168 -65443 -30932
rect -65207 -31168 -65103 -30932
rect -64867 -31168 -64783 -30932
rect -64547 -31168 -64443 -30932
rect -64207 -31168 -64103 -30932
rect -63867 -31168 -63783 -30932
rect -63547 -31168 -63443 -30932
rect -63207 -31168 -63103 -30932
rect -62867 -31168 -62783 -30932
rect -62547 -31168 -62443 -30932
rect -62207 -31168 -62103 -30932
rect -61867 -31168 -61783 -30932
rect -61547 -31168 -61443 -30932
rect -61207 -31168 -61103 -30932
rect -60867 -31168 -60783 -30932
rect -60547 -31168 -60443 -30932
rect -60207 -31168 -60103 -30932
rect -59867 -31168 -59783 -30932
rect -59547 -31168 -59443 -30932
rect -59207 -31168 -59103 -30932
rect -58867 -31168 -58783 -30932
rect -58547 -31168 -58443 -30932
rect -58207 -31168 -58103 -30932
rect -57867 -31168 -57783 -30932
rect -57547 -31168 -57443 -30932
rect -57207 -31168 -57103 -30932
rect -56867 -31168 -56783 -30932
rect -56547 -31168 -56443 -30932
rect -56207 -31168 -56103 -30932
rect -55867 -31168 -55783 -30932
rect -55547 -31168 -55443 -30932
rect -55207 -31168 -55103 -30932
rect -54867 -31168 -54783 -30932
rect -54547 -31168 -54443 -30932
rect -54207 -31168 -54103 -30932
rect -53867 -31168 -53783 -30932
rect -53547 -31168 -53443 -30932
rect -53207 -31168 -53103 -30932
rect -52867 -31168 -52783 -30932
rect -52547 -31168 -52443 -30932
rect -52207 -31168 -52103 -30932
rect -51867 -31168 -51783 -30932
rect -51547 -31168 -51443 -30932
rect -51207 -31168 -51103 -30932
rect -50867 -31168 -50783 -30932
rect -50547 -31168 -50443 -30932
rect -50207 -31168 -50103 -30932
rect -49867 -31168 -49783 -30932
rect -49547 -31168 -49443 -30932
rect -49207 -31168 -49103 -30932
rect -48867 -31168 -48825 -30932
rect -74825 -31210 -48825 -31168
tri -42785 -31210 -42465 -30890 se
rect -42465 -31210 -34785 -30890
tri -34785 -31210 -34465 -30890 nw
rect -74485 -31272 -74165 -31210
rect -74485 -31508 -74443 -31272
rect -74207 -31508 -74165 -31272
rect -74485 -31592 -74165 -31508
rect -74485 -31828 -74443 -31592
rect -74207 -31828 -74165 -31592
rect -74485 -31890 -74165 -31828
rect -73485 -31272 -73165 -31210
rect -73485 -31508 -73443 -31272
rect -73207 -31508 -73165 -31272
rect -73485 -31592 -73165 -31508
rect -73485 -31828 -73443 -31592
rect -73207 -31828 -73165 -31592
rect -73485 -31890 -73165 -31828
rect -72485 -31272 -72165 -31210
rect -72485 -31508 -72443 -31272
rect -72207 -31508 -72165 -31272
rect -72485 -31592 -72165 -31508
rect -72485 -31828 -72443 -31592
rect -72207 -31828 -72165 -31592
rect -72485 -31890 -72165 -31828
rect -71485 -31272 -71165 -31210
rect -71485 -31508 -71443 -31272
rect -71207 -31508 -71165 -31272
rect -71485 -31592 -71165 -31508
rect -71485 -31828 -71443 -31592
rect -71207 -31828 -71165 -31592
rect -71485 -31890 -71165 -31828
rect -70485 -31272 -70165 -31210
rect -70485 -31508 -70443 -31272
rect -70207 -31508 -70165 -31272
rect -70485 -31592 -70165 -31508
rect -70485 -31828 -70443 -31592
rect -70207 -31828 -70165 -31592
rect -70485 -31890 -70165 -31828
rect -69485 -31272 -69165 -31210
rect -69485 -31508 -69443 -31272
rect -69207 -31508 -69165 -31272
rect -69485 -31592 -69165 -31508
rect -69485 -31828 -69443 -31592
rect -69207 -31828 -69165 -31592
rect -69485 -31890 -69165 -31828
rect -68485 -31272 -68165 -31210
rect -68485 -31508 -68443 -31272
rect -68207 -31508 -68165 -31272
rect -68485 -31592 -68165 -31508
rect -68485 -31828 -68443 -31592
rect -68207 -31828 -68165 -31592
rect -68485 -31890 -68165 -31828
rect -67485 -31272 -67165 -31210
rect -67485 -31508 -67443 -31272
rect -67207 -31508 -67165 -31272
rect -67485 -31592 -67165 -31508
rect -67485 -31828 -67443 -31592
rect -67207 -31828 -67165 -31592
rect -67485 -31890 -67165 -31828
rect -66485 -31272 -66165 -31210
rect -66485 -31508 -66443 -31272
rect -66207 -31508 -66165 -31272
rect -66485 -31592 -66165 -31508
rect -66485 -31828 -66443 -31592
rect -66207 -31828 -66165 -31592
rect -66485 -31890 -66165 -31828
rect -65485 -31272 -65165 -31210
rect -65485 -31508 -65443 -31272
rect -65207 -31508 -65165 -31272
rect -65485 -31592 -65165 -31508
rect -65485 -31828 -65443 -31592
rect -65207 -31828 -65165 -31592
rect -65485 -31890 -65165 -31828
rect -64485 -31272 -64165 -31210
rect -64485 -31508 -64443 -31272
rect -64207 -31508 -64165 -31272
rect -64485 -31592 -64165 -31508
rect -64485 -31828 -64443 -31592
rect -64207 -31828 -64165 -31592
rect -64485 -31890 -64165 -31828
rect -63485 -31272 -63165 -31210
rect -63485 -31508 -63443 -31272
rect -63207 -31508 -63165 -31272
rect -63485 -31592 -63165 -31508
rect -63485 -31828 -63443 -31592
rect -63207 -31828 -63165 -31592
rect -63485 -31890 -63165 -31828
rect -62485 -31272 -62165 -31210
rect -62485 -31508 -62443 -31272
rect -62207 -31508 -62165 -31272
rect -62485 -31592 -62165 -31508
rect -62485 -31828 -62443 -31592
rect -62207 -31828 -62165 -31592
rect -62485 -31890 -62165 -31828
rect -61485 -31272 -61165 -31210
rect -61485 -31508 -61443 -31272
rect -61207 -31508 -61165 -31272
rect -61485 -31592 -61165 -31508
rect -61485 -31828 -61443 -31592
rect -61207 -31828 -61165 -31592
rect -61485 -31890 -61165 -31828
rect -60485 -31272 -60165 -31210
rect -60485 -31508 -60443 -31272
rect -60207 -31508 -60165 -31272
rect -60485 -31592 -60165 -31508
rect -60485 -31828 -60443 -31592
rect -60207 -31828 -60165 -31592
rect -60485 -31890 -60165 -31828
rect -59485 -31272 -59165 -31210
rect -59485 -31508 -59443 -31272
rect -59207 -31508 -59165 -31272
rect -59485 -31592 -59165 -31508
rect -59485 -31828 -59443 -31592
rect -59207 -31828 -59165 -31592
rect -59485 -31890 -59165 -31828
rect -58485 -31272 -58165 -31210
rect -58485 -31508 -58443 -31272
rect -58207 -31508 -58165 -31272
rect -58485 -31592 -58165 -31508
rect -58485 -31828 -58443 -31592
rect -58207 -31828 -58165 -31592
rect -58485 -31890 -58165 -31828
rect -57485 -31272 -57165 -31210
rect -57485 -31508 -57443 -31272
rect -57207 -31508 -57165 -31272
rect -57485 -31592 -57165 -31508
rect -57485 -31828 -57443 -31592
rect -57207 -31828 -57165 -31592
rect -57485 -31890 -57165 -31828
rect -56485 -31272 -56165 -31210
rect -56485 -31508 -56443 -31272
rect -56207 -31508 -56165 -31272
rect -56485 -31592 -56165 -31508
rect -56485 -31828 -56443 -31592
rect -56207 -31828 -56165 -31592
rect -56485 -31890 -56165 -31828
rect -55485 -31272 -55165 -31210
rect -55485 -31508 -55443 -31272
rect -55207 -31508 -55165 -31272
rect -55485 -31592 -55165 -31508
rect -55485 -31828 -55443 -31592
rect -55207 -31828 -55165 -31592
rect -55485 -31890 -55165 -31828
rect -54485 -31272 -54165 -31210
rect -54485 -31508 -54443 -31272
rect -54207 -31508 -54165 -31272
rect -54485 -31592 -54165 -31508
rect -54485 -31828 -54443 -31592
rect -54207 -31828 -54165 -31592
rect -54485 -31890 -54165 -31828
rect -53485 -31272 -53165 -31210
rect -53485 -31508 -53443 -31272
rect -53207 -31508 -53165 -31272
rect -53485 -31592 -53165 -31508
rect -53485 -31828 -53443 -31592
rect -53207 -31828 -53165 -31592
rect -53485 -31890 -53165 -31828
rect -52485 -31272 -52165 -31210
rect -52485 -31508 -52443 -31272
rect -52207 -31508 -52165 -31272
rect -52485 -31592 -52165 -31508
rect -52485 -31828 -52443 -31592
rect -52207 -31828 -52165 -31592
rect -52485 -31890 -52165 -31828
rect -51485 -31272 -51165 -31210
rect -51485 -31508 -51443 -31272
rect -51207 -31508 -51165 -31272
rect -51485 -31592 -51165 -31508
rect -51485 -31828 -51443 -31592
rect -51207 -31828 -51165 -31592
rect -51485 -31890 -51165 -31828
rect -50485 -31272 -50165 -31210
rect -50485 -31508 -50443 -31272
rect -50207 -31508 -50165 -31272
rect -50485 -31592 -50165 -31508
rect -50485 -31828 -50443 -31592
rect -50207 -31828 -50165 -31592
rect -50485 -31890 -50165 -31828
rect -49485 -31272 -49165 -31210
rect -49485 -31508 -49443 -31272
rect -49207 -31508 -49165 -31272
rect -49485 -31592 -49165 -31508
rect -49485 -31828 -49443 -31592
rect -49207 -31828 -49165 -31592
rect -49485 -31890 -49165 -31828
tri -43465 -31890 -42785 -31210 se
rect -42785 -31890 -35465 -31210
tri -35465 -31890 -34785 -31210 nw
rect -74825 -31932 -48825 -31890
rect -74825 -32168 -74783 -31932
rect -74547 -32168 -74443 -31932
rect -74207 -32168 -74103 -31932
rect -73867 -32168 -73783 -31932
rect -73547 -32168 -73443 -31932
rect -73207 -32168 -73103 -31932
rect -72867 -32168 -72783 -31932
rect -72547 -32168 -72443 -31932
rect -72207 -32168 -72103 -31932
rect -71867 -32168 -71783 -31932
rect -71547 -32168 -71443 -31932
rect -71207 -32168 -71103 -31932
rect -70867 -32168 -70783 -31932
rect -70547 -32168 -70443 -31932
rect -70207 -32168 -70103 -31932
rect -69867 -32168 -69783 -31932
rect -69547 -32168 -69443 -31932
rect -69207 -32168 -69103 -31932
rect -68867 -32168 -68783 -31932
rect -68547 -32168 -68443 -31932
rect -68207 -32168 -68103 -31932
rect -67867 -32168 -67783 -31932
rect -67547 -32168 -67443 -31932
rect -67207 -32168 -67103 -31932
rect -66867 -32168 -66783 -31932
rect -66547 -32168 -66443 -31932
rect -66207 -32168 -66103 -31932
rect -65867 -32168 -65783 -31932
rect -65547 -32168 -65443 -31932
rect -65207 -32168 -65103 -31932
rect -64867 -32168 -64783 -31932
rect -64547 -32168 -64443 -31932
rect -64207 -32168 -64103 -31932
rect -63867 -32168 -63783 -31932
rect -63547 -32168 -63443 -31932
rect -63207 -32168 -63103 -31932
rect -62867 -32168 -62783 -31932
rect -62547 -32168 -62443 -31932
rect -62207 -32168 -62103 -31932
rect -61867 -32168 -61783 -31932
rect -61547 -32168 -61443 -31932
rect -61207 -32168 -61103 -31932
rect -60867 -32168 -60783 -31932
rect -60547 -32168 -60443 -31932
rect -60207 -32168 -60103 -31932
rect -59867 -32168 -59783 -31932
rect -59547 -32168 -59443 -31932
rect -59207 -32168 -59103 -31932
rect -58867 -32168 -58783 -31932
rect -58547 -32168 -58443 -31932
rect -58207 -32168 -58103 -31932
rect -57867 -32168 -57783 -31932
rect -57547 -32168 -57443 -31932
rect -57207 -32168 -57103 -31932
rect -56867 -32168 -56783 -31932
rect -56547 -32168 -56443 -31932
rect -56207 -32168 -56103 -31932
rect -55867 -32168 -55783 -31932
rect -55547 -32168 -55443 -31932
rect -55207 -32168 -55103 -31932
rect -54867 -32168 -54783 -31932
rect -54547 -32168 -54443 -31932
rect -54207 -32168 -54103 -31932
rect -53867 -32168 -53783 -31932
rect -53547 -32168 -53443 -31932
rect -53207 -32168 -53103 -31932
rect -52867 -32168 -52783 -31932
rect -52547 -32168 -52443 -31932
rect -52207 -32168 -52103 -31932
rect -51867 -32168 -51783 -31932
rect -51547 -32168 -51443 -31932
rect -51207 -32168 -51103 -31932
rect -50867 -32168 -50783 -31932
rect -50547 -32168 -50443 -31932
rect -50207 -32168 -50103 -31932
rect -49867 -32168 -49783 -31932
rect -49547 -32168 -49443 -31932
rect -49207 -32168 -49103 -31932
rect -48867 -32168 -48825 -31932
rect -74825 -32210 -48825 -32168
tri -43785 -32210 -43465 -31890 se
rect -43465 -32210 -35785 -31890
tri -35785 -32210 -35465 -31890 nw
rect -74485 -32272 -74165 -32210
rect -74485 -32508 -74443 -32272
rect -74207 -32508 -74165 -32272
rect -74485 -32592 -74165 -32508
rect -74485 -32828 -74443 -32592
rect -74207 -32828 -74165 -32592
rect -74485 -32890 -74165 -32828
rect -73485 -32272 -73165 -32210
rect -73485 -32508 -73443 -32272
rect -73207 -32508 -73165 -32272
rect -73485 -32592 -73165 -32508
rect -73485 -32828 -73443 -32592
rect -73207 -32828 -73165 -32592
rect -73485 -32890 -73165 -32828
rect -72485 -32272 -72165 -32210
rect -72485 -32508 -72443 -32272
rect -72207 -32508 -72165 -32272
rect -72485 -32592 -72165 -32508
rect -72485 -32828 -72443 -32592
rect -72207 -32828 -72165 -32592
rect -72485 -32890 -72165 -32828
rect -71485 -32272 -71165 -32210
rect -71485 -32508 -71443 -32272
rect -71207 -32508 -71165 -32272
rect -71485 -32592 -71165 -32508
rect -71485 -32828 -71443 -32592
rect -71207 -32828 -71165 -32592
rect -71485 -32890 -71165 -32828
rect -70485 -32272 -70165 -32210
rect -70485 -32508 -70443 -32272
rect -70207 -32508 -70165 -32272
rect -70485 -32592 -70165 -32508
rect -70485 -32828 -70443 -32592
rect -70207 -32828 -70165 -32592
rect -70485 -32890 -70165 -32828
rect -69485 -32272 -69165 -32210
rect -69485 -32508 -69443 -32272
rect -69207 -32508 -69165 -32272
rect -69485 -32592 -69165 -32508
rect -69485 -32828 -69443 -32592
rect -69207 -32828 -69165 -32592
rect -69485 -32890 -69165 -32828
rect -68485 -32272 -68165 -32210
rect -68485 -32508 -68443 -32272
rect -68207 -32508 -68165 -32272
rect -68485 -32592 -68165 -32508
rect -68485 -32828 -68443 -32592
rect -68207 -32828 -68165 -32592
rect -68485 -32890 -68165 -32828
rect -67485 -32272 -67165 -32210
rect -67485 -32508 -67443 -32272
rect -67207 -32508 -67165 -32272
rect -67485 -32592 -67165 -32508
rect -67485 -32828 -67443 -32592
rect -67207 -32828 -67165 -32592
rect -67485 -32890 -67165 -32828
rect -66485 -32272 -66165 -32210
rect -66485 -32508 -66443 -32272
rect -66207 -32508 -66165 -32272
rect -66485 -32592 -66165 -32508
rect -66485 -32828 -66443 -32592
rect -66207 -32828 -66165 -32592
rect -66485 -32890 -66165 -32828
rect -65485 -32272 -65165 -32210
rect -65485 -32508 -65443 -32272
rect -65207 -32508 -65165 -32272
rect -65485 -32592 -65165 -32508
rect -65485 -32828 -65443 -32592
rect -65207 -32828 -65165 -32592
rect -65485 -32890 -65165 -32828
rect -64485 -32272 -64165 -32210
rect -64485 -32508 -64443 -32272
rect -64207 -32508 -64165 -32272
rect -64485 -32592 -64165 -32508
rect -64485 -32828 -64443 -32592
rect -64207 -32828 -64165 -32592
rect -64485 -32890 -64165 -32828
rect -63485 -32272 -63165 -32210
rect -63485 -32508 -63443 -32272
rect -63207 -32508 -63165 -32272
rect -63485 -32592 -63165 -32508
rect -63485 -32828 -63443 -32592
rect -63207 -32828 -63165 -32592
rect -63485 -32890 -63165 -32828
rect -62485 -32272 -62165 -32210
rect -62485 -32508 -62443 -32272
rect -62207 -32508 -62165 -32272
rect -62485 -32592 -62165 -32508
rect -62485 -32828 -62443 -32592
rect -62207 -32828 -62165 -32592
rect -62485 -32890 -62165 -32828
rect -61485 -32272 -61165 -32210
rect -61485 -32508 -61443 -32272
rect -61207 -32508 -61165 -32272
rect -61485 -32592 -61165 -32508
rect -61485 -32828 -61443 -32592
rect -61207 -32828 -61165 -32592
rect -61485 -32890 -61165 -32828
rect -60485 -32272 -60165 -32210
rect -60485 -32508 -60443 -32272
rect -60207 -32508 -60165 -32272
rect -60485 -32592 -60165 -32508
rect -60485 -32828 -60443 -32592
rect -60207 -32828 -60165 -32592
rect -60485 -32890 -60165 -32828
rect -59485 -32272 -59165 -32210
rect -59485 -32508 -59443 -32272
rect -59207 -32508 -59165 -32272
rect -59485 -32592 -59165 -32508
rect -59485 -32828 -59443 -32592
rect -59207 -32828 -59165 -32592
rect -59485 -32890 -59165 -32828
rect -58485 -32272 -58165 -32210
rect -58485 -32508 -58443 -32272
rect -58207 -32508 -58165 -32272
rect -58485 -32592 -58165 -32508
rect -58485 -32828 -58443 -32592
rect -58207 -32828 -58165 -32592
rect -58485 -32890 -58165 -32828
rect -57485 -32272 -57165 -32210
rect -57485 -32508 -57443 -32272
rect -57207 -32508 -57165 -32272
rect -57485 -32592 -57165 -32508
rect -57485 -32828 -57443 -32592
rect -57207 -32828 -57165 -32592
rect -57485 -32890 -57165 -32828
rect -56485 -32272 -56165 -32210
rect -56485 -32508 -56443 -32272
rect -56207 -32508 -56165 -32272
rect -56485 -32592 -56165 -32508
rect -56485 -32828 -56443 -32592
rect -56207 -32828 -56165 -32592
rect -56485 -32890 -56165 -32828
rect -55485 -32272 -55165 -32210
rect -55485 -32508 -55443 -32272
rect -55207 -32508 -55165 -32272
rect -55485 -32592 -55165 -32508
rect -55485 -32828 -55443 -32592
rect -55207 -32828 -55165 -32592
rect -55485 -32890 -55165 -32828
rect -54485 -32272 -54165 -32210
rect -54485 -32508 -54443 -32272
rect -54207 -32508 -54165 -32272
rect -54485 -32592 -54165 -32508
rect -54485 -32828 -54443 -32592
rect -54207 -32828 -54165 -32592
rect -54485 -32890 -54165 -32828
rect -53485 -32272 -53165 -32210
rect -53485 -32508 -53443 -32272
rect -53207 -32508 -53165 -32272
rect -53485 -32592 -53165 -32508
rect -53485 -32828 -53443 -32592
rect -53207 -32828 -53165 -32592
rect -53485 -32890 -53165 -32828
rect -52485 -32272 -52165 -32210
rect -52485 -32508 -52443 -32272
rect -52207 -32508 -52165 -32272
rect -52485 -32592 -52165 -32508
rect -52485 -32828 -52443 -32592
rect -52207 -32828 -52165 -32592
rect -52485 -32890 -52165 -32828
rect -51485 -32272 -51165 -32210
rect -51485 -32508 -51443 -32272
rect -51207 -32508 -51165 -32272
rect -51485 -32592 -51165 -32508
rect -51485 -32828 -51443 -32592
rect -51207 -32828 -51165 -32592
rect -51485 -32890 -51165 -32828
rect -50485 -32272 -50165 -32210
rect -50485 -32508 -50443 -32272
rect -50207 -32508 -50165 -32272
rect -50485 -32592 -50165 -32508
rect -50485 -32828 -50443 -32592
rect -50207 -32828 -50165 -32592
rect -50485 -32890 -50165 -32828
rect -49485 -32272 -49165 -32210
rect -49485 -32508 -49443 -32272
rect -49207 -32508 -49165 -32272
rect -49485 -32592 -49165 -32508
tri -44125 -32550 -43785 -32210 se
rect -43785 -32550 -36125 -32210
tri -36125 -32550 -35785 -32210 nw
rect -22625 -32550 -17925 -2350
rect 20275 -2600 32275 -2350
tri 20275 -4600 22275 -2600 ne
rect 22275 -4600 30275 -2600
tri 30275 -4600 32275 -2600 nw
rect -12425 -7880 12275 -7850
tri 12275 -7880 12305 -7850 sw
rect -12425 -8012 12305 -7880
rect -12425 -8026 242 -8012
rect -12425 -13702 -12323 -8026
rect -11127 -13688 242 -8026
rect 1758 -13688 12305 -8012
rect -11127 -13702 12305 -13688
rect -12425 -13820 12305 -13702
tri 12305 -13820 18245 -7880 sw
rect -12425 -13830 18245 -13820
tri 18245 -13830 18255 -13820 sw
rect -12425 -13839 18255 -13830
tri 18255 -13839 18264 -13830 sw
rect -12425 -13850 18264 -13839
tri 18264 -13850 18275 -13839 sw
rect -12425 -23850 -6425 -13850
tri 10275 -15850 12275 -13850 ne
rect 12275 -15850 18275 -13850
tri 18275 -15850 20275 -13850 sw
tri 12275 -16000 12425 -15850 ne
rect 12425 -16000 20275 -15850
tri 20275 -16000 20425 -15850 sw
tri 12425 -16030 12455 -16000 ne
rect 12455 -16030 32275 -16000
tri 12455 -21850 18275 -16030 ne
rect 18275 -16082 32275 -16030
rect 18275 -21850 20392 -16082
tri 18275 -22550 18975 -21850 ne
rect 18975 -22550 20392 -21850
tri -6425 -23850 -5125 -22550 sw
tri 18975 -23850 20275 -22550 ne
rect -12425 -24550 -5125 -23850
tri -5125 -24550 -4425 -23850 sw
tri -12425 -25970 -11005 -24550 ne
rect -11005 -25970 -4425 -24550
tri -4425 -25970 -3005 -24550 sw
rect 20275 -25918 20392 -22550
rect 32148 -25918 32275 -16082
tri -11005 -26000 -10975 -25970 ne
rect -10975 -26000 -3005 -25970
tri -10975 -28550 -8425 -26000 ne
rect -8425 -28550 -3005 -26000
tri -8425 -28890 -8085 -28550 ne
rect -8085 -28890 -3005 -28550
tri -8085 -29210 -7765 -28890 ne
rect -7765 -29210 -3005 -28890
tri -7765 -29890 -7085 -29210 ne
rect -7085 -29890 -3005 -29210
tri -7085 -30210 -6765 -29890 ne
rect -6765 -30210 -3005 -29890
tri -6765 -30890 -6085 -30210 ne
rect -6085 -30890 -3005 -30210
tri -6085 -31210 -5765 -30890 ne
rect -5765 -31210 -3005 -30890
tri -5765 -31890 -5085 -31210 ne
rect -5085 -31890 -3005 -31210
tri -5085 -32210 -4765 -31890 ne
rect -4765 -32210 -3005 -31890
tri -4765 -32550 -4425 -32210 ne
rect -4425 -32550 -3005 -32210
tri -3005 -32550 3575 -25970 sw
rect 20275 -26000 32275 -25918
rect 8615 -28592 8935 -28550
rect 8615 -28828 8657 -28592
rect 8893 -28828 8935 -28592
rect 8615 -28890 8935 -28828
rect 9615 -28592 9935 -28550
rect 9615 -28828 9657 -28592
rect 9893 -28828 9935 -28592
rect 9615 -28890 9935 -28828
rect 10615 -28592 10935 -28550
rect 10615 -28828 10657 -28592
rect 10893 -28828 10935 -28592
rect 10615 -28890 10935 -28828
rect 11615 -28592 11935 -28550
rect 11615 -28828 11657 -28592
rect 11893 -28828 11935 -28592
rect 11615 -28890 11935 -28828
rect 12615 -28592 12935 -28550
rect 12615 -28828 12657 -28592
rect 12893 -28828 12935 -28592
rect 12615 -28890 12935 -28828
rect 13615 -28592 13935 -28550
rect 13615 -28828 13657 -28592
rect 13893 -28828 13935 -28592
rect 13615 -28890 13935 -28828
rect 14615 -28592 14935 -28550
rect 14615 -28828 14657 -28592
rect 14893 -28828 14935 -28592
rect 14615 -28890 14935 -28828
rect 15615 -28592 15935 -28550
rect 15615 -28828 15657 -28592
rect 15893 -28828 15935 -28592
rect 15615 -28890 15935 -28828
rect 16615 -28592 16935 -28550
rect 16615 -28828 16657 -28592
rect 16893 -28828 16935 -28592
rect 16615 -28890 16935 -28828
rect 17615 -28592 17935 -28550
rect 17615 -28828 17657 -28592
rect 17893 -28828 17935 -28592
rect 17615 -28890 17935 -28828
rect 18615 -28592 18935 -28550
rect 18615 -28828 18657 -28592
rect 18893 -28828 18935 -28592
rect 18615 -28890 18935 -28828
rect 19615 -28592 19935 -28550
rect 19615 -28828 19657 -28592
rect 19893 -28828 19935 -28592
rect 19615 -28890 19935 -28828
rect 20615 -28592 20935 -28550
rect 20615 -28828 20657 -28592
rect 20893 -28828 20935 -28592
rect 20615 -28890 20935 -28828
rect 21615 -28592 21935 -28550
rect 21615 -28828 21657 -28592
rect 21893 -28828 21935 -28592
rect 21615 -28890 21935 -28828
rect 22615 -28592 22935 -28550
rect 22615 -28828 22657 -28592
rect 22893 -28828 22935 -28592
rect 22615 -28890 22935 -28828
rect 23615 -28592 23935 -28550
rect 23615 -28828 23657 -28592
rect 23893 -28828 23935 -28592
rect 23615 -28890 23935 -28828
rect 24615 -28592 24935 -28550
rect 24615 -28828 24657 -28592
rect 24893 -28828 24935 -28592
rect 24615 -28890 24935 -28828
rect 25615 -28592 25935 -28550
rect 25615 -28828 25657 -28592
rect 25893 -28828 25935 -28592
rect 25615 -28890 25935 -28828
rect 26615 -28592 26935 -28550
rect 26615 -28828 26657 -28592
rect 26893 -28828 26935 -28592
rect 26615 -28890 26935 -28828
rect 27615 -28592 27935 -28550
rect 27615 -28828 27657 -28592
rect 27893 -28828 27935 -28592
rect 27615 -28890 27935 -28828
rect 28615 -28592 28935 -28550
rect 28615 -28828 28657 -28592
rect 28893 -28828 28935 -28592
rect 28615 -28890 28935 -28828
rect 29615 -28592 29935 -28550
rect 29615 -28828 29657 -28592
rect 29893 -28828 29935 -28592
rect 29615 -28890 29935 -28828
rect 30615 -28592 30935 -28550
rect 30615 -28828 30657 -28592
rect 30893 -28828 30935 -28592
rect 30615 -28890 30935 -28828
rect 31615 -28592 31935 -28550
rect 31615 -28828 31657 -28592
rect 31893 -28828 31935 -28592
rect 31615 -28890 31935 -28828
rect 32615 -28592 32935 -28550
rect 32615 -28828 32657 -28592
rect 32893 -28828 32935 -28592
rect 32615 -28890 32935 -28828
rect 33615 -28592 33935 -28550
rect 33615 -28828 33657 -28592
rect 33893 -28828 33935 -28592
rect 33615 -28890 33935 -28828
rect 8275 -28932 34275 -28890
rect 8275 -29168 8317 -28932
rect 8553 -29168 8657 -28932
rect 8893 -29168 8997 -28932
rect 9233 -29168 9317 -28932
rect 9553 -29168 9657 -28932
rect 9893 -29168 9997 -28932
rect 10233 -29168 10317 -28932
rect 10553 -29168 10657 -28932
rect 10893 -29168 10997 -28932
rect 11233 -29168 11317 -28932
rect 11553 -29168 11657 -28932
rect 11893 -29168 11997 -28932
rect 12233 -29168 12317 -28932
rect 12553 -29168 12657 -28932
rect 12893 -29168 12997 -28932
rect 13233 -29168 13317 -28932
rect 13553 -29168 13657 -28932
rect 13893 -29168 13997 -28932
rect 14233 -29168 14317 -28932
rect 14553 -29168 14657 -28932
rect 14893 -29168 14997 -28932
rect 15233 -29168 15317 -28932
rect 15553 -29168 15657 -28932
rect 15893 -29168 15997 -28932
rect 16233 -29168 16317 -28932
rect 16553 -29168 16657 -28932
rect 16893 -29168 16997 -28932
rect 17233 -29168 17317 -28932
rect 17553 -29168 17657 -28932
rect 17893 -29168 17997 -28932
rect 18233 -29168 18317 -28932
rect 18553 -29168 18657 -28932
rect 18893 -29168 18997 -28932
rect 19233 -29168 19317 -28932
rect 19553 -29168 19657 -28932
rect 19893 -29168 19997 -28932
rect 20233 -29168 20317 -28932
rect 20553 -29168 20657 -28932
rect 20893 -29168 20997 -28932
rect 21233 -29168 21317 -28932
rect 21553 -29168 21657 -28932
rect 21893 -29168 21997 -28932
rect 22233 -29168 22317 -28932
rect 22553 -29168 22657 -28932
rect 22893 -29168 22997 -28932
rect 23233 -29168 23317 -28932
rect 23553 -29168 23657 -28932
rect 23893 -29168 23997 -28932
rect 24233 -29168 24317 -28932
rect 24553 -29168 24657 -28932
rect 24893 -29168 24997 -28932
rect 25233 -29168 25317 -28932
rect 25553 -29168 25657 -28932
rect 25893 -29168 25997 -28932
rect 26233 -29168 26317 -28932
rect 26553 -29168 26657 -28932
rect 26893 -29168 26997 -28932
rect 27233 -29168 27317 -28932
rect 27553 -29168 27657 -28932
rect 27893 -29168 27997 -28932
rect 28233 -29168 28317 -28932
rect 28553 -29168 28657 -28932
rect 28893 -29168 28997 -28932
rect 29233 -29168 29317 -28932
rect 29553 -29168 29657 -28932
rect 29893 -29168 29997 -28932
rect 30233 -29168 30317 -28932
rect 30553 -29168 30657 -28932
rect 30893 -29168 30997 -28932
rect 31233 -29168 31317 -28932
rect 31553 -29168 31657 -28932
rect 31893 -29168 31997 -28932
rect 32233 -29168 32317 -28932
rect 32553 -29168 32657 -28932
rect 32893 -29168 32997 -28932
rect 33233 -29168 33317 -28932
rect 33553 -29168 33657 -28932
rect 33893 -29168 33997 -28932
rect 34233 -29168 34275 -28932
rect 8275 -29210 34275 -29168
rect 8615 -29272 8935 -29210
rect 8615 -29508 8657 -29272
rect 8893 -29508 8935 -29272
rect 8615 -29592 8935 -29508
rect 8615 -29828 8657 -29592
rect 8893 -29828 8935 -29592
rect 8615 -29890 8935 -29828
rect 9615 -29272 9935 -29210
rect 9615 -29508 9657 -29272
rect 9893 -29508 9935 -29272
rect 9615 -29592 9935 -29508
rect 9615 -29828 9657 -29592
rect 9893 -29828 9935 -29592
rect 9615 -29890 9935 -29828
rect 10615 -29272 10935 -29210
rect 10615 -29508 10657 -29272
rect 10893 -29508 10935 -29272
rect 10615 -29592 10935 -29508
rect 10615 -29828 10657 -29592
rect 10893 -29828 10935 -29592
rect 10615 -29890 10935 -29828
rect 11615 -29272 11935 -29210
rect 11615 -29508 11657 -29272
rect 11893 -29508 11935 -29272
rect 11615 -29592 11935 -29508
rect 11615 -29828 11657 -29592
rect 11893 -29828 11935 -29592
rect 11615 -29890 11935 -29828
rect 12615 -29272 12935 -29210
rect 12615 -29508 12657 -29272
rect 12893 -29508 12935 -29272
rect 12615 -29592 12935 -29508
rect 12615 -29828 12657 -29592
rect 12893 -29828 12935 -29592
rect 12615 -29890 12935 -29828
rect 13615 -29272 13935 -29210
rect 13615 -29508 13657 -29272
rect 13893 -29508 13935 -29272
rect 13615 -29592 13935 -29508
rect 13615 -29828 13657 -29592
rect 13893 -29828 13935 -29592
rect 13615 -29890 13935 -29828
rect 14615 -29272 14935 -29210
rect 14615 -29508 14657 -29272
rect 14893 -29508 14935 -29272
rect 14615 -29592 14935 -29508
rect 14615 -29828 14657 -29592
rect 14893 -29828 14935 -29592
rect 14615 -29890 14935 -29828
rect 15615 -29272 15935 -29210
rect 15615 -29508 15657 -29272
rect 15893 -29508 15935 -29272
rect 15615 -29592 15935 -29508
rect 15615 -29828 15657 -29592
rect 15893 -29828 15935 -29592
rect 15615 -29890 15935 -29828
rect 16615 -29272 16935 -29210
rect 16615 -29508 16657 -29272
rect 16893 -29508 16935 -29272
rect 16615 -29592 16935 -29508
rect 16615 -29828 16657 -29592
rect 16893 -29828 16935 -29592
rect 16615 -29890 16935 -29828
rect 17615 -29272 17935 -29210
rect 17615 -29508 17657 -29272
rect 17893 -29508 17935 -29272
rect 17615 -29592 17935 -29508
rect 17615 -29828 17657 -29592
rect 17893 -29828 17935 -29592
rect 17615 -29890 17935 -29828
rect 18615 -29272 18935 -29210
rect 18615 -29508 18657 -29272
rect 18893 -29508 18935 -29272
rect 18615 -29592 18935 -29508
rect 18615 -29828 18657 -29592
rect 18893 -29828 18935 -29592
rect 18615 -29890 18935 -29828
rect 19615 -29272 19935 -29210
rect 19615 -29508 19657 -29272
rect 19893 -29508 19935 -29272
rect 19615 -29592 19935 -29508
rect 19615 -29828 19657 -29592
rect 19893 -29828 19935 -29592
rect 19615 -29890 19935 -29828
rect 20615 -29272 20935 -29210
rect 20615 -29508 20657 -29272
rect 20893 -29508 20935 -29272
rect 20615 -29592 20935 -29508
rect 20615 -29828 20657 -29592
rect 20893 -29828 20935 -29592
rect 20615 -29890 20935 -29828
rect 21615 -29272 21935 -29210
rect 21615 -29508 21657 -29272
rect 21893 -29508 21935 -29272
rect 21615 -29592 21935 -29508
rect 21615 -29828 21657 -29592
rect 21893 -29828 21935 -29592
rect 21615 -29890 21935 -29828
rect 22615 -29272 22935 -29210
rect 22615 -29508 22657 -29272
rect 22893 -29508 22935 -29272
rect 22615 -29592 22935 -29508
rect 22615 -29828 22657 -29592
rect 22893 -29828 22935 -29592
rect 22615 -29890 22935 -29828
rect 23615 -29272 23935 -29210
rect 23615 -29508 23657 -29272
rect 23893 -29508 23935 -29272
rect 23615 -29592 23935 -29508
rect 23615 -29828 23657 -29592
rect 23893 -29828 23935 -29592
rect 23615 -29890 23935 -29828
rect 24615 -29272 24935 -29210
rect 24615 -29508 24657 -29272
rect 24893 -29508 24935 -29272
rect 24615 -29592 24935 -29508
rect 24615 -29828 24657 -29592
rect 24893 -29828 24935 -29592
rect 24615 -29890 24935 -29828
rect 25615 -29272 25935 -29210
rect 25615 -29508 25657 -29272
rect 25893 -29508 25935 -29272
rect 25615 -29592 25935 -29508
rect 25615 -29828 25657 -29592
rect 25893 -29828 25935 -29592
rect 25615 -29890 25935 -29828
rect 26615 -29272 26935 -29210
rect 26615 -29508 26657 -29272
rect 26893 -29508 26935 -29272
rect 26615 -29592 26935 -29508
rect 26615 -29828 26657 -29592
rect 26893 -29828 26935 -29592
rect 26615 -29890 26935 -29828
rect 27615 -29272 27935 -29210
rect 27615 -29508 27657 -29272
rect 27893 -29508 27935 -29272
rect 27615 -29592 27935 -29508
rect 27615 -29828 27657 -29592
rect 27893 -29828 27935 -29592
rect 27615 -29890 27935 -29828
rect 28615 -29272 28935 -29210
rect 28615 -29508 28657 -29272
rect 28893 -29508 28935 -29272
rect 28615 -29592 28935 -29508
rect 28615 -29828 28657 -29592
rect 28893 -29828 28935 -29592
rect 28615 -29890 28935 -29828
rect 29615 -29272 29935 -29210
rect 29615 -29508 29657 -29272
rect 29893 -29508 29935 -29272
rect 29615 -29592 29935 -29508
rect 29615 -29828 29657 -29592
rect 29893 -29828 29935 -29592
rect 29615 -29890 29935 -29828
rect 30615 -29272 30935 -29210
rect 30615 -29508 30657 -29272
rect 30893 -29508 30935 -29272
rect 30615 -29592 30935 -29508
rect 30615 -29828 30657 -29592
rect 30893 -29828 30935 -29592
rect 30615 -29890 30935 -29828
rect 31615 -29272 31935 -29210
rect 31615 -29508 31657 -29272
rect 31893 -29508 31935 -29272
rect 31615 -29592 31935 -29508
rect 31615 -29828 31657 -29592
rect 31893 -29828 31935 -29592
rect 31615 -29890 31935 -29828
rect 32615 -29272 32935 -29210
rect 32615 -29508 32657 -29272
rect 32893 -29508 32935 -29272
rect 32615 -29592 32935 -29508
rect 32615 -29828 32657 -29592
rect 32893 -29828 32935 -29592
rect 32615 -29890 32935 -29828
rect 33615 -29272 33935 -29210
rect 33615 -29508 33657 -29272
rect 33893 -29508 33935 -29272
rect 33615 -29592 33935 -29508
rect 33615 -29828 33657 -29592
rect 33893 -29828 33935 -29592
rect 33615 -29890 33935 -29828
rect 8275 -29932 34275 -29890
rect 8275 -30168 8317 -29932
rect 8553 -30168 8657 -29932
rect 8893 -30168 8997 -29932
rect 9233 -30168 9317 -29932
rect 9553 -30168 9657 -29932
rect 9893 -30168 9997 -29932
rect 10233 -30168 10317 -29932
rect 10553 -30168 10657 -29932
rect 10893 -30168 10997 -29932
rect 11233 -30168 11317 -29932
rect 11553 -30168 11657 -29932
rect 11893 -30168 11997 -29932
rect 12233 -30168 12317 -29932
rect 12553 -30168 12657 -29932
rect 12893 -30168 12997 -29932
rect 13233 -30168 13317 -29932
rect 13553 -30168 13657 -29932
rect 13893 -30168 13997 -29932
rect 14233 -30168 14317 -29932
rect 14553 -30168 14657 -29932
rect 14893 -30168 14997 -29932
rect 15233 -30168 15317 -29932
rect 15553 -30168 15657 -29932
rect 15893 -30168 15997 -29932
rect 16233 -30168 16317 -29932
rect 16553 -30168 16657 -29932
rect 16893 -30168 16997 -29932
rect 17233 -30168 17317 -29932
rect 17553 -30168 17657 -29932
rect 17893 -30168 17997 -29932
rect 18233 -30168 18317 -29932
rect 18553 -30168 18657 -29932
rect 18893 -30168 18997 -29932
rect 19233 -30168 19317 -29932
rect 19553 -30168 19657 -29932
rect 19893 -30168 19997 -29932
rect 20233 -30168 20317 -29932
rect 20553 -30168 20657 -29932
rect 20893 -30168 20997 -29932
rect 21233 -30168 21317 -29932
rect 21553 -30168 21657 -29932
rect 21893 -30168 21997 -29932
rect 22233 -30168 22317 -29932
rect 22553 -30168 22657 -29932
rect 22893 -30168 22997 -29932
rect 23233 -30168 23317 -29932
rect 23553 -30168 23657 -29932
rect 23893 -30168 23997 -29932
rect 24233 -30168 24317 -29932
rect 24553 -30168 24657 -29932
rect 24893 -30168 24997 -29932
rect 25233 -30168 25317 -29932
rect 25553 -30168 25657 -29932
rect 25893 -30168 25997 -29932
rect 26233 -30168 26317 -29932
rect 26553 -30168 26657 -29932
rect 26893 -30168 26997 -29932
rect 27233 -30168 27317 -29932
rect 27553 -30168 27657 -29932
rect 27893 -30168 27997 -29932
rect 28233 -30168 28317 -29932
rect 28553 -30168 28657 -29932
rect 28893 -30168 28997 -29932
rect 29233 -30168 29317 -29932
rect 29553 -30168 29657 -29932
rect 29893 -30168 29997 -29932
rect 30233 -30168 30317 -29932
rect 30553 -30168 30657 -29932
rect 30893 -30168 30997 -29932
rect 31233 -30168 31317 -29932
rect 31553 -30168 31657 -29932
rect 31893 -30168 31997 -29932
rect 32233 -30168 32317 -29932
rect 32553 -30168 32657 -29932
rect 32893 -30168 32997 -29932
rect 33233 -30168 33317 -29932
rect 33553 -30168 33657 -29932
rect 33893 -30168 33997 -29932
rect 34233 -30168 34275 -29932
rect 8275 -30210 34275 -30168
rect 8615 -30272 8935 -30210
rect 8615 -30508 8657 -30272
rect 8893 -30508 8935 -30272
rect 8615 -30592 8935 -30508
rect 8615 -30828 8657 -30592
rect 8893 -30828 8935 -30592
rect 8615 -30890 8935 -30828
rect 9615 -30272 9935 -30210
rect 9615 -30508 9657 -30272
rect 9893 -30508 9935 -30272
rect 9615 -30592 9935 -30508
rect 9615 -30828 9657 -30592
rect 9893 -30828 9935 -30592
rect 9615 -30890 9935 -30828
rect 10615 -30272 10935 -30210
rect 10615 -30508 10657 -30272
rect 10893 -30508 10935 -30272
rect 10615 -30592 10935 -30508
rect 10615 -30828 10657 -30592
rect 10893 -30828 10935 -30592
rect 10615 -30890 10935 -30828
rect 11615 -30272 11935 -30210
rect 11615 -30508 11657 -30272
rect 11893 -30508 11935 -30272
rect 11615 -30592 11935 -30508
rect 11615 -30828 11657 -30592
rect 11893 -30828 11935 -30592
rect 11615 -30890 11935 -30828
rect 12615 -30272 12935 -30210
rect 12615 -30508 12657 -30272
rect 12893 -30508 12935 -30272
rect 12615 -30592 12935 -30508
rect 12615 -30828 12657 -30592
rect 12893 -30828 12935 -30592
rect 12615 -30890 12935 -30828
rect 13615 -30272 13935 -30210
rect 13615 -30508 13657 -30272
rect 13893 -30508 13935 -30272
rect 13615 -30592 13935 -30508
rect 13615 -30828 13657 -30592
rect 13893 -30828 13935 -30592
rect 13615 -30890 13935 -30828
rect 14615 -30272 14935 -30210
rect 14615 -30508 14657 -30272
rect 14893 -30508 14935 -30272
rect 14615 -30592 14935 -30508
rect 14615 -30828 14657 -30592
rect 14893 -30828 14935 -30592
rect 14615 -30890 14935 -30828
rect 15615 -30272 15935 -30210
rect 15615 -30508 15657 -30272
rect 15893 -30508 15935 -30272
rect 15615 -30592 15935 -30508
rect 15615 -30828 15657 -30592
rect 15893 -30828 15935 -30592
rect 15615 -30890 15935 -30828
rect 16615 -30272 16935 -30210
rect 16615 -30508 16657 -30272
rect 16893 -30508 16935 -30272
rect 16615 -30592 16935 -30508
rect 16615 -30828 16657 -30592
rect 16893 -30828 16935 -30592
rect 16615 -30890 16935 -30828
rect 17615 -30272 17935 -30210
rect 17615 -30508 17657 -30272
rect 17893 -30508 17935 -30272
rect 17615 -30592 17935 -30508
rect 17615 -30828 17657 -30592
rect 17893 -30828 17935 -30592
rect 17615 -30890 17935 -30828
rect 18615 -30272 18935 -30210
rect 18615 -30508 18657 -30272
rect 18893 -30508 18935 -30272
rect 18615 -30592 18935 -30508
rect 18615 -30828 18657 -30592
rect 18893 -30828 18935 -30592
rect 18615 -30890 18935 -30828
rect 19615 -30272 19935 -30210
rect 19615 -30508 19657 -30272
rect 19893 -30508 19935 -30272
rect 19615 -30592 19935 -30508
rect 19615 -30828 19657 -30592
rect 19893 -30828 19935 -30592
rect 19615 -30890 19935 -30828
rect 20615 -30272 20935 -30210
rect 20615 -30508 20657 -30272
rect 20893 -30508 20935 -30272
rect 20615 -30592 20935 -30508
rect 20615 -30828 20657 -30592
rect 20893 -30828 20935 -30592
rect 20615 -30890 20935 -30828
rect 21615 -30272 21935 -30210
rect 21615 -30508 21657 -30272
rect 21893 -30508 21935 -30272
rect 21615 -30592 21935 -30508
rect 21615 -30828 21657 -30592
rect 21893 -30828 21935 -30592
rect 21615 -30890 21935 -30828
rect 22615 -30272 22935 -30210
rect 22615 -30508 22657 -30272
rect 22893 -30508 22935 -30272
rect 22615 -30592 22935 -30508
rect 22615 -30828 22657 -30592
rect 22893 -30828 22935 -30592
rect 22615 -30890 22935 -30828
rect 23615 -30272 23935 -30210
rect 23615 -30508 23657 -30272
rect 23893 -30508 23935 -30272
rect 23615 -30592 23935 -30508
rect 23615 -30828 23657 -30592
rect 23893 -30828 23935 -30592
rect 23615 -30890 23935 -30828
rect 24615 -30272 24935 -30210
rect 24615 -30508 24657 -30272
rect 24893 -30508 24935 -30272
rect 24615 -30592 24935 -30508
rect 24615 -30828 24657 -30592
rect 24893 -30828 24935 -30592
rect 24615 -30890 24935 -30828
rect 25615 -30272 25935 -30210
rect 25615 -30508 25657 -30272
rect 25893 -30508 25935 -30272
rect 25615 -30592 25935 -30508
rect 25615 -30828 25657 -30592
rect 25893 -30828 25935 -30592
rect 25615 -30890 25935 -30828
rect 26615 -30272 26935 -30210
rect 26615 -30508 26657 -30272
rect 26893 -30508 26935 -30272
rect 26615 -30592 26935 -30508
rect 26615 -30828 26657 -30592
rect 26893 -30828 26935 -30592
rect 26615 -30890 26935 -30828
rect 27615 -30272 27935 -30210
rect 27615 -30508 27657 -30272
rect 27893 -30508 27935 -30272
rect 27615 -30592 27935 -30508
rect 27615 -30828 27657 -30592
rect 27893 -30828 27935 -30592
rect 27615 -30890 27935 -30828
rect 28615 -30272 28935 -30210
rect 28615 -30508 28657 -30272
rect 28893 -30508 28935 -30272
rect 28615 -30592 28935 -30508
rect 28615 -30828 28657 -30592
rect 28893 -30828 28935 -30592
rect 28615 -30890 28935 -30828
rect 29615 -30272 29935 -30210
rect 29615 -30508 29657 -30272
rect 29893 -30508 29935 -30272
rect 29615 -30592 29935 -30508
rect 29615 -30828 29657 -30592
rect 29893 -30828 29935 -30592
rect 29615 -30890 29935 -30828
rect 30615 -30272 30935 -30210
rect 30615 -30508 30657 -30272
rect 30893 -30508 30935 -30272
rect 30615 -30592 30935 -30508
rect 30615 -30828 30657 -30592
rect 30893 -30828 30935 -30592
rect 30615 -30890 30935 -30828
rect 31615 -30272 31935 -30210
rect 31615 -30508 31657 -30272
rect 31893 -30508 31935 -30272
rect 31615 -30592 31935 -30508
rect 31615 -30828 31657 -30592
rect 31893 -30828 31935 -30592
rect 31615 -30890 31935 -30828
rect 32615 -30272 32935 -30210
rect 32615 -30508 32657 -30272
rect 32893 -30508 32935 -30272
rect 32615 -30592 32935 -30508
rect 32615 -30828 32657 -30592
rect 32893 -30828 32935 -30592
rect 32615 -30890 32935 -30828
rect 33615 -30272 33935 -30210
rect 33615 -30508 33657 -30272
rect 33893 -30508 33935 -30272
rect 33615 -30592 33935 -30508
rect 33615 -30828 33657 -30592
rect 33893 -30828 33935 -30592
rect 33615 -30890 33935 -30828
rect 8275 -30932 34275 -30890
rect 8275 -31168 8317 -30932
rect 8553 -31168 8657 -30932
rect 8893 -31168 8997 -30932
rect 9233 -31168 9317 -30932
rect 9553 -31168 9657 -30932
rect 9893 -31168 9997 -30932
rect 10233 -31168 10317 -30932
rect 10553 -31168 10657 -30932
rect 10893 -31168 10997 -30932
rect 11233 -31168 11317 -30932
rect 11553 -31168 11657 -30932
rect 11893 -31168 11997 -30932
rect 12233 -31168 12317 -30932
rect 12553 -31168 12657 -30932
rect 12893 -31168 12997 -30932
rect 13233 -31168 13317 -30932
rect 13553 -31168 13657 -30932
rect 13893 -31168 13997 -30932
rect 14233 -31168 14317 -30932
rect 14553 -31168 14657 -30932
rect 14893 -31168 14997 -30932
rect 15233 -31168 15317 -30932
rect 15553 -31168 15657 -30932
rect 15893 -31168 15997 -30932
rect 16233 -31168 16317 -30932
rect 16553 -31168 16657 -30932
rect 16893 -31168 16997 -30932
rect 17233 -31168 17317 -30932
rect 17553 -31168 17657 -30932
rect 17893 -31168 17997 -30932
rect 18233 -31168 18317 -30932
rect 18553 -31168 18657 -30932
rect 18893 -31168 18997 -30932
rect 19233 -31168 19317 -30932
rect 19553 -31168 19657 -30932
rect 19893 -31168 19997 -30932
rect 20233 -31168 20317 -30932
rect 20553 -31168 20657 -30932
rect 20893 -31168 20997 -30932
rect 21233 -31168 21317 -30932
rect 21553 -31168 21657 -30932
rect 21893 -31168 21997 -30932
rect 22233 -31168 22317 -30932
rect 22553 -31168 22657 -30932
rect 22893 -31168 22997 -30932
rect 23233 -31168 23317 -30932
rect 23553 -31168 23657 -30932
rect 23893 -31168 23997 -30932
rect 24233 -31168 24317 -30932
rect 24553 -31168 24657 -30932
rect 24893 -31168 24997 -30932
rect 25233 -31168 25317 -30932
rect 25553 -31168 25657 -30932
rect 25893 -31168 25997 -30932
rect 26233 -31168 26317 -30932
rect 26553 -31168 26657 -30932
rect 26893 -31168 26997 -30932
rect 27233 -31168 27317 -30932
rect 27553 -31168 27657 -30932
rect 27893 -31168 27997 -30932
rect 28233 -31168 28317 -30932
rect 28553 -31168 28657 -30932
rect 28893 -31168 28997 -30932
rect 29233 -31168 29317 -30932
rect 29553 -31168 29657 -30932
rect 29893 -31168 29997 -30932
rect 30233 -31168 30317 -30932
rect 30553 -31168 30657 -30932
rect 30893 -31168 30997 -30932
rect 31233 -31168 31317 -30932
rect 31553 -31168 31657 -30932
rect 31893 -31168 31997 -30932
rect 32233 -31168 32317 -30932
rect 32553 -31168 32657 -30932
rect 32893 -31168 32997 -30932
rect 33233 -31168 33317 -30932
rect 33553 -31168 33657 -30932
rect 33893 -31168 33997 -30932
rect 34233 -31168 34275 -30932
rect 8275 -31210 34275 -31168
rect 8615 -31272 8935 -31210
rect 8615 -31508 8657 -31272
rect 8893 -31508 8935 -31272
rect 8615 -31592 8935 -31508
rect 8615 -31828 8657 -31592
rect 8893 -31828 8935 -31592
rect 8615 -31890 8935 -31828
rect 9615 -31272 9935 -31210
rect 9615 -31508 9657 -31272
rect 9893 -31508 9935 -31272
rect 9615 -31592 9935 -31508
rect 9615 -31828 9657 -31592
rect 9893 -31828 9935 -31592
rect 9615 -31890 9935 -31828
rect 10615 -31272 10935 -31210
rect 10615 -31508 10657 -31272
rect 10893 -31508 10935 -31272
rect 10615 -31592 10935 -31508
rect 10615 -31828 10657 -31592
rect 10893 -31828 10935 -31592
rect 10615 -31890 10935 -31828
rect 11615 -31272 11935 -31210
rect 11615 -31508 11657 -31272
rect 11893 -31508 11935 -31272
rect 11615 -31592 11935 -31508
rect 11615 -31828 11657 -31592
rect 11893 -31828 11935 -31592
rect 11615 -31890 11935 -31828
rect 12615 -31272 12935 -31210
rect 12615 -31508 12657 -31272
rect 12893 -31508 12935 -31272
rect 12615 -31592 12935 -31508
rect 12615 -31828 12657 -31592
rect 12893 -31828 12935 -31592
rect 12615 -31890 12935 -31828
rect 13615 -31272 13935 -31210
rect 13615 -31508 13657 -31272
rect 13893 -31508 13935 -31272
rect 13615 -31592 13935 -31508
rect 13615 -31828 13657 -31592
rect 13893 -31828 13935 -31592
rect 13615 -31890 13935 -31828
rect 14615 -31272 14935 -31210
rect 14615 -31508 14657 -31272
rect 14893 -31508 14935 -31272
rect 14615 -31592 14935 -31508
rect 14615 -31828 14657 -31592
rect 14893 -31828 14935 -31592
rect 14615 -31890 14935 -31828
rect 15615 -31272 15935 -31210
rect 15615 -31508 15657 -31272
rect 15893 -31508 15935 -31272
rect 15615 -31592 15935 -31508
rect 15615 -31828 15657 -31592
rect 15893 -31828 15935 -31592
rect 15615 -31890 15935 -31828
rect 16615 -31272 16935 -31210
rect 16615 -31508 16657 -31272
rect 16893 -31508 16935 -31272
rect 16615 -31592 16935 -31508
rect 16615 -31828 16657 -31592
rect 16893 -31828 16935 -31592
rect 16615 -31890 16935 -31828
rect 17615 -31272 17935 -31210
rect 17615 -31508 17657 -31272
rect 17893 -31508 17935 -31272
rect 17615 -31592 17935 -31508
rect 17615 -31828 17657 -31592
rect 17893 -31828 17935 -31592
rect 17615 -31890 17935 -31828
rect 18615 -31272 18935 -31210
rect 18615 -31508 18657 -31272
rect 18893 -31508 18935 -31272
rect 18615 -31592 18935 -31508
rect 18615 -31828 18657 -31592
rect 18893 -31828 18935 -31592
rect 18615 -31890 18935 -31828
rect 19615 -31272 19935 -31210
rect 19615 -31508 19657 -31272
rect 19893 -31508 19935 -31272
rect 19615 -31592 19935 -31508
rect 19615 -31828 19657 -31592
rect 19893 -31828 19935 -31592
rect 19615 -31890 19935 -31828
rect 20615 -31272 20935 -31210
rect 20615 -31508 20657 -31272
rect 20893 -31508 20935 -31272
rect 20615 -31592 20935 -31508
rect 20615 -31828 20657 -31592
rect 20893 -31828 20935 -31592
rect 20615 -31890 20935 -31828
rect 21615 -31272 21935 -31210
rect 21615 -31508 21657 -31272
rect 21893 -31508 21935 -31272
rect 21615 -31592 21935 -31508
rect 21615 -31828 21657 -31592
rect 21893 -31828 21935 -31592
rect 21615 -31890 21935 -31828
rect 22615 -31272 22935 -31210
rect 22615 -31508 22657 -31272
rect 22893 -31508 22935 -31272
rect 22615 -31592 22935 -31508
rect 22615 -31828 22657 -31592
rect 22893 -31828 22935 -31592
rect 22615 -31890 22935 -31828
rect 23615 -31272 23935 -31210
rect 23615 -31508 23657 -31272
rect 23893 -31508 23935 -31272
rect 23615 -31592 23935 -31508
rect 23615 -31828 23657 -31592
rect 23893 -31828 23935 -31592
rect 23615 -31890 23935 -31828
rect 24615 -31272 24935 -31210
rect 24615 -31508 24657 -31272
rect 24893 -31508 24935 -31272
rect 24615 -31592 24935 -31508
rect 24615 -31828 24657 -31592
rect 24893 -31828 24935 -31592
rect 24615 -31890 24935 -31828
rect 25615 -31272 25935 -31210
rect 25615 -31508 25657 -31272
rect 25893 -31508 25935 -31272
rect 25615 -31592 25935 -31508
rect 25615 -31828 25657 -31592
rect 25893 -31828 25935 -31592
rect 25615 -31890 25935 -31828
rect 26615 -31272 26935 -31210
rect 26615 -31508 26657 -31272
rect 26893 -31508 26935 -31272
rect 26615 -31592 26935 -31508
rect 26615 -31828 26657 -31592
rect 26893 -31828 26935 -31592
rect 26615 -31890 26935 -31828
rect 27615 -31272 27935 -31210
rect 27615 -31508 27657 -31272
rect 27893 -31508 27935 -31272
rect 27615 -31592 27935 -31508
rect 27615 -31828 27657 -31592
rect 27893 -31828 27935 -31592
rect 27615 -31890 27935 -31828
rect 28615 -31272 28935 -31210
rect 28615 -31508 28657 -31272
rect 28893 -31508 28935 -31272
rect 28615 -31592 28935 -31508
rect 28615 -31828 28657 -31592
rect 28893 -31828 28935 -31592
rect 28615 -31890 28935 -31828
rect 29615 -31272 29935 -31210
rect 29615 -31508 29657 -31272
rect 29893 -31508 29935 -31272
rect 29615 -31592 29935 -31508
rect 29615 -31828 29657 -31592
rect 29893 -31828 29935 -31592
rect 29615 -31890 29935 -31828
rect 30615 -31272 30935 -31210
rect 30615 -31508 30657 -31272
rect 30893 -31508 30935 -31272
rect 30615 -31592 30935 -31508
rect 30615 -31828 30657 -31592
rect 30893 -31828 30935 -31592
rect 30615 -31890 30935 -31828
rect 31615 -31272 31935 -31210
rect 31615 -31508 31657 -31272
rect 31893 -31508 31935 -31272
rect 31615 -31592 31935 -31508
rect 31615 -31828 31657 -31592
rect 31893 -31828 31935 -31592
rect 31615 -31890 31935 -31828
rect 32615 -31272 32935 -31210
rect 32615 -31508 32657 -31272
rect 32893 -31508 32935 -31272
rect 32615 -31592 32935 -31508
rect 32615 -31828 32657 -31592
rect 32893 -31828 32935 -31592
rect 32615 -31890 32935 -31828
rect 33615 -31272 33935 -31210
rect 33615 -31508 33657 -31272
rect 33893 -31508 33935 -31272
rect 33615 -31592 33935 -31508
rect 33615 -31828 33657 -31592
rect 33893 -31828 33935 -31592
rect 33615 -31890 33935 -31828
rect 8275 -31932 34275 -31890
rect 8275 -32168 8317 -31932
rect 8553 -32168 8657 -31932
rect 8893 -32168 8997 -31932
rect 9233 -32168 9317 -31932
rect 9553 -32168 9657 -31932
rect 9893 -32168 9997 -31932
rect 10233 -32168 10317 -31932
rect 10553 -32168 10657 -31932
rect 10893 -32168 10997 -31932
rect 11233 -32168 11317 -31932
rect 11553 -32168 11657 -31932
rect 11893 -32168 11997 -31932
rect 12233 -32168 12317 -31932
rect 12553 -32168 12657 -31932
rect 12893 -32168 12997 -31932
rect 13233 -32168 13317 -31932
rect 13553 -32168 13657 -31932
rect 13893 -32168 13997 -31932
rect 14233 -32168 14317 -31932
rect 14553 -32168 14657 -31932
rect 14893 -32168 14997 -31932
rect 15233 -32168 15317 -31932
rect 15553 -32168 15657 -31932
rect 15893 -32168 15997 -31932
rect 16233 -32168 16317 -31932
rect 16553 -32168 16657 -31932
rect 16893 -32168 16997 -31932
rect 17233 -32168 17317 -31932
rect 17553 -32168 17657 -31932
rect 17893 -32168 17997 -31932
rect 18233 -32168 18317 -31932
rect 18553 -32168 18657 -31932
rect 18893 -32168 18997 -31932
rect 19233 -32168 19317 -31932
rect 19553 -32168 19657 -31932
rect 19893 -32168 19997 -31932
rect 20233 -32168 20317 -31932
rect 20553 -32168 20657 -31932
rect 20893 -32168 20997 -31932
rect 21233 -32168 21317 -31932
rect 21553 -32168 21657 -31932
rect 21893 -32168 21997 -31932
rect 22233 -32168 22317 -31932
rect 22553 -32168 22657 -31932
rect 22893 -32168 22997 -31932
rect 23233 -32168 23317 -31932
rect 23553 -32168 23657 -31932
rect 23893 -32168 23997 -31932
rect 24233 -32168 24317 -31932
rect 24553 -32168 24657 -31932
rect 24893 -32168 24997 -31932
rect 25233 -32168 25317 -31932
rect 25553 -32168 25657 -31932
rect 25893 -32168 25997 -31932
rect 26233 -32168 26317 -31932
rect 26553 -32168 26657 -31932
rect 26893 -32168 26997 -31932
rect 27233 -32168 27317 -31932
rect 27553 -32168 27657 -31932
rect 27893 -32168 27997 -31932
rect 28233 -32168 28317 -31932
rect 28553 -32168 28657 -31932
rect 28893 -32168 28997 -31932
rect 29233 -32168 29317 -31932
rect 29553 -32168 29657 -31932
rect 29893 -32168 29997 -31932
rect 30233 -32168 30317 -31932
rect 30553 -32168 30657 -31932
rect 30893 -32168 30997 -31932
rect 31233 -32168 31317 -31932
rect 31553 -32168 31657 -31932
rect 31893 -32168 31997 -31932
rect 32233 -32168 32317 -31932
rect 32553 -32168 32657 -31932
rect 32893 -32168 32997 -31932
rect 33233 -32168 33317 -31932
rect 33553 -32168 33657 -31932
rect 33893 -32168 33997 -31932
rect 34233 -32168 34275 -31932
rect 8275 -32210 34275 -32168
rect 8615 -32272 8935 -32210
rect 8615 -32508 8657 -32272
rect 8893 -32508 8935 -32272
rect -49485 -32828 -49443 -32592
rect -49207 -32828 -49165 -32592
rect -49485 -32890 -49165 -32828
rect -46275 -32580 -36155 -32550
tri -36155 -32580 -36125 -32550 nw
tri -22905 -32580 -22875 -32550 se
rect -22875 -32580 -17675 -32550
tri -17675 -32580 -17645 -32550 sw
tri -4425 -32580 -4395 -32550 ne
rect -4395 -32580 5725 -32550
rect -46275 -32672 -36275 -32580
rect -74825 -32932 -48825 -32890
rect -74825 -33168 -74783 -32932
rect -74547 -33168 -74443 -32932
rect -74207 -33168 -74103 -32932
rect -73867 -33168 -73783 -32932
rect -73547 -33168 -73443 -32932
rect -73207 -33168 -73103 -32932
rect -72867 -33168 -72783 -32932
rect -72547 -33168 -72443 -32932
rect -72207 -33168 -72103 -32932
rect -71867 -33168 -71783 -32932
rect -71547 -33168 -71443 -32932
rect -71207 -33168 -71103 -32932
rect -70867 -33168 -70783 -32932
rect -70547 -33168 -70443 -32932
rect -70207 -33168 -70103 -32932
rect -69867 -33168 -69783 -32932
rect -69547 -33168 -69443 -32932
rect -69207 -33168 -69103 -32932
rect -68867 -33168 -68783 -32932
rect -68547 -33168 -68443 -32932
rect -68207 -33168 -68103 -32932
rect -67867 -33168 -67783 -32932
rect -67547 -33168 -67443 -32932
rect -67207 -33168 -67103 -32932
rect -66867 -33168 -66783 -32932
rect -66547 -33168 -66443 -32932
rect -66207 -33168 -66103 -32932
rect -65867 -33168 -65783 -32932
rect -65547 -33168 -65443 -32932
rect -65207 -33168 -65103 -32932
rect -64867 -33168 -64783 -32932
rect -64547 -33168 -64443 -32932
rect -64207 -33168 -64103 -32932
rect -63867 -33168 -63783 -32932
rect -63547 -33168 -63443 -32932
rect -63207 -33168 -63103 -32932
rect -62867 -33168 -62783 -32932
rect -62547 -33168 -62443 -32932
rect -62207 -33168 -62103 -32932
rect -61867 -33168 -61783 -32932
rect -61547 -33168 -61443 -32932
rect -61207 -33168 -61103 -32932
rect -60867 -33168 -60783 -32932
rect -60547 -33168 -60443 -32932
rect -60207 -33168 -60103 -32932
rect -59867 -33168 -59783 -32932
rect -59547 -33168 -59443 -32932
rect -59207 -33168 -59103 -32932
rect -58867 -33168 -58783 -32932
rect -58547 -33168 -58443 -32932
rect -58207 -33168 -58103 -32932
rect -57867 -33168 -57783 -32932
rect -57547 -33168 -57443 -32932
rect -57207 -33168 -57103 -32932
rect -56867 -33168 -56783 -32932
rect -56547 -33168 -56443 -32932
rect -56207 -33168 -56103 -32932
rect -55867 -33168 -55783 -32932
rect -55547 -33168 -55443 -32932
rect -55207 -33168 -55103 -32932
rect -54867 -33168 -54783 -32932
rect -54547 -33168 -54443 -32932
rect -54207 -33168 -54103 -32932
rect -53867 -33168 -53783 -32932
rect -53547 -33168 -53443 -32932
rect -53207 -33168 -53103 -32932
rect -52867 -33168 -52783 -32932
rect -52547 -33168 -52443 -32932
rect -52207 -33168 -52103 -32932
rect -51867 -33168 -51783 -32932
rect -51547 -33168 -51443 -32932
rect -51207 -33168 -51103 -32932
rect -50867 -33168 -50783 -32932
rect -50547 -33168 -50443 -32932
rect -50207 -33168 -50103 -32932
rect -49867 -33168 -49783 -32932
rect -49547 -33168 -49443 -32932
rect -49207 -33168 -49103 -32932
rect -48867 -33168 -48825 -32932
rect -74825 -33210 -48825 -33168
rect -74485 -33272 -74165 -33210
rect -74485 -33508 -74443 -33272
rect -74207 -33508 -74165 -33272
rect -74485 -33592 -74165 -33508
rect -74485 -33828 -74443 -33592
rect -74207 -33828 -74165 -33592
rect -74485 -33890 -74165 -33828
rect -73485 -33272 -73165 -33210
rect -73485 -33508 -73443 -33272
rect -73207 -33508 -73165 -33272
rect -73485 -33592 -73165 -33508
rect -73485 -33828 -73443 -33592
rect -73207 -33828 -73165 -33592
rect -73485 -33890 -73165 -33828
rect -72485 -33272 -72165 -33210
rect -72485 -33508 -72443 -33272
rect -72207 -33508 -72165 -33272
rect -72485 -33592 -72165 -33508
rect -72485 -33828 -72443 -33592
rect -72207 -33828 -72165 -33592
rect -72485 -33890 -72165 -33828
rect -71485 -33272 -71165 -33210
rect -71485 -33508 -71443 -33272
rect -71207 -33508 -71165 -33272
rect -71485 -33592 -71165 -33508
rect -71485 -33828 -71443 -33592
rect -71207 -33828 -71165 -33592
rect -71485 -33890 -71165 -33828
rect -70485 -33272 -70165 -33210
rect -70485 -33508 -70443 -33272
rect -70207 -33508 -70165 -33272
rect -70485 -33592 -70165 -33508
rect -70485 -33828 -70443 -33592
rect -70207 -33828 -70165 -33592
rect -70485 -33890 -70165 -33828
rect -69485 -33272 -69165 -33210
rect -69485 -33508 -69443 -33272
rect -69207 -33508 -69165 -33272
rect -69485 -33592 -69165 -33508
rect -69485 -33828 -69443 -33592
rect -69207 -33828 -69165 -33592
rect -69485 -33890 -69165 -33828
rect -68485 -33272 -68165 -33210
rect -68485 -33508 -68443 -33272
rect -68207 -33508 -68165 -33272
rect -68485 -33592 -68165 -33508
rect -68485 -33828 -68443 -33592
rect -68207 -33828 -68165 -33592
rect -68485 -33890 -68165 -33828
rect -67485 -33272 -67165 -33210
rect -67485 -33508 -67443 -33272
rect -67207 -33508 -67165 -33272
rect -67485 -33592 -67165 -33508
rect -67485 -33828 -67443 -33592
rect -67207 -33828 -67165 -33592
rect -67485 -33890 -67165 -33828
rect -66485 -33272 -66165 -33210
rect -66485 -33508 -66443 -33272
rect -66207 -33508 -66165 -33272
rect -66485 -33592 -66165 -33508
rect -66485 -33828 -66443 -33592
rect -66207 -33828 -66165 -33592
rect -66485 -33890 -66165 -33828
rect -65485 -33272 -65165 -33210
rect -65485 -33508 -65443 -33272
rect -65207 -33508 -65165 -33272
rect -65485 -33592 -65165 -33508
rect -65485 -33828 -65443 -33592
rect -65207 -33828 -65165 -33592
rect -65485 -33890 -65165 -33828
rect -64485 -33272 -64165 -33210
rect -64485 -33508 -64443 -33272
rect -64207 -33508 -64165 -33272
rect -64485 -33592 -64165 -33508
rect -64485 -33828 -64443 -33592
rect -64207 -33828 -64165 -33592
rect -64485 -33890 -64165 -33828
rect -63485 -33272 -63165 -33210
rect -63485 -33508 -63443 -33272
rect -63207 -33508 -63165 -33272
rect -63485 -33592 -63165 -33508
rect -63485 -33828 -63443 -33592
rect -63207 -33828 -63165 -33592
rect -63485 -33890 -63165 -33828
rect -62485 -33272 -62165 -33210
rect -62485 -33508 -62443 -33272
rect -62207 -33508 -62165 -33272
rect -62485 -33592 -62165 -33508
rect -62485 -33828 -62443 -33592
rect -62207 -33828 -62165 -33592
rect -62485 -33890 -62165 -33828
rect -61485 -33272 -61165 -33210
rect -61485 -33508 -61443 -33272
rect -61207 -33508 -61165 -33272
rect -61485 -33592 -61165 -33508
rect -61485 -33828 -61443 -33592
rect -61207 -33828 -61165 -33592
rect -61485 -33890 -61165 -33828
rect -60485 -33272 -60165 -33210
rect -60485 -33508 -60443 -33272
rect -60207 -33508 -60165 -33272
rect -60485 -33592 -60165 -33508
rect -60485 -33828 -60443 -33592
rect -60207 -33828 -60165 -33592
rect -60485 -33890 -60165 -33828
rect -59485 -33272 -59165 -33210
rect -59485 -33508 -59443 -33272
rect -59207 -33508 -59165 -33272
rect -59485 -33592 -59165 -33508
rect -59485 -33828 -59443 -33592
rect -59207 -33828 -59165 -33592
rect -59485 -33890 -59165 -33828
rect -58485 -33272 -58165 -33210
rect -58485 -33508 -58443 -33272
rect -58207 -33508 -58165 -33272
rect -58485 -33592 -58165 -33508
rect -58485 -33828 -58443 -33592
rect -58207 -33828 -58165 -33592
rect -58485 -33890 -58165 -33828
rect -57485 -33272 -57165 -33210
rect -57485 -33508 -57443 -33272
rect -57207 -33508 -57165 -33272
rect -57485 -33592 -57165 -33508
rect -57485 -33828 -57443 -33592
rect -57207 -33828 -57165 -33592
rect -57485 -33890 -57165 -33828
rect -56485 -33272 -56165 -33210
rect -56485 -33508 -56443 -33272
rect -56207 -33508 -56165 -33272
rect -56485 -33592 -56165 -33508
rect -56485 -33828 -56443 -33592
rect -56207 -33828 -56165 -33592
rect -56485 -33890 -56165 -33828
rect -55485 -33272 -55165 -33210
rect -55485 -33508 -55443 -33272
rect -55207 -33508 -55165 -33272
rect -55485 -33592 -55165 -33508
rect -55485 -33828 -55443 -33592
rect -55207 -33828 -55165 -33592
rect -55485 -33890 -55165 -33828
rect -54485 -33272 -54165 -33210
rect -54485 -33508 -54443 -33272
rect -54207 -33508 -54165 -33272
rect -54485 -33592 -54165 -33508
rect -54485 -33828 -54443 -33592
rect -54207 -33828 -54165 -33592
rect -54485 -33890 -54165 -33828
rect -53485 -33272 -53165 -33210
rect -53485 -33508 -53443 -33272
rect -53207 -33508 -53165 -33272
rect -53485 -33592 -53165 -33508
rect -53485 -33828 -53443 -33592
rect -53207 -33828 -53165 -33592
rect -53485 -33890 -53165 -33828
rect -52485 -33272 -52165 -33210
rect -52485 -33508 -52443 -33272
rect -52207 -33508 -52165 -33272
rect -52485 -33592 -52165 -33508
rect -52485 -33828 -52443 -33592
rect -52207 -33828 -52165 -33592
rect -52485 -33890 -52165 -33828
rect -51485 -33272 -51165 -33210
rect -51485 -33508 -51443 -33272
rect -51207 -33508 -51165 -33272
rect -51485 -33592 -51165 -33508
rect -51485 -33828 -51443 -33592
rect -51207 -33828 -51165 -33592
rect -51485 -33890 -51165 -33828
rect -50485 -33272 -50165 -33210
rect -50485 -33508 -50443 -33272
rect -50207 -33508 -50165 -33272
rect -50485 -33592 -50165 -33508
rect -50485 -33828 -50443 -33592
rect -50207 -33828 -50165 -33592
rect -50485 -33890 -50165 -33828
rect -49485 -33272 -49165 -33210
rect -49485 -33508 -49443 -33272
rect -49207 -33508 -49165 -33272
rect -49485 -33592 -49165 -33508
rect -49485 -33828 -49443 -33592
rect -49207 -33828 -49165 -33592
rect -49485 -33890 -49165 -33828
rect -74825 -33932 -48825 -33890
rect -74825 -34168 -74783 -33932
rect -74547 -34168 -74443 -33932
rect -74207 -34168 -74103 -33932
rect -73867 -34168 -73783 -33932
rect -73547 -34168 -73443 -33932
rect -73207 -34168 -73103 -33932
rect -72867 -34168 -72783 -33932
rect -72547 -34168 -72443 -33932
rect -72207 -34168 -72103 -33932
rect -71867 -34168 -71783 -33932
rect -71547 -34168 -71443 -33932
rect -71207 -34168 -71103 -33932
rect -70867 -34168 -70783 -33932
rect -70547 -34168 -70443 -33932
rect -70207 -34168 -70103 -33932
rect -69867 -34168 -69783 -33932
rect -69547 -34168 -69443 -33932
rect -69207 -34168 -69103 -33932
rect -68867 -34168 -68783 -33932
rect -68547 -34168 -68443 -33932
rect -68207 -34168 -68103 -33932
rect -67867 -34168 -67783 -33932
rect -67547 -34168 -67443 -33932
rect -67207 -34168 -67103 -33932
rect -66867 -34168 -66783 -33932
rect -66547 -34168 -66443 -33932
rect -66207 -34168 -66103 -33932
rect -65867 -34168 -65783 -33932
rect -65547 -34168 -65443 -33932
rect -65207 -34168 -65103 -33932
rect -64867 -34168 -64783 -33932
rect -64547 -34168 -64443 -33932
rect -64207 -34168 -64103 -33932
rect -63867 -34168 -63783 -33932
rect -63547 -34168 -63443 -33932
rect -63207 -34168 -63103 -33932
rect -62867 -34168 -62783 -33932
rect -62547 -34168 -62443 -33932
rect -62207 -34168 -62103 -33932
rect -61867 -34168 -61783 -33932
rect -61547 -34168 -61443 -33932
rect -61207 -34168 -61103 -33932
rect -60867 -34168 -60783 -33932
rect -60547 -34168 -60443 -33932
rect -60207 -34168 -60103 -33932
rect -59867 -34168 -59783 -33932
rect -59547 -34168 -59443 -33932
rect -59207 -34168 -59103 -33932
rect -58867 -34168 -58783 -33932
rect -58547 -34168 -58443 -33932
rect -58207 -34168 -58103 -33932
rect -57867 -34168 -57783 -33932
rect -57547 -34168 -57443 -33932
rect -57207 -34168 -57103 -33932
rect -56867 -34168 -56783 -33932
rect -56547 -34168 -56443 -33932
rect -56207 -34168 -56103 -33932
rect -55867 -34168 -55783 -33932
rect -55547 -34168 -55443 -33932
rect -55207 -34168 -55103 -33932
rect -54867 -34168 -54783 -33932
rect -54547 -34168 -54443 -33932
rect -54207 -34168 -54103 -33932
rect -53867 -34168 -53783 -33932
rect -53547 -34168 -53443 -33932
rect -53207 -34168 -53103 -33932
rect -52867 -34168 -52783 -33932
rect -52547 -34168 -52443 -33932
rect -52207 -34168 -52103 -33932
rect -51867 -34168 -51783 -33932
rect -51547 -34168 -51443 -33932
rect -51207 -34168 -51103 -33932
rect -50867 -34168 -50783 -33932
rect -50547 -34168 -50443 -33932
rect -50207 -34168 -50103 -33932
rect -49867 -34168 -49783 -33932
rect -49547 -34168 -49443 -33932
rect -49207 -34168 -49103 -33932
rect -48867 -34168 -48825 -33932
rect -74825 -34210 -48825 -34168
rect -74485 -34272 -74165 -34210
rect -74485 -34508 -74443 -34272
rect -74207 -34508 -74165 -34272
rect -74485 -34592 -74165 -34508
rect -74485 -34828 -74443 -34592
rect -74207 -34828 -74165 -34592
rect -74485 -34890 -74165 -34828
rect -73485 -34272 -73165 -34210
rect -73485 -34508 -73443 -34272
rect -73207 -34508 -73165 -34272
rect -73485 -34592 -73165 -34508
rect -73485 -34828 -73443 -34592
rect -73207 -34828 -73165 -34592
rect -73485 -34890 -73165 -34828
rect -72485 -34272 -72165 -34210
rect -72485 -34508 -72443 -34272
rect -72207 -34508 -72165 -34272
rect -72485 -34592 -72165 -34508
rect -72485 -34828 -72443 -34592
rect -72207 -34828 -72165 -34592
rect -72485 -34890 -72165 -34828
rect -71485 -34272 -71165 -34210
rect -71485 -34508 -71443 -34272
rect -71207 -34508 -71165 -34272
rect -71485 -34592 -71165 -34508
rect -71485 -34828 -71443 -34592
rect -71207 -34828 -71165 -34592
rect -71485 -34890 -71165 -34828
rect -70485 -34272 -70165 -34210
rect -70485 -34508 -70443 -34272
rect -70207 -34508 -70165 -34272
rect -70485 -34592 -70165 -34508
rect -70485 -34828 -70443 -34592
rect -70207 -34828 -70165 -34592
rect -70485 -34890 -70165 -34828
rect -69485 -34272 -69165 -34210
rect -69485 -34508 -69443 -34272
rect -69207 -34508 -69165 -34272
rect -69485 -34592 -69165 -34508
rect -69485 -34828 -69443 -34592
rect -69207 -34828 -69165 -34592
rect -69485 -34890 -69165 -34828
rect -68485 -34272 -68165 -34210
rect -68485 -34508 -68443 -34272
rect -68207 -34508 -68165 -34272
rect -68485 -34592 -68165 -34508
rect -68485 -34828 -68443 -34592
rect -68207 -34828 -68165 -34592
rect -68485 -34890 -68165 -34828
rect -67485 -34272 -67165 -34210
rect -67485 -34508 -67443 -34272
rect -67207 -34508 -67165 -34272
rect -67485 -34592 -67165 -34508
rect -67485 -34828 -67443 -34592
rect -67207 -34828 -67165 -34592
rect -67485 -34890 -67165 -34828
rect -66485 -34272 -66165 -34210
rect -66485 -34508 -66443 -34272
rect -66207 -34508 -66165 -34272
rect -66485 -34592 -66165 -34508
rect -66485 -34828 -66443 -34592
rect -66207 -34828 -66165 -34592
rect -66485 -34890 -66165 -34828
rect -65485 -34272 -65165 -34210
rect -65485 -34508 -65443 -34272
rect -65207 -34508 -65165 -34272
rect -65485 -34592 -65165 -34508
rect -65485 -34828 -65443 -34592
rect -65207 -34828 -65165 -34592
rect -65485 -34890 -65165 -34828
rect -64485 -34272 -64165 -34210
rect -64485 -34508 -64443 -34272
rect -64207 -34508 -64165 -34272
rect -64485 -34592 -64165 -34508
rect -64485 -34828 -64443 -34592
rect -64207 -34828 -64165 -34592
rect -64485 -34890 -64165 -34828
rect -63485 -34272 -63165 -34210
rect -63485 -34508 -63443 -34272
rect -63207 -34508 -63165 -34272
rect -63485 -34592 -63165 -34508
rect -63485 -34828 -63443 -34592
rect -63207 -34828 -63165 -34592
rect -63485 -34890 -63165 -34828
rect -62485 -34272 -62165 -34210
rect -62485 -34508 -62443 -34272
rect -62207 -34508 -62165 -34272
rect -62485 -34592 -62165 -34508
rect -62485 -34828 -62443 -34592
rect -62207 -34828 -62165 -34592
rect -62485 -34890 -62165 -34828
rect -61485 -34272 -61165 -34210
rect -61485 -34508 -61443 -34272
rect -61207 -34508 -61165 -34272
rect -61485 -34592 -61165 -34508
rect -61485 -34828 -61443 -34592
rect -61207 -34828 -61165 -34592
rect -61485 -34890 -61165 -34828
rect -60485 -34272 -60165 -34210
rect -60485 -34508 -60443 -34272
rect -60207 -34508 -60165 -34272
rect -60485 -34592 -60165 -34508
rect -60485 -34828 -60443 -34592
rect -60207 -34828 -60165 -34592
rect -60485 -34890 -60165 -34828
rect -59485 -34272 -59165 -34210
rect -59485 -34508 -59443 -34272
rect -59207 -34508 -59165 -34272
rect -59485 -34592 -59165 -34508
rect -59485 -34828 -59443 -34592
rect -59207 -34828 -59165 -34592
rect -59485 -34890 -59165 -34828
rect -58485 -34272 -58165 -34210
rect -58485 -34508 -58443 -34272
rect -58207 -34508 -58165 -34272
rect -58485 -34592 -58165 -34508
rect -58485 -34828 -58443 -34592
rect -58207 -34828 -58165 -34592
rect -58485 -34890 -58165 -34828
rect -57485 -34272 -57165 -34210
rect -57485 -34508 -57443 -34272
rect -57207 -34508 -57165 -34272
rect -57485 -34592 -57165 -34508
rect -57485 -34828 -57443 -34592
rect -57207 -34828 -57165 -34592
rect -57485 -34890 -57165 -34828
rect -56485 -34272 -56165 -34210
rect -56485 -34508 -56443 -34272
rect -56207 -34508 -56165 -34272
rect -56485 -34592 -56165 -34508
rect -56485 -34828 -56443 -34592
rect -56207 -34828 -56165 -34592
rect -56485 -34890 -56165 -34828
rect -55485 -34272 -55165 -34210
rect -55485 -34508 -55443 -34272
rect -55207 -34508 -55165 -34272
rect -55485 -34592 -55165 -34508
rect -55485 -34828 -55443 -34592
rect -55207 -34828 -55165 -34592
rect -55485 -34890 -55165 -34828
rect -54485 -34272 -54165 -34210
rect -54485 -34508 -54443 -34272
rect -54207 -34508 -54165 -34272
rect -54485 -34592 -54165 -34508
rect -54485 -34828 -54443 -34592
rect -54207 -34828 -54165 -34592
rect -54485 -34890 -54165 -34828
rect -53485 -34272 -53165 -34210
rect -53485 -34508 -53443 -34272
rect -53207 -34508 -53165 -34272
rect -53485 -34592 -53165 -34508
rect -53485 -34828 -53443 -34592
rect -53207 -34828 -53165 -34592
rect -53485 -34890 -53165 -34828
rect -52485 -34272 -52165 -34210
rect -52485 -34508 -52443 -34272
rect -52207 -34508 -52165 -34272
rect -52485 -34592 -52165 -34508
rect -52485 -34828 -52443 -34592
rect -52207 -34828 -52165 -34592
rect -52485 -34890 -52165 -34828
rect -51485 -34272 -51165 -34210
rect -51485 -34508 -51443 -34272
rect -51207 -34508 -51165 -34272
rect -51485 -34592 -51165 -34508
rect -51485 -34828 -51443 -34592
rect -51207 -34828 -51165 -34592
rect -51485 -34890 -51165 -34828
rect -50485 -34272 -50165 -34210
rect -50485 -34508 -50443 -34272
rect -50207 -34508 -50165 -34272
rect -50485 -34592 -50165 -34508
rect -50485 -34828 -50443 -34592
rect -50207 -34828 -50165 -34592
rect -50485 -34890 -50165 -34828
rect -49485 -34272 -49165 -34210
rect -49485 -34508 -49443 -34272
rect -49207 -34508 -49165 -34272
rect -49485 -34592 -49165 -34508
rect -49485 -34828 -49443 -34592
rect -49207 -34828 -49165 -34592
rect -49485 -34890 -49165 -34828
rect -74825 -34932 -48825 -34890
rect -74825 -35168 -74783 -34932
rect -74547 -35168 -74443 -34932
rect -74207 -35168 -74103 -34932
rect -73867 -35168 -73783 -34932
rect -73547 -35168 -73443 -34932
rect -73207 -35168 -73103 -34932
rect -72867 -35168 -72783 -34932
rect -72547 -35168 -72443 -34932
rect -72207 -35168 -72103 -34932
rect -71867 -35168 -71783 -34932
rect -71547 -35168 -71443 -34932
rect -71207 -35168 -71103 -34932
rect -70867 -35168 -70783 -34932
rect -70547 -35168 -70443 -34932
rect -70207 -35168 -70103 -34932
rect -69867 -35168 -69783 -34932
rect -69547 -35168 -69443 -34932
rect -69207 -35168 -69103 -34932
rect -68867 -35168 -68783 -34932
rect -68547 -35168 -68443 -34932
rect -68207 -35168 -68103 -34932
rect -67867 -35168 -67783 -34932
rect -67547 -35168 -67443 -34932
rect -67207 -35168 -67103 -34932
rect -66867 -35168 -66783 -34932
rect -66547 -35168 -66443 -34932
rect -66207 -35168 -66103 -34932
rect -65867 -35168 -65783 -34932
rect -65547 -35168 -65443 -34932
rect -65207 -35168 -65103 -34932
rect -64867 -35168 -64783 -34932
rect -64547 -35168 -64443 -34932
rect -64207 -35168 -64103 -34932
rect -63867 -35168 -63783 -34932
rect -63547 -35168 -63443 -34932
rect -63207 -35168 -63103 -34932
rect -62867 -35168 -62783 -34932
rect -62547 -35168 -62443 -34932
rect -62207 -35168 -62103 -34932
rect -61867 -35168 -61783 -34932
rect -61547 -35168 -61443 -34932
rect -61207 -35168 -61103 -34932
rect -60867 -35168 -60783 -34932
rect -60547 -35168 -60443 -34932
rect -60207 -35168 -60103 -34932
rect -59867 -35168 -59783 -34932
rect -59547 -35168 -59443 -34932
rect -59207 -35168 -59103 -34932
rect -58867 -35168 -58783 -34932
rect -58547 -35168 -58443 -34932
rect -58207 -35168 -58103 -34932
rect -57867 -35168 -57783 -34932
rect -57547 -35168 -57443 -34932
rect -57207 -35168 -57103 -34932
rect -56867 -35168 -56783 -34932
rect -56547 -35168 -56443 -34932
rect -56207 -35168 -56103 -34932
rect -55867 -35168 -55783 -34932
rect -55547 -35168 -55443 -34932
rect -55207 -35168 -55103 -34932
rect -54867 -35168 -54783 -34932
rect -54547 -35168 -54443 -34932
rect -54207 -35168 -54103 -34932
rect -53867 -35168 -53783 -34932
rect -53547 -35168 -53443 -34932
rect -53207 -35168 -53103 -34932
rect -52867 -35168 -52783 -34932
rect -52547 -35168 -52443 -34932
rect -52207 -35168 -52103 -34932
rect -51867 -35168 -51783 -34932
rect -51547 -35168 -51443 -34932
rect -51207 -35168 -51103 -34932
rect -50867 -35168 -50783 -34932
rect -50547 -35168 -50443 -34932
rect -50207 -35168 -50103 -34932
rect -49867 -35168 -49783 -34932
rect -49547 -35168 -49443 -34932
rect -49207 -35168 -49103 -34932
rect -48867 -35168 -48825 -34932
rect -74825 -35210 -48825 -35168
rect -74485 -35272 -74165 -35210
rect -74485 -35508 -74443 -35272
rect -74207 -35508 -74165 -35272
rect -74485 -35592 -74165 -35508
rect -74485 -35828 -74443 -35592
rect -74207 -35828 -74165 -35592
rect -74485 -35890 -74165 -35828
rect -73485 -35272 -73165 -35210
rect -73485 -35508 -73443 -35272
rect -73207 -35508 -73165 -35272
rect -73485 -35592 -73165 -35508
rect -73485 -35828 -73443 -35592
rect -73207 -35828 -73165 -35592
rect -73485 -35890 -73165 -35828
rect -72485 -35272 -72165 -35210
rect -72485 -35508 -72443 -35272
rect -72207 -35508 -72165 -35272
rect -72485 -35592 -72165 -35508
rect -72485 -35828 -72443 -35592
rect -72207 -35828 -72165 -35592
rect -72485 -35890 -72165 -35828
rect -71485 -35272 -71165 -35210
rect -71485 -35508 -71443 -35272
rect -71207 -35508 -71165 -35272
rect -71485 -35592 -71165 -35508
rect -71485 -35828 -71443 -35592
rect -71207 -35828 -71165 -35592
rect -71485 -35890 -71165 -35828
rect -70485 -35272 -70165 -35210
rect -70485 -35508 -70443 -35272
rect -70207 -35508 -70165 -35272
rect -70485 -35592 -70165 -35508
rect -70485 -35828 -70443 -35592
rect -70207 -35828 -70165 -35592
rect -70485 -35890 -70165 -35828
rect -69485 -35272 -69165 -35210
rect -69485 -35508 -69443 -35272
rect -69207 -35508 -69165 -35272
rect -69485 -35592 -69165 -35508
rect -69485 -35828 -69443 -35592
rect -69207 -35828 -69165 -35592
rect -69485 -35890 -69165 -35828
rect -68485 -35272 -68165 -35210
rect -68485 -35508 -68443 -35272
rect -68207 -35508 -68165 -35272
rect -68485 -35592 -68165 -35508
rect -68485 -35828 -68443 -35592
rect -68207 -35828 -68165 -35592
rect -68485 -35890 -68165 -35828
rect -67485 -35272 -67165 -35210
rect -67485 -35508 -67443 -35272
rect -67207 -35508 -67165 -35272
rect -67485 -35592 -67165 -35508
rect -67485 -35828 -67443 -35592
rect -67207 -35828 -67165 -35592
rect -67485 -35890 -67165 -35828
rect -66485 -35272 -66165 -35210
rect -66485 -35508 -66443 -35272
rect -66207 -35508 -66165 -35272
rect -66485 -35592 -66165 -35508
rect -66485 -35828 -66443 -35592
rect -66207 -35828 -66165 -35592
rect -66485 -35890 -66165 -35828
rect -65485 -35272 -65165 -35210
rect -65485 -35508 -65443 -35272
rect -65207 -35508 -65165 -35272
rect -65485 -35592 -65165 -35508
rect -65485 -35828 -65443 -35592
rect -65207 -35828 -65165 -35592
rect -65485 -35890 -65165 -35828
rect -64485 -35272 -64165 -35210
rect -64485 -35508 -64443 -35272
rect -64207 -35508 -64165 -35272
rect -64485 -35592 -64165 -35508
rect -64485 -35828 -64443 -35592
rect -64207 -35828 -64165 -35592
rect -64485 -35890 -64165 -35828
rect -63485 -35272 -63165 -35210
rect -63485 -35508 -63443 -35272
rect -63207 -35508 -63165 -35272
rect -63485 -35592 -63165 -35508
rect -63485 -35828 -63443 -35592
rect -63207 -35828 -63165 -35592
rect -63485 -35890 -63165 -35828
rect -62485 -35272 -62165 -35210
rect -62485 -35508 -62443 -35272
rect -62207 -35508 -62165 -35272
rect -62485 -35592 -62165 -35508
rect -62485 -35828 -62443 -35592
rect -62207 -35828 -62165 -35592
rect -62485 -35890 -62165 -35828
rect -61485 -35272 -61165 -35210
rect -61485 -35508 -61443 -35272
rect -61207 -35508 -61165 -35272
rect -61485 -35592 -61165 -35508
rect -61485 -35828 -61443 -35592
rect -61207 -35828 -61165 -35592
rect -61485 -35890 -61165 -35828
rect -60485 -35272 -60165 -35210
rect -60485 -35508 -60443 -35272
rect -60207 -35508 -60165 -35272
rect -60485 -35592 -60165 -35508
rect -60485 -35828 -60443 -35592
rect -60207 -35828 -60165 -35592
rect -60485 -35890 -60165 -35828
rect -59485 -35272 -59165 -35210
rect -59485 -35508 -59443 -35272
rect -59207 -35508 -59165 -35272
rect -59485 -35592 -59165 -35508
rect -59485 -35828 -59443 -35592
rect -59207 -35828 -59165 -35592
rect -59485 -35890 -59165 -35828
rect -58485 -35272 -58165 -35210
rect -58485 -35508 -58443 -35272
rect -58207 -35508 -58165 -35272
rect -58485 -35592 -58165 -35508
rect -58485 -35828 -58443 -35592
rect -58207 -35828 -58165 -35592
rect -58485 -35890 -58165 -35828
rect -57485 -35272 -57165 -35210
rect -57485 -35508 -57443 -35272
rect -57207 -35508 -57165 -35272
rect -57485 -35592 -57165 -35508
rect -57485 -35828 -57443 -35592
rect -57207 -35828 -57165 -35592
rect -57485 -35890 -57165 -35828
rect -56485 -35272 -56165 -35210
rect -56485 -35508 -56443 -35272
rect -56207 -35508 -56165 -35272
rect -56485 -35592 -56165 -35508
rect -56485 -35828 -56443 -35592
rect -56207 -35828 -56165 -35592
rect -56485 -35890 -56165 -35828
rect -55485 -35272 -55165 -35210
rect -55485 -35508 -55443 -35272
rect -55207 -35508 -55165 -35272
rect -55485 -35592 -55165 -35508
rect -55485 -35828 -55443 -35592
rect -55207 -35828 -55165 -35592
rect -55485 -35890 -55165 -35828
rect -54485 -35272 -54165 -35210
rect -54485 -35508 -54443 -35272
rect -54207 -35508 -54165 -35272
rect -54485 -35592 -54165 -35508
rect -54485 -35828 -54443 -35592
rect -54207 -35828 -54165 -35592
rect -54485 -35890 -54165 -35828
rect -53485 -35272 -53165 -35210
rect -53485 -35508 -53443 -35272
rect -53207 -35508 -53165 -35272
rect -53485 -35592 -53165 -35508
rect -53485 -35828 -53443 -35592
rect -53207 -35828 -53165 -35592
rect -53485 -35890 -53165 -35828
rect -52485 -35272 -52165 -35210
rect -52485 -35508 -52443 -35272
rect -52207 -35508 -52165 -35272
rect -52485 -35592 -52165 -35508
rect -52485 -35828 -52443 -35592
rect -52207 -35828 -52165 -35592
rect -52485 -35890 -52165 -35828
rect -51485 -35272 -51165 -35210
rect -51485 -35508 -51443 -35272
rect -51207 -35508 -51165 -35272
rect -51485 -35592 -51165 -35508
rect -51485 -35828 -51443 -35592
rect -51207 -35828 -51165 -35592
rect -51485 -35890 -51165 -35828
rect -50485 -35272 -50165 -35210
rect -50485 -35508 -50443 -35272
rect -50207 -35508 -50165 -35272
rect -50485 -35592 -50165 -35508
rect -50485 -35828 -50443 -35592
rect -50207 -35828 -50165 -35592
rect -50485 -35890 -50165 -35828
rect -49485 -35272 -49165 -35210
rect -49485 -35508 -49443 -35272
rect -49207 -35508 -49165 -35272
rect -49485 -35592 -49165 -35508
rect -49485 -35828 -49443 -35592
rect -49207 -35828 -49165 -35592
rect -49485 -35890 -49165 -35828
rect -74825 -35932 -48825 -35890
rect -74825 -36168 -74783 -35932
rect -74547 -36168 -74443 -35932
rect -74207 -36168 -74103 -35932
rect -73867 -36168 -73783 -35932
rect -73547 -36168 -73443 -35932
rect -73207 -36168 -73103 -35932
rect -72867 -36168 -72783 -35932
rect -72547 -36168 -72443 -35932
rect -72207 -36168 -72103 -35932
rect -71867 -36168 -71783 -35932
rect -71547 -36168 -71443 -35932
rect -71207 -36168 -71103 -35932
rect -70867 -36168 -70783 -35932
rect -70547 -36168 -70443 -35932
rect -70207 -36168 -70103 -35932
rect -69867 -36168 -69783 -35932
rect -69547 -36168 -69443 -35932
rect -69207 -36168 -69103 -35932
rect -68867 -36168 -68783 -35932
rect -68547 -36168 -68443 -35932
rect -68207 -36168 -68103 -35932
rect -67867 -36168 -67783 -35932
rect -67547 -36168 -67443 -35932
rect -67207 -36168 -67103 -35932
rect -66867 -36168 -66783 -35932
rect -66547 -36168 -66443 -35932
rect -66207 -36168 -66103 -35932
rect -65867 -36168 -65783 -35932
rect -65547 -36168 -65443 -35932
rect -65207 -36168 -65103 -35932
rect -64867 -36168 -64783 -35932
rect -64547 -36168 -64443 -35932
rect -64207 -36168 -64103 -35932
rect -63867 -36168 -63783 -35932
rect -63547 -36168 -63443 -35932
rect -63207 -36168 -63103 -35932
rect -62867 -36168 -62783 -35932
rect -62547 -36168 -62443 -35932
rect -62207 -36168 -62103 -35932
rect -61867 -36168 -61783 -35932
rect -61547 -36168 -61443 -35932
rect -61207 -36168 -61103 -35932
rect -60867 -36168 -60783 -35932
rect -60547 -36168 -60443 -35932
rect -60207 -36168 -60103 -35932
rect -59867 -36168 -59783 -35932
rect -59547 -36168 -59443 -35932
rect -59207 -36168 -59103 -35932
rect -58867 -36168 -58783 -35932
rect -58547 -36168 -58443 -35932
rect -58207 -36168 -58103 -35932
rect -57867 -36168 -57783 -35932
rect -57547 -36168 -57443 -35932
rect -57207 -36168 -57103 -35932
rect -56867 -36168 -56783 -35932
rect -56547 -36168 -56443 -35932
rect -56207 -36168 -56103 -35932
rect -55867 -36168 -55783 -35932
rect -55547 -36168 -55443 -35932
rect -55207 -36168 -55103 -35932
rect -54867 -36168 -54783 -35932
rect -54547 -36168 -54443 -35932
rect -54207 -36168 -54103 -35932
rect -53867 -36168 -53783 -35932
rect -53547 -36168 -53443 -35932
rect -53207 -36168 -53103 -35932
rect -52867 -36168 -52783 -35932
rect -52547 -36168 -52443 -35932
rect -52207 -36168 -52103 -35932
rect -51867 -36168 -51783 -35932
rect -51547 -36168 -51443 -35932
rect -51207 -36168 -51103 -35932
rect -50867 -36168 -50783 -35932
rect -50547 -36168 -50443 -35932
rect -50207 -36168 -50103 -35932
rect -49867 -36168 -49783 -35932
rect -49547 -36168 -49443 -35932
rect -49207 -36168 -49103 -35932
rect -48867 -36168 -48825 -35932
rect -74825 -36210 -48825 -36168
rect -74485 -36272 -74165 -36210
rect -74485 -36508 -74443 -36272
rect -74207 -36508 -74165 -36272
rect -74485 -36592 -74165 -36508
rect -74485 -36828 -74443 -36592
rect -74207 -36828 -74165 -36592
rect -74485 -36890 -74165 -36828
rect -73485 -36272 -73165 -36210
rect -73485 -36508 -73443 -36272
rect -73207 -36508 -73165 -36272
rect -73485 -36592 -73165 -36508
rect -73485 -36828 -73443 -36592
rect -73207 -36828 -73165 -36592
rect -73485 -36890 -73165 -36828
rect -72485 -36272 -72165 -36210
rect -72485 -36508 -72443 -36272
rect -72207 -36508 -72165 -36272
rect -72485 -36592 -72165 -36508
rect -72485 -36828 -72443 -36592
rect -72207 -36828 -72165 -36592
rect -72485 -36890 -72165 -36828
rect -71485 -36272 -71165 -36210
rect -71485 -36508 -71443 -36272
rect -71207 -36508 -71165 -36272
rect -71485 -36592 -71165 -36508
rect -71485 -36828 -71443 -36592
rect -71207 -36828 -71165 -36592
rect -71485 -36890 -71165 -36828
rect -70485 -36272 -70165 -36210
rect -70485 -36508 -70443 -36272
rect -70207 -36508 -70165 -36272
rect -70485 -36592 -70165 -36508
rect -70485 -36828 -70443 -36592
rect -70207 -36828 -70165 -36592
rect -70485 -36890 -70165 -36828
rect -69485 -36272 -69165 -36210
rect -69485 -36508 -69443 -36272
rect -69207 -36508 -69165 -36272
rect -69485 -36592 -69165 -36508
rect -69485 -36828 -69443 -36592
rect -69207 -36828 -69165 -36592
rect -69485 -36890 -69165 -36828
rect -68485 -36272 -68165 -36210
rect -68485 -36508 -68443 -36272
rect -68207 -36508 -68165 -36272
rect -68485 -36592 -68165 -36508
rect -68485 -36828 -68443 -36592
rect -68207 -36828 -68165 -36592
rect -68485 -36890 -68165 -36828
rect -67485 -36272 -67165 -36210
rect -67485 -36508 -67443 -36272
rect -67207 -36508 -67165 -36272
rect -67485 -36592 -67165 -36508
rect -67485 -36828 -67443 -36592
rect -67207 -36828 -67165 -36592
rect -67485 -36890 -67165 -36828
rect -66485 -36272 -66165 -36210
rect -66485 -36508 -66443 -36272
rect -66207 -36508 -66165 -36272
rect -66485 -36592 -66165 -36508
rect -66485 -36828 -66443 -36592
rect -66207 -36828 -66165 -36592
rect -66485 -36890 -66165 -36828
rect -65485 -36272 -65165 -36210
rect -65485 -36508 -65443 -36272
rect -65207 -36508 -65165 -36272
rect -65485 -36592 -65165 -36508
rect -65485 -36828 -65443 -36592
rect -65207 -36828 -65165 -36592
rect -65485 -36890 -65165 -36828
rect -64485 -36272 -64165 -36210
rect -64485 -36508 -64443 -36272
rect -64207 -36508 -64165 -36272
rect -64485 -36592 -64165 -36508
rect -64485 -36828 -64443 -36592
rect -64207 -36828 -64165 -36592
rect -64485 -36890 -64165 -36828
rect -63485 -36272 -63165 -36210
rect -63485 -36508 -63443 -36272
rect -63207 -36508 -63165 -36272
rect -63485 -36592 -63165 -36508
rect -63485 -36828 -63443 -36592
rect -63207 -36828 -63165 -36592
rect -63485 -36890 -63165 -36828
rect -62485 -36272 -62165 -36210
rect -62485 -36508 -62443 -36272
rect -62207 -36508 -62165 -36272
rect -62485 -36592 -62165 -36508
rect -62485 -36828 -62443 -36592
rect -62207 -36828 -62165 -36592
rect -62485 -36890 -62165 -36828
rect -61485 -36272 -61165 -36210
rect -61485 -36508 -61443 -36272
rect -61207 -36508 -61165 -36272
rect -61485 -36592 -61165 -36508
rect -61485 -36828 -61443 -36592
rect -61207 -36828 -61165 -36592
rect -61485 -36890 -61165 -36828
rect -60485 -36272 -60165 -36210
rect -60485 -36508 -60443 -36272
rect -60207 -36508 -60165 -36272
rect -60485 -36592 -60165 -36508
rect -60485 -36828 -60443 -36592
rect -60207 -36828 -60165 -36592
rect -60485 -36890 -60165 -36828
rect -59485 -36272 -59165 -36210
rect -59485 -36508 -59443 -36272
rect -59207 -36508 -59165 -36272
rect -59485 -36592 -59165 -36508
rect -59485 -36828 -59443 -36592
rect -59207 -36828 -59165 -36592
rect -59485 -36890 -59165 -36828
rect -58485 -36272 -58165 -36210
rect -58485 -36508 -58443 -36272
rect -58207 -36508 -58165 -36272
rect -58485 -36592 -58165 -36508
rect -58485 -36828 -58443 -36592
rect -58207 -36828 -58165 -36592
rect -58485 -36890 -58165 -36828
rect -57485 -36272 -57165 -36210
rect -57485 -36508 -57443 -36272
rect -57207 -36508 -57165 -36272
rect -57485 -36592 -57165 -36508
rect -57485 -36828 -57443 -36592
rect -57207 -36828 -57165 -36592
rect -57485 -36890 -57165 -36828
rect -56485 -36272 -56165 -36210
rect -56485 -36508 -56443 -36272
rect -56207 -36508 -56165 -36272
rect -56485 -36592 -56165 -36508
rect -56485 -36828 -56443 -36592
rect -56207 -36828 -56165 -36592
rect -56485 -36890 -56165 -36828
rect -55485 -36272 -55165 -36210
rect -55485 -36508 -55443 -36272
rect -55207 -36508 -55165 -36272
rect -55485 -36592 -55165 -36508
rect -55485 -36828 -55443 -36592
rect -55207 -36828 -55165 -36592
rect -55485 -36890 -55165 -36828
rect -54485 -36272 -54165 -36210
rect -54485 -36508 -54443 -36272
rect -54207 -36508 -54165 -36272
rect -54485 -36592 -54165 -36508
rect -54485 -36828 -54443 -36592
rect -54207 -36828 -54165 -36592
rect -54485 -36890 -54165 -36828
rect -53485 -36272 -53165 -36210
rect -53485 -36508 -53443 -36272
rect -53207 -36508 -53165 -36272
rect -53485 -36592 -53165 -36508
rect -53485 -36828 -53443 -36592
rect -53207 -36828 -53165 -36592
rect -53485 -36890 -53165 -36828
rect -52485 -36272 -52165 -36210
rect -52485 -36508 -52443 -36272
rect -52207 -36508 -52165 -36272
rect -52485 -36592 -52165 -36508
rect -52485 -36828 -52443 -36592
rect -52207 -36828 -52165 -36592
rect -52485 -36890 -52165 -36828
rect -51485 -36272 -51165 -36210
rect -51485 -36508 -51443 -36272
rect -51207 -36508 -51165 -36272
rect -51485 -36592 -51165 -36508
rect -51485 -36828 -51443 -36592
rect -51207 -36828 -51165 -36592
rect -51485 -36890 -51165 -36828
rect -50485 -36272 -50165 -36210
rect -50485 -36508 -50443 -36272
rect -50207 -36508 -50165 -36272
rect -50485 -36592 -50165 -36508
rect -50485 -36828 -50443 -36592
rect -50207 -36828 -50165 -36592
rect -50485 -36890 -50165 -36828
rect -49485 -36272 -49165 -36210
rect -49485 -36508 -49443 -36272
rect -49207 -36508 -49165 -36272
rect -49485 -36592 -49165 -36508
rect -49485 -36828 -49443 -36592
rect -49207 -36828 -49165 -36592
rect -49485 -36890 -49165 -36828
rect -74825 -36932 -48825 -36890
rect -74825 -37168 -74783 -36932
rect -74547 -37168 -74443 -36932
rect -74207 -37168 -74103 -36932
rect -73867 -37168 -73783 -36932
rect -73547 -37168 -73443 -36932
rect -73207 -37168 -73103 -36932
rect -72867 -37168 -72783 -36932
rect -72547 -37168 -72443 -36932
rect -72207 -37168 -72103 -36932
rect -71867 -37168 -71783 -36932
rect -71547 -37168 -71443 -36932
rect -71207 -37168 -71103 -36932
rect -70867 -37168 -70783 -36932
rect -70547 -37168 -70443 -36932
rect -70207 -37168 -70103 -36932
rect -69867 -37168 -69783 -36932
rect -69547 -37168 -69443 -36932
rect -69207 -37168 -69103 -36932
rect -68867 -37168 -68783 -36932
rect -68547 -37168 -68443 -36932
rect -68207 -37168 -68103 -36932
rect -67867 -37168 -67783 -36932
rect -67547 -37168 -67443 -36932
rect -67207 -37168 -67103 -36932
rect -66867 -37168 -66783 -36932
rect -66547 -37168 -66443 -36932
rect -66207 -37168 -66103 -36932
rect -65867 -37168 -65783 -36932
rect -65547 -37168 -65443 -36932
rect -65207 -37168 -65103 -36932
rect -64867 -37168 -64783 -36932
rect -64547 -37168 -64443 -36932
rect -64207 -37168 -64103 -36932
rect -63867 -37168 -63783 -36932
rect -63547 -37168 -63443 -36932
rect -63207 -37168 -63103 -36932
rect -62867 -37168 -62783 -36932
rect -62547 -37168 -62443 -36932
rect -62207 -37168 -62103 -36932
rect -61867 -37168 -61783 -36932
rect -61547 -37168 -61443 -36932
rect -61207 -37168 -61103 -36932
rect -60867 -37168 -60783 -36932
rect -60547 -37168 -60443 -36932
rect -60207 -37168 -60103 -36932
rect -59867 -37168 -59783 -36932
rect -59547 -37168 -59443 -36932
rect -59207 -37168 -59103 -36932
rect -58867 -37168 -58783 -36932
rect -58547 -37168 -58443 -36932
rect -58207 -37168 -58103 -36932
rect -57867 -37168 -57783 -36932
rect -57547 -37168 -57443 -36932
rect -57207 -37168 -57103 -36932
rect -56867 -37168 -56783 -36932
rect -56547 -37168 -56443 -36932
rect -56207 -37168 -56103 -36932
rect -55867 -37168 -55783 -36932
rect -55547 -37168 -55443 -36932
rect -55207 -37168 -55103 -36932
rect -54867 -37168 -54783 -36932
rect -54547 -37168 -54443 -36932
rect -54207 -37168 -54103 -36932
rect -53867 -37168 -53783 -36932
rect -53547 -37168 -53443 -36932
rect -53207 -37168 -53103 -36932
rect -52867 -37168 -52783 -36932
rect -52547 -37168 -52443 -36932
rect -52207 -37168 -52103 -36932
rect -51867 -37168 -51783 -36932
rect -51547 -37168 -51443 -36932
rect -51207 -37168 -51103 -36932
rect -50867 -37168 -50783 -36932
rect -50547 -37168 -50443 -36932
rect -50207 -37168 -50103 -36932
rect -49867 -37168 -49783 -36932
rect -49547 -37168 -49443 -36932
rect -49207 -37168 -49103 -36932
rect -48867 -37168 -48825 -36932
rect -74825 -37210 -48825 -37168
rect -74485 -37272 -74165 -37210
rect -74485 -37508 -74443 -37272
rect -74207 -37508 -74165 -37272
rect -74485 -37592 -74165 -37508
rect -74485 -37828 -74443 -37592
rect -74207 -37828 -74165 -37592
rect -74485 -37890 -74165 -37828
rect -73485 -37272 -73165 -37210
rect -73485 -37508 -73443 -37272
rect -73207 -37508 -73165 -37272
rect -73485 -37592 -73165 -37508
rect -73485 -37828 -73443 -37592
rect -73207 -37828 -73165 -37592
rect -73485 -37890 -73165 -37828
rect -72485 -37272 -72165 -37210
rect -72485 -37508 -72443 -37272
rect -72207 -37508 -72165 -37272
rect -72485 -37592 -72165 -37508
rect -72485 -37828 -72443 -37592
rect -72207 -37828 -72165 -37592
rect -72485 -37890 -72165 -37828
rect -71485 -37272 -71165 -37210
rect -71485 -37508 -71443 -37272
rect -71207 -37508 -71165 -37272
rect -71485 -37592 -71165 -37508
rect -71485 -37828 -71443 -37592
rect -71207 -37828 -71165 -37592
rect -71485 -37890 -71165 -37828
rect -70485 -37272 -70165 -37210
rect -70485 -37508 -70443 -37272
rect -70207 -37508 -70165 -37272
rect -70485 -37592 -70165 -37508
rect -70485 -37828 -70443 -37592
rect -70207 -37828 -70165 -37592
rect -70485 -37890 -70165 -37828
rect -69485 -37272 -69165 -37210
rect -69485 -37508 -69443 -37272
rect -69207 -37508 -69165 -37272
rect -69485 -37592 -69165 -37508
rect -69485 -37828 -69443 -37592
rect -69207 -37828 -69165 -37592
rect -69485 -37890 -69165 -37828
rect -68485 -37272 -68165 -37210
rect -68485 -37508 -68443 -37272
rect -68207 -37508 -68165 -37272
rect -68485 -37592 -68165 -37508
rect -68485 -37828 -68443 -37592
rect -68207 -37828 -68165 -37592
rect -68485 -37890 -68165 -37828
rect -67485 -37272 -67165 -37210
rect -67485 -37508 -67443 -37272
rect -67207 -37508 -67165 -37272
rect -67485 -37592 -67165 -37508
rect -67485 -37828 -67443 -37592
rect -67207 -37828 -67165 -37592
rect -67485 -37890 -67165 -37828
rect -66485 -37272 -66165 -37210
rect -66485 -37508 -66443 -37272
rect -66207 -37508 -66165 -37272
rect -66485 -37592 -66165 -37508
rect -66485 -37828 -66443 -37592
rect -66207 -37828 -66165 -37592
rect -66485 -37890 -66165 -37828
rect -65485 -37272 -65165 -37210
rect -65485 -37508 -65443 -37272
rect -65207 -37508 -65165 -37272
rect -65485 -37592 -65165 -37508
rect -65485 -37828 -65443 -37592
rect -65207 -37828 -65165 -37592
rect -65485 -37890 -65165 -37828
rect -64485 -37272 -64165 -37210
rect -64485 -37508 -64443 -37272
rect -64207 -37508 -64165 -37272
rect -64485 -37592 -64165 -37508
rect -64485 -37828 -64443 -37592
rect -64207 -37828 -64165 -37592
rect -64485 -37890 -64165 -37828
rect -63485 -37272 -63165 -37210
rect -63485 -37508 -63443 -37272
rect -63207 -37508 -63165 -37272
rect -63485 -37592 -63165 -37508
rect -63485 -37828 -63443 -37592
rect -63207 -37828 -63165 -37592
rect -63485 -37890 -63165 -37828
rect -62485 -37272 -62165 -37210
rect -62485 -37508 -62443 -37272
rect -62207 -37508 -62165 -37272
rect -62485 -37592 -62165 -37508
rect -62485 -37828 -62443 -37592
rect -62207 -37828 -62165 -37592
rect -62485 -37890 -62165 -37828
rect -61485 -37272 -61165 -37210
rect -61485 -37508 -61443 -37272
rect -61207 -37508 -61165 -37272
rect -61485 -37592 -61165 -37508
rect -61485 -37828 -61443 -37592
rect -61207 -37828 -61165 -37592
rect -61485 -37890 -61165 -37828
rect -60485 -37272 -60165 -37210
rect -60485 -37508 -60443 -37272
rect -60207 -37508 -60165 -37272
rect -60485 -37592 -60165 -37508
rect -60485 -37828 -60443 -37592
rect -60207 -37828 -60165 -37592
rect -60485 -37890 -60165 -37828
rect -59485 -37272 -59165 -37210
rect -59485 -37508 -59443 -37272
rect -59207 -37508 -59165 -37272
rect -59485 -37592 -59165 -37508
rect -59485 -37828 -59443 -37592
rect -59207 -37828 -59165 -37592
rect -59485 -37890 -59165 -37828
rect -58485 -37272 -58165 -37210
rect -58485 -37508 -58443 -37272
rect -58207 -37508 -58165 -37272
rect -58485 -37592 -58165 -37508
rect -58485 -37828 -58443 -37592
rect -58207 -37828 -58165 -37592
rect -58485 -37890 -58165 -37828
rect -57485 -37272 -57165 -37210
rect -57485 -37508 -57443 -37272
rect -57207 -37508 -57165 -37272
rect -57485 -37592 -57165 -37508
rect -57485 -37828 -57443 -37592
rect -57207 -37828 -57165 -37592
rect -57485 -37890 -57165 -37828
rect -56485 -37272 -56165 -37210
rect -56485 -37508 -56443 -37272
rect -56207 -37508 -56165 -37272
rect -56485 -37592 -56165 -37508
rect -56485 -37828 -56443 -37592
rect -56207 -37828 -56165 -37592
rect -56485 -37890 -56165 -37828
rect -55485 -37272 -55165 -37210
rect -55485 -37508 -55443 -37272
rect -55207 -37508 -55165 -37272
rect -55485 -37592 -55165 -37508
rect -55485 -37828 -55443 -37592
rect -55207 -37828 -55165 -37592
rect -55485 -37890 -55165 -37828
rect -54485 -37272 -54165 -37210
rect -54485 -37508 -54443 -37272
rect -54207 -37508 -54165 -37272
rect -54485 -37592 -54165 -37508
rect -54485 -37828 -54443 -37592
rect -54207 -37828 -54165 -37592
rect -54485 -37890 -54165 -37828
rect -53485 -37272 -53165 -37210
rect -53485 -37508 -53443 -37272
rect -53207 -37508 -53165 -37272
rect -53485 -37592 -53165 -37508
rect -53485 -37828 -53443 -37592
rect -53207 -37828 -53165 -37592
rect -53485 -37890 -53165 -37828
rect -52485 -37272 -52165 -37210
rect -52485 -37508 -52443 -37272
rect -52207 -37508 -52165 -37272
rect -52485 -37592 -52165 -37508
rect -52485 -37828 -52443 -37592
rect -52207 -37828 -52165 -37592
rect -52485 -37890 -52165 -37828
rect -51485 -37272 -51165 -37210
rect -51485 -37508 -51443 -37272
rect -51207 -37508 -51165 -37272
rect -51485 -37592 -51165 -37508
rect -51485 -37828 -51443 -37592
rect -51207 -37828 -51165 -37592
rect -51485 -37890 -51165 -37828
rect -50485 -37272 -50165 -37210
rect -50485 -37508 -50443 -37272
rect -50207 -37508 -50165 -37272
rect -50485 -37592 -50165 -37508
rect -50485 -37828 -50443 -37592
rect -50207 -37828 -50165 -37592
rect -50485 -37890 -50165 -37828
rect -49485 -37272 -49165 -37210
rect -49485 -37508 -49443 -37272
rect -49207 -37508 -49165 -37272
rect -49485 -37592 -49165 -37508
rect -49485 -37828 -49443 -37592
rect -49207 -37828 -49165 -37592
rect -49485 -37890 -49165 -37828
rect -74825 -37932 -48825 -37890
rect -74825 -38168 -74783 -37932
rect -74547 -38168 -74443 -37932
rect -74207 -38168 -74103 -37932
rect -73867 -38168 -73783 -37932
rect -73547 -38168 -73443 -37932
rect -73207 -38168 -73103 -37932
rect -72867 -38168 -72783 -37932
rect -72547 -38168 -72443 -37932
rect -72207 -38168 -72103 -37932
rect -71867 -38168 -71783 -37932
rect -71547 -38168 -71443 -37932
rect -71207 -38168 -71103 -37932
rect -70867 -38168 -70783 -37932
rect -70547 -38168 -70443 -37932
rect -70207 -38168 -70103 -37932
rect -69867 -38168 -69783 -37932
rect -69547 -38168 -69443 -37932
rect -69207 -38168 -69103 -37932
rect -68867 -38168 -68783 -37932
rect -68547 -38168 -68443 -37932
rect -68207 -38168 -68103 -37932
rect -67867 -38168 -67783 -37932
rect -67547 -38168 -67443 -37932
rect -67207 -38168 -67103 -37932
rect -66867 -38168 -66783 -37932
rect -66547 -38168 -66443 -37932
rect -66207 -38168 -66103 -37932
rect -65867 -38168 -65783 -37932
rect -65547 -38168 -65443 -37932
rect -65207 -38168 -65103 -37932
rect -64867 -38168 -64783 -37932
rect -64547 -38168 -64443 -37932
rect -64207 -38168 -64103 -37932
rect -63867 -38168 -63783 -37932
rect -63547 -38168 -63443 -37932
rect -63207 -38168 -63103 -37932
rect -62867 -38168 -62783 -37932
rect -62547 -38168 -62443 -37932
rect -62207 -38168 -62103 -37932
rect -61867 -38168 -61783 -37932
rect -61547 -38168 -61443 -37932
rect -61207 -38168 -61103 -37932
rect -60867 -38168 -60783 -37932
rect -60547 -38168 -60443 -37932
rect -60207 -38168 -60103 -37932
rect -59867 -38168 -59783 -37932
rect -59547 -38168 -59443 -37932
rect -59207 -38168 -59103 -37932
rect -58867 -38168 -58783 -37932
rect -58547 -38168 -58443 -37932
rect -58207 -38168 -58103 -37932
rect -57867 -38168 -57783 -37932
rect -57547 -38168 -57443 -37932
rect -57207 -38168 -57103 -37932
rect -56867 -38168 -56783 -37932
rect -56547 -38168 -56443 -37932
rect -56207 -38168 -56103 -37932
rect -55867 -38168 -55783 -37932
rect -55547 -38168 -55443 -37932
rect -55207 -38168 -55103 -37932
rect -54867 -38168 -54783 -37932
rect -54547 -38168 -54443 -37932
rect -54207 -38168 -54103 -37932
rect -53867 -38168 -53783 -37932
rect -53547 -38168 -53443 -37932
rect -53207 -38168 -53103 -37932
rect -52867 -38168 -52783 -37932
rect -52547 -38168 -52443 -37932
rect -52207 -38168 -52103 -37932
rect -51867 -38168 -51783 -37932
rect -51547 -38168 -51443 -37932
rect -51207 -38168 -51103 -37932
rect -50867 -38168 -50783 -37932
rect -50547 -38168 -50443 -37932
rect -50207 -38168 -50103 -37932
rect -49867 -38168 -49783 -37932
rect -49547 -38168 -49443 -37932
rect -49207 -38168 -49103 -37932
rect -48867 -38168 -48825 -37932
rect -74825 -38210 -48825 -38168
rect -74485 -38272 -74165 -38210
rect -74485 -38508 -74443 -38272
rect -74207 -38508 -74165 -38272
rect -74485 -38592 -74165 -38508
rect -74485 -38828 -74443 -38592
rect -74207 -38828 -74165 -38592
rect -74485 -38890 -74165 -38828
rect -73485 -38272 -73165 -38210
rect -73485 -38508 -73443 -38272
rect -73207 -38508 -73165 -38272
rect -73485 -38592 -73165 -38508
rect -73485 -38828 -73443 -38592
rect -73207 -38828 -73165 -38592
rect -73485 -38890 -73165 -38828
rect -72485 -38272 -72165 -38210
rect -72485 -38508 -72443 -38272
rect -72207 -38508 -72165 -38272
rect -72485 -38592 -72165 -38508
rect -72485 -38828 -72443 -38592
rect -72207 -38828 -72165 -38592
rect -72485 -38890 -72165 -38828
rect -71485 -38272 -71165 -38210
rect -71485 -38508 -71443 -38272
rect -71207 -38508 -71165 -38272
rect -71485 -38592 -71165 -38508
rect -71485 -38828 -71443 -38592
rect -71207 -38828 -71165 -38592
rect -71485 -38890 -71165 -38828
rect -70485 -38272 -70165 -38210
rect -70485 -38508 -70443 -38272
rect -70207 -38508 -70165 -38272
rect -70485 -38592 -70165 -38508
rect -70485 -38828 -70443 -38592
rect -70207 -38828 -70165 -38592
rect -70485 -38890 -70165 -38828
rect -69485 -38272 -69165 -38210
rect -69485 -38508 -69443 -38272
rect -69207 -38508 -69165 -38272
rect -69485 -38592 -69165 -38508
rect -69485 -38828 -69443 -38592
rect -69207 -38828 -69165 -38592
rect -69485 -38890 -69165 -38828
rect -68485 -38272 -68165 -38210
rect -68485 -38508 -68443 -38272
rect -68207 -38508 -68165 -38272
rect -68485 -38592 -68165 -38508
rect -68485 -38828 -68443 -38592
rect -68207 -38828 -68165 -38592
rect -68485 -38890 -68165 -38828
rect -67485 -38272 -67165 -38210
rect -67485 -38508 -67443 -38272
rect -67207 -38508 -67165 -38272
rect -67485 -38592 -67165 -38508
rect -67485 -38828 -67443 -38592
rect -67207 -38828 -67165 -38592
rect -67485 -38890 -67165 -38828
rect -66485 -38272 -66165 -38210
rect -66485 -38508 -66443 -38272
rect -66207 -38508 -66165 -38272
rect -66485 -38592 -66165 -38508
rect -66485 -38828 -66443 -38592
rect -66207 -38828 -66165 -38592
rect -66485 -38890 -66165 -38828
rect -65485 -38272 -65165 -38210
rect -65485 -38508 -65443 -38272
rect -65207 -38508 -65165 -38272
rect -65485 -38592 -65165 -38508
rect -65485 -38828 -65443 -38592
rect -65207 -38828 -65165 -38592
rect -65485 -38890 -65165 -38828
rect -64485 -38272 -64165 -38210
rect -64485 -38508 -64443 -38272
rect -64207 -38508 -64165 -38272
rect -64485 -38592 -64165 -38508
rect -64485 -38828 -64443 -38592
rect -64207 -38828 -64165 -38592
rect -64485 -38890 -64165 -38828
rect -63485 -38272 -63165 -38210
rect -63485 -38508 -63443 -38272
rect -63207 -38508 -63165 -38272
rect -63485 -38592 -63165 -38508
rect -63485 -38828 -63443 -38592
rect -63207 -38828 -63165 -38592
rect -63485 -38890 -63165 -38828
rect -62485 -38272 -62165 -38210
rect -62485 -38508 -62443 -38272
rect -62207 -38508 -62165 -38272
rect -62485 -38592 -62165 -38508
rect -62485 -38828 -62443 -38592
rect -62207 -38828 -62165 -38592
rect -62485 -38890 -62165 -38828
rect -61485 -38272 -61165 -38210
rect -61485 -38508 -61443 -38272
rect -61207 -38508 -61165 -38272
rect -61485 -38592 -61165 -38508
rect -61485 -38828 -61443 -38592
rect -61207 -38828 -61165 -38592
rect -61485 -38890 -61165 -38828
rect -60485 -38272 -60165 -38210
rect -60485 -38508 -60443 -38272
rect -60207 -38508 -60165 -38272
rect -60485 -38592 -60165 -38508
rect -60485 -38828 -60443 -38592
rect -60207 -38828 -60165 -38592
rect -60485 -38890 -60165 -38828
rect -59485 -38272 -59165 -38210
rect -59485 -38508 -59443 -38272
rect -59207 -38508 -59165 -38272
rect -59485 -38592 -59165 -38508
rect -59485 -38828 -59443 -38592
rect -59207 -38828 -59165 -38592
rect -59485 -38890 -59165 -38828
rect -58485 -38272 -58165 -38210
rect -58485 -38508 -58443 -38272
rect -58207 -38508 -58165 -38272
rect -58485 -38592 -58165 -38508
rect -58485 -38828 -58443 -38592
rect -58207 -38828 -58165 -38592
rect -58485 -38890 -58165 -38828
rect -57485 -38272 -57165 -38210
rect -57485 -38508 -57443 -38272
rect -57207 -38508 -57165 -38272
rect -57485 -38592 -57165 -38508
rect -57485 -38828 -57443 -38592
rect -57207 -38828 -57165 -38592
rect -57485 -38890 -57165 -38828
rect -56485 -38272 -56165 -38210
rect -56485 -38508 -56443 -38272
rect -56207 -38508 -56165 -38272
rect -56485 -38592 -56165 -38508
rect -56485 -38828 -56443 -38592
rect -56207 -38828 -56165 -38592
rect -56485 -38890 -56165 -38828
rect -55485 -38272 -55165 -38210
rect -55485 -38508 -55443 -38272
rect -55207 -38508 -55165 -38272
rect -55485 -38592 -55165 -38508
rect -55485 -38828 -55443 -38592
rect -55207 -38828 -55165 -38592
rect -55485 -38890 -55165 -38828
rect -54485 -38272 -54165 -38210
rect -54485 -38508 -54443 -38272
rect -54207 -38508 -54165 -38272
rect -54485 -38592 -54165 -38508
rect -54485 -38828 -54443 -38592
rect -54207 -38828 -54165 -38592
rect -54485 -38890 -54165 -38828
rect -53485 -38272 -53165 -38210
rect -53485 -38508 -53443 -38272
rect -53207 -38508 -53165 -38272
rect -53485 -38592 -53165 -38508
rect -53485 -38828 -53443 -38592
rect -53207 -38828 -53165 -38592
rect -53485 -38890 -53165 -38828
rect -52485 -38272 -52165 -38210
rect -52485 -38508 -52443 -38272
rect -52207 -38508 -52165 -38272
rect -52485 -38592 -52165 -38508
rect -52485 -38828 -52443 -38592
rect -52207 -38828 -52165 -38592
rect -52485 -38890 -52165 -38828
rect -51485 -38272 -51165 -38210
rect -51485 -38508 -51443 -38272
rect -51207 -38508 -51165 -38272
rect -51485 -38592 -51165 -38508
rect -51485 -38828 -51443 -38592
rect -51207 -38828 -51165 -38592
rect -51485 -38890 -51165 -38828
rect -50485 -38272 -50165 -38210
rect -50485 -38508 -50443 -38272
rect -50207 -38508 -50165 -38272
rect -50485 -38592 -50165 -38508
rect -50485 -38828 -50443 -38592
rect -50207 -38828 -50165 -38592
rect -50485 -38890 -50165 -38828
rect -49485 -38272 -49165 -38210
rect -49485 -38508 -49443 -38272
rect -49207 -38508 -49165 -38272
rect -49485 -38592 -49165 -38508
rect -49485 -38828 -49443 -38592
rect -49207 -38828 -49165 -38592
rect -49485 -38890 -49165 -38828
rect -74825 -38932 -48825 -38890
rect -74825 -39168 -74783 -38932
rect -74547 -39168 -74443 -38932
rect -74207 -39168 -74103 -38932
rect -73867 -39168 -73783 -38932
rect -73547 -39168 -73443 -38932
rect -73207 -39168 -73103 -38932
rect -72867 -39168 -72783 -38932
rect -72547 -39168 -72443 -38932
rect -72207 -39168 -72103 -38932
rect -71867 -39168 -71783 -38932
rect -71547 -39168 -71443 -38932
rect -71207 -39168 -71103 -38932
rect -70867 -39168 -70783 -38932
rect -70547 -39168 -70443 -38932
rect -70207 -39168 -70103 -38932
rect -69867 -39168 -69783 -38932
rect -69547 -39168 -69443 -38932
rect -69207 -39168 -69103 -38932
rect -68867 -39168 -68783 -38932
rect -68547 -39168 -68443 -38932
rect -68207 -39168 -68103 -38932
rect -67867 -39168 -67783 -38932
rect -67547 -39168 -67443 -38932
rect -67207 -39168 -67103 -38932
rect -66867 -39168 -66783 -38932
rect -66547 -39168 -66443 -38932
rect -66207 -39168 -66103 -38932
rect -65867 -39168 -65783 -38932
rect -65547 -39168 -65443 -38932
rect -65207 -39168 -65103 -38932
rect -64867 -39168 -64783 -38932
rect -64547 -39168 -64443 -38932
rect -64207 -39168 -64103 -38932
rect -63867 -39168 -63783 -38932
rect -63547 -39168 -63443 -38932
rect -63207 -39168 -63103 -38932
rect -62867 -39168 -62783 -38932
rect -62547 -39168 -62443 -38932
rect -62207 -39168 -62103 -38932
rect -61867 -39168 -61783 -38932
rect -61547 -39168 -61443 -38932
rect -61207 -39168 -61103 -38932
rect -60867 -39168 -60783 -38932
rect -60547 -39168 -60443 -38932
rect -60207 -39168 -60103 -38932
rect -59867 -39168 -59783 -38932
rect -59547 -39168 -59443 -38932
rect -59207 -39168 -59103 -38932
rect -58867 -39168 -58783 -38932
rect -58547 -39168 -58443 -38932
rect -58207 -39168 -58103 -38932
rect -57867 -39168 -57783 -38932
rect -57547 -39168 -57443 -38932
rect -57207 -39168 -57103 -38932
rect -56867 -39168 -56783 -38932
rect -56547 -39168 -56443 -38932
rect -56207 -39168 -56103 -38932
rect -55867 -39168 -55783 -38932
rect -55547 -39168 -55443 -38932
rect -55207 -39168 -55103 -38932
rect -54867 -39168 -54783 -38932
rect -54547 -39168 -54443 -38932
rect -54207 -39168 -54103 -38932
rect -53867 -39168 -53783 -38932
rect -53547 -39168 -53443 -38932
rect -53207 -39168 -53103 -38932
rect -52867 -39168 -52783 -38932
rect -52547 -39168 -52443 -38932
rect -52207 -39168 -52103 -38932
rect -51867 -39168 -51783 -38932
rect -51547 -39168 -51443 -38932
rect -51207 -39168 -51103 -38932
rect -50867 -39168 -50783 -38932
rect -50547 -39168 -50443 -38932
rect -50207 -39168 -50103 -38932
rect -49867 -39168 -49783 -38932
rect -49547 -39168 -49443 -38932
rect -49207 -39168 -49103 -38932
rect -48867 -39168 -48825 -38932
rect -74825 -39210 -48825 -39168
rect -74485 -39272 -74165 -39210
rect -74485 -39508 -74443 -39272
rect -74207 -39508 -74165 -39272
rect -74485 -39592 -74165 -39508
rect -74485 -39828 -74443 -39592
rect -74207 -39828 -74165 -39592
rect -74485 -39890 -74165 -39828
rect -73485 -39272 -73165 -39210
rect -73485 -39508 -73443 -39272
rect -73207 -39508 -73165 -39272
rect -73485 -39592 -73165 -39508
rect -73485 -39828 -73443 -39592
rect -73207 -39828 -73165 -39592
rect -73485 -39890 -73165 -39828
rect -72485 -39272 -72165 -39210
rect -72485 -39508 -72443 -39272
rect -72207 -39508 -72165 -39272
rect -72485 -39592 -72165 -39508
rect -72485 -39828 -72443 -39592
rect -72207 -39828 -72165 -39592
rect -72485 -39890 -72165 -39828
rect -71485 -39272 -71165 -39210
rect -71485 -39508 -71443 -39272
rect -71207 -39508 -71165 -39272
rect -71485 -39592 -71165 -39508
rect -71485 -39828 -71443 -39592
rect -71207 -39828 -71165 -39592
rect -71485 -39890 -71165 -39828
rect -70485 -39272 -70165 -39210
rect -70485 -39508 -70443 -39272
rect -70207 -39508 -70165 -39272
rect -70485 -39592 -70165 -39508
rect -70485 -39828 -70443 -39592
rect -70207 -39828 -70165 -39592
rect -70485 -39890 -70165 -39828
rect -69485 -39272 -69165 -39210
rect -69485 -39508 -69443 -39272
rect -69207 -39508 -69165 -39272
rect -69485 -39592 -69165 -39508
rect -69485 -39828 -69443 -39592
rect -69207 -39828 -69165 -39592
rect -69485 -39890 -69165 -39828
rect -68485 -39272 -68165 -39210
rect -68485 -39508 -68443 -39272
rect -68207 -39508 -68165 -39272
rect -68485 -39592 -68165 -39508
rect -68485 -39828 -68443 -39592
rect -68207 -39828 -68165 -39592
rect -68485 -39890 -68165 -39828
rect -67485 -39272 -67165 -39210
rect -67485 -39508 -67443 -39272
rect -67207 -39508 -67165 -39272
rect -67485 -39592 -67165 -39508
rect -67485 -39828 -67443 -39592
rect -67207 -39828 -67165 -39592
rect -67485 -39890 -67165 -39828
rect -66485 -39272 -66165 -39210
rect -66485 -39508 -66443 -39272
rect -66207 -39508 -66165 -39272
rect -66485 -39592 -66165 -39508
rect -66485 -39828 -66443 -39592
rect -66207 -39828 -66165 -39592
rect -66485 -39890 -66165 -39828
rect -65485 -39272 -65165 -39210
rect -65485 -39508 -65443 -39272
rect -65207 -39508 -65165 -39272
rect -65485 -39592 -65165 -39508
rect -65485 -39828 -65443 -39592
rect -65207 -39828 -65165 -39592
rect -65485 -39890 -65165 -39828
rect -64485 -39272 -64165 -39210
rect -64485 -39508 -64443 -39272
rect -64207 -39508 -64165 -39272
rect -64485 -39592 -64165 -39508
rect -64485 -39828 -64443 -39592
rect -64207 -39828 -64165 -39592
rect -64485 -39890 -64165 -39828
rect -63485 -39272 -63165 -39210
rect -63485 -39508 -63443 -39272
rect -63207 -39508 -63165 -39272
rect -63485 -39592 -63165 -39508
rect -63485 -39828 -63443 -39592
rect -63207 -39828 -63165 -39592
rect -63485 -39890 -63165 -39828
rect -62485 -39272 -62165 -39210
rect -62485 -39508 -62443 -39272
rect -62207 -39508 -62165 -39272
rect -62485 -39592 -62165 -39508
rect -62485 -39828 -62443 -39592
rect -62207 -39828 -62165 -39592
rect -62485 -39890 -62165 -39828
rect -61485 -39272 -61165 -39210
rect -61485 -39508 -61443 -39272
rect -61207 -39508 -61165 -39272
rect -61485 -39592 -61165 -39508
rect -61485 -39828 -61443 -39592
rect -61207 -39828 -61165 -39592
rect -61485 -39890 -61165 -39828
rect -60485 -39272 -60165 -39210
rect -60485 -39508 -60443 -39272
rect -60207 -39508 -60165 -39272
rect -60485 -39592 -60165 -39508
rect -60485 -39828 -60443 -39592
rect -60207 -39828 -60165 -39592
rect -60485 -39890 -60165 -39828
rect -59485 -39272 -59165 -39210
rect -59485 -39508 -59443 -39272
rect -59207 -39508 -59165 -39272
rect -59485 -39592 -59165 -39508
rect -59485 -39828 -59443 -39592
rect -59207 -39828 -59165 -39592
rect -59485 -39890 -59165 -39828
rect -58485 -39272 -58165 -39210
rect -58485 -39508 -58443 -39272
rect -58207 -39508 -58165 -39272
rect -58485 -39592 -58165 -39508
rect -58485 -39828 -58443 -39592
rect -58207 -39828 -58165 -39592
rect -58485 -39890 -58165 -39828
rect -57485 -39272 -57165 -39210
rect -57485 -39508 -57443 -39272
rect -57207 -39508 -57165 -39272
rect -57485 -39592 -57165 -39508
rect -57485 -39828 -57443 -39592
rect -57207 -39828 -57165 -39592
rect -57485 -39890 -57165 -39828
rect -56485 -39272 -56165 -39210
rect -56485 -39508 -56443 -39272
rect -56207 -39508 -56165 -39272
rect -56485 -39592 -56165 -39508
rect -56485 -39828 -56443 -39592
rect -56207 -39828 -56165 -39592
rect -56485 -39890 -56165 -39828
rect -55485 -39272 -55165 -39210
rect -55485 -39508 -55443 -39272
rect -55207 -39508 -55165 -39272
rect -55485 -39592 -55165 -39508
rect -55485 -39828 -55443 -39592
rect -55207 -39828 -55165 -39592
rect -55485 -39890 -55165 -39828
rect -54485 -39272 -54165 -39210
rect -54485 -39508 -54443 -39272
rect -54207 -39508 -54165 -39272
rect -54485 -39592 -54165 -39508
rect -54485 -39828 -54443 -39592
rect -54207 -39828 -54165 -39592
rect -54485 -39890 -54165 -39828
rect -53485 -39272 -53165 -39210
rect -53485 -39508 -53443 -39272
rect -53207 -39508 -53165 -39272
rect -53485 -39592 -53165 -39508
rect -53485 -39828 -53443 -39592
rect -53207 -39828 -53165 -39592
rect -53485 -39890 -53165 -39828
rect -52485 -39272 -52165 -39210
rect -52485 -39508 -52443 -39272
rect -52207 -39508 -52165 -39272
rect -52485 -39592 -52165 -39508
rect -52485 -39828 -52443 -39592
rect -52207 -39828 -52165 -39592
rect -52485 -39890 -52165 -39828
rect -51485 -39272 -51165 -39210
rect -51485 -39508 -51443 -39272
rect -51207 -39508 -51165 -39272
rect -51485 -39592 -51165 -39508
rect -51485 -39828 -51443 -39592
rect -51207 -39828 -51165 -39592
rect -51485 -39890 -51165 -39828
rect -50485 -39272 -50165 -39210
rect -50485 -39508 -50443 -39272
rect -50207 -39508 -50165 -39272
rect -50485 -39592 -50165 -39508
rect -50485 -39828 -50443 -39592
rect -50207 -39828 -50165 -39592
rect -50485 -39890 -50165 -39828
rect -49485 -39272 -49165 -39210
rect -49485 -39508 -49443 -39272
rect -49207 -39508 -49165 -39272
rect -49485 -39592 -49165 -39508
rect -49485 -39828 -49443 -39592
rect -49207 -39828 -49165 -39592
rect -49485 -39890 -49165 -39828
rect -74825 -39932 -48825 -39890
rect -74825 -40168 -74783 -39932
rect -74547 -40168 -74443 -39932
rect -74207 -40168 -74103 -39932
rect -73867 -40168 -73783 -39932
rect -73547 -40168 -73443 -39932
rect -73207 -40168 -73103 -39932
rect -72867 -40168 -72783 -39932
rect -72547 -40168 -72443 -39932
rect -72207 -40168 -72103 -39932
rect -71867 -40168 -71783 -39932
rect -71547 -40168 -71443 -39932
rect -71207 -40168 -71103 -39932
rect -70867 -40168 -70783 -39932
rect -70547 -40168 -70443 -39932
rect -70207 -40168 -70103 -39932
rect -69867 -40168 -69783 -39932
rect -69547 -40168 -69443 -39932
rect -69207 -40168 -69103 -39932
rect -68867 -40168 -68783 -39932
rect -68547 -40168 -68443 -39932
rect -68207 -40168 -68103 -39932
rect -67867 -40168 -67783 -39932
rect -67547 -40168 -67443 -39932
rect -67207 -40168 -67103 -39932
rect -66867 -40168 -66783 -39932
rect -66547 -40168 -66443 -39932
rect -66207 -40168 -66103 -39932
rect -65867 -40168 -65783 -39932
rect -65547 -40168 -65443 -39932
rect -65207 -40168 -65103 -39932
rect -64867 -40168 -64783 -39932
rect -64547 -40168 -64443 -39932
rect -64207 -40168 -64103 -39932
rect -63867 -40168 -63783 -39932
rect -63547 -40168 -63443 -39932
rect -63207 -40168 -63103 -39932
rect -62867 -40168 -62783 -39932
rect -62547 -40168 -62443 -39932
rect -62207 -40168 -62103 -39932
rect -61867 -40168 -61783 -39932
rect -61547 -40168 -61443 -39932
rect -61207 -40168 -61103 -39932
rect -60867 -40168 -60783 -39932
rect -60547 -40168 -60443 -39932
rect -60207 -40168 -60103 -39932
rect -59867 -40168 -59783 -39932
rect -59547 -40168 -59443 -39932
rect -59207 -40168 -59103 -39932
rect -58867 -40168 -58783 -39932
rect -58547 -40168 -58443 -39932
rect -58207 -40168 -58103 -39932
rect -57867 -40168 -57783 -39932
rect -57547 -40168 -57443 -39932
rect -57207 -40168 -57103 -39932
rect -56867 -40168 -56783 -39932
rect -56547 -40168 -56443 -39932
rect -56207 -40168 -56103 -39932
rect -55867 -40168 -55783 -39932
rect -55547 -40168 -55443 -39932
rect -55207 -40168 -55103 -39932
rect -54867 -40168 -54783 -39932
rect -54547 -40168 -54443 -39932
rect -54207 -40168 -54103 -39932
rect -53867 -40168 -53783 -39932
rect -53547 -40168 -53443 -39932
rect -53207 -40168 -53103 -39932
rect -52867 -40168 -52783 -39932
rect -52547 -40168 -52443 -39932
rect -52207 -40168 -52103 -39932
rect -51867 -40168 -51783 -39932
rect -51547 -40168 -51443 -39932
rect -51207 -40168 -51103 -39932
rect -50867 -40168 -50783 -39932
rect -50547 -40168 -50443 -39932
rect -50207 -40168 -50103 -39932
rect -49867 -40168 -49783 -39932
rect -49547 -40168 -49443 -39932
rect -49207 -40168 -49103 -39932
rect -48867 -40168 -48825 -39932
rect -74825 -40210 -48825 -40168
rect -74485 -40272 -74165 -40210
rect -74485 -40508 -74443 -40272
rect -74207 -40508 -74165 -40272
rect -74485 -40592 -74165 -40508
rect -74485 -40828 -74443 -40592
rect -74207 -40828 -74165 -40592
rect -74485 -40890 -74165 -40828
rect -73485 -40272 -73165 -40210
rect -73485 -40508 -73443 -40272
rect -73207 -40508 -73165 -40272
rect -73485 -40592 -73165 -40508
rect -73485 -40828 -73443 -40592
rect -73207 -40828 -73165 -40592
rect -73485 -40890 -73165 -40828
rect -72485 -40272 -72165 -40210
rect -72485 -40508 -72443 -40272
rect -72207 -40508 -72165 -40272
rect -72485 -40592 -72165 -40508
rect -72485 -40828 -72443 -40592
rect -72207 -40828 -72165 -40592
rect -72485 -40890 -72165 -40828
rect -71485 -40272 -71165 -40210
rect -71485 -40508 -71443 -40272
rect -71207 -40508 -71165 -40272
rect -71485 -40592 -71165 -40508
rect -71485 -40828 -71443 -40592
rect -71207 -40828 -71165 -40592
rect -71485 -40890 -71165 -40828
rect -70485 -40272 -70165 -40210
rect -70485 -40508 -70443 -40272
rect -70207 -40508 -70165 -40272
rect -70485 -40592 -70165 -40508
rect -70485 -40828 -70443 -40592
rect -70207 -40828 -70165 -40592
rect -70485 -40890 -70165 -40828
rect -69485 -40272 -69165 -40210
rect -69485 -40508 -69443 -40272
rect -69207 -40508 -69165 -40272
rect -69485 -40592 -69165 -40508
rect -69485 -40828 -69443 -40592
rect -69207 -40828 -69165 -40592
rect -69485 -40890 -69165 -40828
rect -68485 -40272 -68165 -40210
rect -68485 -40508 -68443 -40272
rect -68207 -40508 -68165 -40272
rect -68485 -40592 -68165 -40508
rect -68485 -40828 -68443 -40592
rect -68207 -40828 -68165 -40592
rect -68485 -40890 -68165 -40828
rect -67485 -40272 -67165 -40210
rect -67485 -40508 -67443 -40272
rect -67207 -40508 -67165 -40272
rect -67485 -40592 -67165 -40508
rect -67485 -40828 -67443 -40592
rect -67207 -40828 -67165 -40592
rect -67485 -40890 -67165 -40828
rect -66485 -40272 -66165 -40210
rect -66485 -40508 -66443 -40272
rect -66207 -40508 -66165 -40272
rect -66485 -40592 -66165 -40508
rect -66485 -40828 -66443 -40592
rect -66207 -40828 -66165 -40592
rect -66485 -40890 -66165 -40828
rect -65485 -40272 -65165 -40210
rect -65485 -40508 -65443 -40272
rect -65207 -40508 -65165 -40272
rect -65485 -40592 -65165 -40508
rect -65485 -40828 -65443 -40592
rect -65207 -40828 -65165 -40592
rect -65485 -40890 -65165 -40828
rect -64485 -40272 -64165 -40210
rect -64485 -40508 -64443 -40272
rect -64207 -40508 -64165 -40272
rect -64485 -40592 -64165 -40508
rect -64485 -40828 -64443 -40592
rect -64207 -40828 -64165 -40592
rect -64485 -40890 -64165 -40828
rect -63485 -40272 -63165 -40210
rect -63485 -40508 -63443 -40272
rect -63207 -40508 -63165 -40272
rect -63485 -40592 -63165 -40508
rect -63485 -40828 -63443 -40592
rect -63207 -40828 -63165 -40592
rect -63485 -40890 -63165 -40828
rect -62485 -40272 -62165 -40210
rect -62485 -40508 -62443 -40272
rect -62207 -40508 -62165 -40272
rect -62485 -40592 -62165 -40508
rect -62485 -40828 -62443 -40592
rect -62207 -40828 -62165 -40592
rect -62485 -40890 -62165 -40828
rect -61485 -40272 -61165 -40210
rect -61485 -40508 -61443 -40272
rect -61207 -40508 -61165 -40272
rect -61485 -40592 -61165 -40508
rect -61485 -40828 -61443 -40592
rect -61207 -40828 -61165 -40592
rect -61485 -40890 -61165 -40828
rect -60485 -40272 -60165 -40210
rect -60485 -40508 -60443 -40272
rect -60207 -40508 -60165 -40272
rect -60485 -40592 -60165 -40508
rect -60485 -40828 -60443 -40592
rect -60207 -40828 -60165 -40592
rect -60485 -40890 -60165 -40828
rect -59485 -40272 -59165 -40210
rect -59485 -40508 -59443 -40272
rect -59207 -40508 -59165 -40272
rect -59485 -40592 -59165 -40508
rect -59485 -40828 -59443 -40592
rect -59207 -40828 -59165 -40592
rect -59485 -40890 -59165 -40828
rect -58485 -40272 -58165 -40210
rect -58485 -40508 -58443 -40272
rect -58207 -40508 -58165 -40272
rect -58485 -40592 -58165 -40508
rect -58485 -40828 -58443 -40592
rect -58207 -40828 -58165 -40592
rect -58485 -40890 -58165 -40828
rect -57485 -40272 -57165 -40210
rect -57485 -40508 -57443 -40272
rect -57207 -40508 -57165 -40272
rect -57485 -40592 -57165 -40508
rect -57485 -40828 -57443 -40592
rect -57207 -40828 -57165 -40592
rect -57485 -40890 -57165 -40828
rect -56485 -40272 -56165 -40210
rect -56485 -40508 -56443 -40272
rect -56207 -40508 -56165 -40272
rect -56485 -40592 -56165 -40508
rect -56485 -40828 -56443 -40592
rect -56207 -40828 -56165 -40592
rect -56485 -40890 -56165 -40828
rect -55485 -40272 -55165 -40210
rect -55485 -40508 -55443 -40272
rect -55207 -40508 -55165 -40272
rect -55485 -40592 -55165 -40508
rect -55485 -40828 -55443 -40592
rect -55207 -40828 -55165 -40592
rect -55485 -40890 -55165 -40828
rect -54485 -40272 -54165 -40210
rect -54485 -40508 -54443 -40272
rect -54207 -40508 -54165 -40272
rect -54485 -40592 -54165 -40508
rect -54485 -40828 -54443 -40592
rect -54207 -40828 -54165 -40592
rect -54485 -40890 -54165 -40828
rect -53485 -40272 -53165 -40210
rect -53485 -40508 -53443 -40272
rect -53207 -40508 -53165 -40272
rect -53485 -40592 -53165 -40508
rect -53485 -40828 -53443 -40592
rect -53207 -40828 -53165 -40592
rect -53485 -40890 -53165 -40828
rect -52485 -40272 -52165 -40210
rect -52485 -40508 -52443 -40272
rect -52207 -40508 -52165 -40272
rect -52485 -40592 -52165 -40508
rect -52485 -40828 -52443 -40592
rect -52207 -40828 -52165 -40592
rect -52485 -40890 -52165 -40828
rect -51485 -40272 -51165 -40210
rect -51485 -40508 -51443 -40272
rect -51207 -40508 -51165 -40272
rect -51485 -40592 -51165 -40508
rect -51485 -40828 -51443 -40592
rect -51207 -40828 -51165 -40592
rect -51485 -40890 -51165 -40828
rect -50485 -40272 -50165 -40210
rect -50485 -40508 -50443 -40272
rect -50207 -40508 -50165 -40272
rect -50485 -40592 -50165 -40508
rect -50485 -40828 -50443 -40592
rect -50207 -40828 -50165 -40592
rect -50485 -40890 -50165 -40828
rect -49485 -40272 -49165 -40210
rect -49485 -40508 -49443 -40272
rect -49207 -40508 -49165 -40272
rect -49485 -40592 -49165 -40508
rect -49485 -40828 -49443 -40592
rect -49207 -40828 -49165 -40592
rect -49485 -40890 -49165 -40828
rect -74825 -40932 -48825 -40890
rect -74825 -41168 -74783 -40932
rect -74547 -41168 -74443 -40932
rect -74207 -41168 -74103 -40932
rect -73867 -41168 -73783 -40932
rect -73547 -41168 -73443 -40932
rect -73207 -41168 -73103 -40932
rect -72867 -41168 -72783 -40932
rect -72547 -41168 -72443 -40932
rect -72207 -41168 -72103 -40932
rect -71867 -41168 -71783 -40932
rect -71547 -41168 -71443 -40932
rect -71207 -41168 -71103 -40932
rect -70867 -41168 -70783 -40932
rect -70547 -41168 -70443 -40932
rect -70207 -41168 -70103 -40932
rect -69867 -41168 -69783 -40932
rect -69547 -41168 -69443 -40932
rect -69207 -41168 -69103 -40932
rect -68867 -41168 -68783 -40932
rect -68547 -41168 -68443 -40932
rect -68207 -41168 -68103 -40932
rect -67867 -41168 -67783 -40932
rect -67547 -41168 -67443 -40932
rect -67207 -41168 -67103 -40932
rect -66867 -41168 -66783 -40932
rect -66547 -41168 -66443 -40932
rect -66207 -41168 -66103 -40932
rect -65867 -41168 -65783 -40932
rect -65547 -41168 -65443 -40932
rect -65207 -41168 -65103 -40932
rect -64867 -41168 -64783 -40932
rect -64547 -41168 -64443 -40932
rect -64207 -41168 -64103 -40932
rect -63867 -41168 -63783 -40932
rect -63547 -41168 -63443 -40932
rect -63207 -41168 -63103 -40932
rect -62867 -41168 -62783 -40932
rect -62547 -41168 -62443 -40932
rect -62207 -41168 -62103 -40932
rect -61867 -41168 -61783 -40932
rect -61547 -41168 -61443 -40932
rect -61207 -41168 -61103 -40932
rect -60867 -41168 -60783 -40932
rect -60547 -41168 -60443 -40932
rect -60207 -41168 -60103 -40932
rect -59867 -41168 -59783 -40932
rect -59547 -41168 -59443 -40932
rect -59207 -41168 -59103 -40932
rect -58867 -41168 -58783 -40932
rect -58547 -41168 -58443 -40932
rect -58207 -41168 -58103 -40932
rect -57867 -41168 -57783 -40932
rect -57547 -41168 -57443 -40932
rect -57207 -41168 -57103 -40932
rect -56867 -41168 -56783 -40932
rect -56547 -41168 -56443 -40932
rect -56207 -41168 -56103 -40932
rect -55867 -41168 -55783 -40932
rect -55547 -41168 -55443 -40932
rect -55207 -41168 -55103 -40932
rect -54867 -41168 -54783 -40932
rect -54547 -41168 -54443 -40932
rect -54207 -41168 -54103 -40932
rect -53867 -41168 -53783 -40932
rect -53547 -41168 -53443 -40932
rect -53207 -41168 -53103 -40932
rect -52867 -41168 -52783 -40932
rect -52547 -41168 -52443 -40932
rect -52207 -41168 -52103 -40932
rect -51867 -41168 -51783 -40932
rect -51547 -41168 -51443 -40932
rect -51207 -41168 -51103 -40932
rect -50867 -41168 -50783 -40932
rect -50547 -41168 -50443 -40932
rect -50207 -41168 -50103 -40932
rect -49867 -41168 -49783 -40932
rect -49547 -41168 -49443 -40932
rect -49207 -41168 -49103 -40932
rect -48867 -41168 -48825 -40932
rect -74825 -41210 -48825 -41168
rect -74485 -41272 -74165 -41210
rect -74485 -41508 -74443 -41272
rect -74207 -41508 -74165 -41272
rect -74485 -41592 -74165 -41508
rect -74485 -41828 -74443 -41592
rect -74207 -41828 -74165 -41592
rect -74485 -41890 -74165 -41828
rect -73485 -41272 -73165 -41210
rect -73485 -41508 -73443 -41272
rect -73207 -41508 -73165 -41272
rect -73485 -41592 -73165 -41508
rect -73485 -41828 -73443 -41592
rect -73207 -41828 -73165 -41592
rect -73485 -41890 -73165 -41828
rect -72485 -41272 -72165 -41210
rect -72485 -41508 -72443 -41272
rect -72207 -41508 -72165 -41272
rect -72485 -41592 -72165 -41508
rect -72485 -41828 -72443 -41592
rect -72207 -41828 -72165 -41592
rect -72485 -41890 -72165 -41828
rect -71485 -41272 -71165 -41210
rect -71485 -41508 -71443 -41272
rect -71207 -41508 -71165 -41272
rect -71485 -41592 -71165 -41508
rect -71485 -41828 -71443 -41592
rect -71207 -41828 -71165 -41592
rect -71485 -41890 -71165 -41828
rect -70485 -41272 -70165 -41210
rect -70485 -41508 -70443 -41272
rect -70207 -41508 -70165 -41272
rect -70485 -41592 -70165 -41508
rect -70485 -41828 -70443 -41592
rect -70207 -41828 -70165 -41592
rect -70485 -41890 -70165 -41828
rect -69485 -41272 -69165 -41210
rect -69485 -41508 -69443 -41272
rect -69207 -41508 -69165 -41272
rect -69485 -41592 -69165 -41508
rect -69485 -41828 -69443 -41592
rect -69207 -41828 -69165 -41592
rect -69485 -41890 -69165 -41828
rect -68485 -41272 -68165 -41210
rect -68485 -41508 -68443 -41272
rect -68207 -41508 -68165 -41272
rect -68485 -41592 -68165 -41508
rect -68485 -41828 -68443 -41592
rect -68207 -41828 -68165 -41592
rect -68485 -41890 -68165 -41828
rect -67485 -41272 -67165 -41210
rect -67485 -41508 -67443 -41272
rect -67207 -41508 -67165 -41272
rect -67485 -41592 -67165 -41508
rect -67485 -41828 -67443 -41592
rect -67207 -41828 -67165 -41592
rect -67485 -41890 -67165 -41828
rect -66485 -41272 -66165 -41210
rect -66485 -41508 -66443 -41272
rect -66207 -41508 -66165 -41272
rect -66485 -41592 -66165 -41508
rect -66485 -41828 -66443 -41592
rect -66207 -41828 -66165 -41592
rect -66485 -41890 -66165 -41828
rect -65485 -41272 -65165 -41210
rect -65485 -41508 -65443 -41272
rect -65207 -41508 -65165 -41272
rect -65485 -41592 -65165 -41508
rect -65485 -41828 -65443 -41592
rect -65207 -41828 -65165 -41592
rect -65485 -41890 -65165 -41828
rect -64485 -41272 -64165 -41210
rect -64485 -41508 -64443 -41272
rect -64207 -41508 -64165 -41272
rect -64485 -41592 -64165 -41508
rect -64485 -41828 -64443 -41592
rect -64207 -41828 -64165 -41592
rect -64485 -41890 -64165 -41828
rect -63485 -41272 -63165 -41210
rect -63485 -41508 -63443 -41272
rect -63207 -41508 -63165 -41272
rect -63485 -41592 -63165 -41508
rect -63485 -41828 -63443 -41592
rect -63207 -41828 -63165 -41592
rect -63485 -41890 -63165 -41828
rect -62485 -41272 -62165 -41210
rect -62485 -41508 -62443 -41272
rect -62207 -41508 -62165 -41272
rect -62485 -41592 -62165 -41508
rect -62485 -41828 -62443 -41592
rect -62207 -41828 -62165 -41592
rect -62485 -41890 -62165 -41828
rect -61485 -41272 -61165 -41210
rect -61485 -41508 -61443 -41272
rect -61207 -41508 -61165 -41272
rect -61485 -41592 -61165 -41508
rect -61485 -41828 -61443 -41592
rect -61207 -41828 -61165 -41592
rect -61485 -41890 -61165 -41828
rect -60485 -41272 -60165 -41210
rect -60485 -41508 -60443 -41272
rect -60207 -41508 -60165 -41272
rect -60485 -41592 -60165 -41508
rect -60485 -41828 -60443 -41592
rect -60207 -41828 -60165 -41592
rect -60485 -41890 -60165 -41828
rect -59485 -41272 -59165 -41210
rect -59485 -41508 -59443 -41272
rect -59207 -41508 -59165 -41272
rect -59485 -41592 -59165 -41508
rect -59485 -41828 -59443 -41592
rect -59207 -41828 -59165 -41592
rect -59485 -41890 -59165 -41828
rect -58485 -41272 -58165 -41210
rect -58485 -41508 -58443 -41272
rect -58207 -41508 -58165 -41272
rect -58485 -41592 -58165 -41508
rect -58485 -41828 -58443 -41592
rect -58207 -41828 -58165 -41592
rect -58485 -41890 -58165 -41828
rect -57485 -41272 -57165 -41210
rect -57485 -41508 -57443 -41272
rect -57207 -41508 -57165 -41272
rect -57485 -41592 -57165 -41508
rect -57485 -41828 -57443 -41592
rect -57207 -41828 -57165 -41592
rect -57485 -41890 -57165 -41828
rect -56485 -41272 -56165 -41210
rect -56485 -41508 -56443 -41272
rect -56207 -41508 -56165 -41272
rect -56485 -41592 -56165 -41508
rect -56485 -41828 -56443 -41592
rect -56207 -41828 -56165 -41592
rect -56485 -41890 -56165 -41828
rect -55485 -41272 -55165 -41210
rect -55485 -41508 -55443 -41272
rect -55207 -41508 -55165 -41272
rect -55485 -41592 -55165 -41508
rect -55485 -41828 -55443 -41592
rect -55207 -41828 -55165 -41592
rect -55485 -41890 -55165 -41828
rect -54485 -41272 -54165 -41210
rect -54485 -41508 -54443 -41272
rect -54207 -41508 -54165 -41272
rect -54485 -41592 -54165 -41508
rect -54485 -41828 -54443 -41592
rect -54207 -41828 -54165 -41592
rect -54485 -41890 -54165 -41828
rect -53485 -41272 -53165 -41210
rect -53485 -41508 -53443 -41272
rect -53207 -41508 -53165 -41272
rect -53485 -41592 -53165 -41508
rect -53485 -41828 -53443 -41592
rect -53207 -41828 -53165 -41592
rect -53485 -41890 -53165 -41828
rect -52485 -41272 -52165 -41210
rect -52485 -41508 -52443 -41272
rect -52207 -41508 -52165 -41272
rect -52485 -41592 -52165 -41508
rect -52485 -41828 -52443 -41592
rect -52207 -41828 -52165 -41592
rect -52485 -41890 -52165 -41828
rect -51485 -41272 -51165 -41210
rect -51485 -41508 -51443 -41272
rect -51207 -41508 -51165 -41272
rect -51485 -41592 -51165 -41508
rect -51485 -41828 -51443 -41592
rect -51207 -41828 -51165 -41592
rect -51485 -41890 -51165 -41828
rect -50485 -41272 -50165 -41210
rect -50485 -41508 -50443 -41272
rect -50207 -41508 -50165 -41272
rect -50485 -41592 -50165 -41508
rect -50485 -41828 -50443 -41592
rect -50207 -41828 -50165 -41592
rect -50485 -41890 -50165 -41828
rect -49485 -41272 -49165 -41210
rect -49485 -41508 -49443 -41272
rect -49207 -41508 -49165 -41272
rect -49485 -41592 -49165 -41508
rect -49485 -41828 -49443 -41592
rect -49207 -41828 -49165 -41592
rect -49485 -41890 -49165 -41828
rect -74825 -41932 -48825 -41890
rect -74825 -42168 -74783 -41932
rect -74547 -42168 -74443 -41932
rect -74207 -42168 -74103 -41932
rect -73867 -42168 -73783 -41932
rect -73547 -42168 -73443 -41932
rect -73207 -42168 -73103 -41932
rect -72867 -42168 -72783 -41932
rect -72547 -42168 -72443 -41932
rect -72207 -42168 -72103 -41932
rect -71867 -42168 -71783 -41932
rect -71547 -42168 -71443 -41932
rect -71207 -42168 -71103 -41932
rect -70867 -42168 -70783 -41932
rect -70547 -42168 -70443 -41932
rect -70207 -42168 -70103 -41932
rect -69867 -42168 -69783 -41932
rect -69547 -42168 -69443 -41932
rect -69207 -42168 -69103 -41932
rect -68867 -42168 -68783 -41932
rect -68547 -42168 -68443 -41932
rect -68207 -42168 -68103 -41932
rect -67867 -42168 -67783 -41932
rect -67547 -42168 -67443 -41932
rect -67207 -42168 -67103 -41932
rect -66867 -42168 -66783 -41932
rect -66547 -42168 -66443 -41932
rect -66207 -42168 -66103 -41932
rect -65867 -42168 -65783 -41932
rect -65547 -42168 -65443 -41932
rect -65207 -42168 -65103 -41932
rect -64867 -42168 -64783 -41932
rect -64547 -42168 -64443 -41932
rect -64207 -42168 -64103 -41932
rect -63867 -42168 -63783 -41932
rect -63547 -42168 -63443 -41932
rect -63207 -42168 -63103 -41932
rect -62867 -42168 -62783 -41932
rect -62547 -42168 -62443 -41932
rect -62207 -42168 -62103 -41932
rect -61867 -42168 -61783 -41932
rect -61547 -42168 -61443 -41932
rect -61207 -42168 -61103 -41932
rect -60867 -42168 -60783 -41932
rect -60547 -42168 -60443 -41932
rect -60207 -42168 -60103 -41932
rect -59867 -42168 -59783 -41932
rect -59547 -42168 -59443 -41932
rect -59207 -42168 -59103 -41932
rect -58867 -42168 -58783 -41932
rect -58547 -42168 -58443 -41932
rect -58207 -42168 -58103 -41932
rect -57867 -42168 -57783 -41932
rect -57547 -42168 -57443 -41932
rect -57207 -42168 -57103 -41932
rect -56867 -42168 -56783 -41932
rect -56547 -42168 -56443 -41932
rect -56207 -42168 -56103 -41932
rect -55867 -42168 -55783 -41932
rect -55547 -42168 -55443 -41932
rect -55207 -42168 -55103 -41932
rect -54867 -42168 -54783 -41932
rect -54547 -42168 -54443 -41932
rect -54207 -42168 -54103 -41932
rect -53867 -42168 -53783 -41932
rect -53547 -42168 -53443 -41932
rect -53207 -42168 -53103 -41932
rect -52867 -42168 -52783 -41932
rect -52547 -42168 -52443 -41932
rect -52207 -42168 -52103 -41932
rect -51867 -42168 -51783 -41932
rect -51547 -42168 -51443 -41932
rect -51207 -42168 -51103 -41932
rect -50867 -42168 -50783 -41932
rect -50547 -42168 -50443 -41932
rect -50207 -42168 -50103 -41932
rect -49867 -42168 -49783 -41932
rect -49547 -42168 -49443 -41932
rect -49207 -42168 -49103 -41932
rect -48867 -42168 -48825 -41932
rect -74825 -42210 -48825 -42168
rect -74485 -42272 -74165 -42210
rect -74485 -42508 -74443 -42272
rect -74207 -42508 -74165 -42272
rect -74485 -42592 -74165 -42508
rect -74485 -42828 -74443 -42592
rect -74207 -42828 -74165 -42592
rect -74485 -42890 -74165 -42828
rect -73485 -42272 -73165 -42210
rect -73485 -42508 -73443 -42272
rect -73207 -42508 -73165 -42272
rect -73485 -42592 -73165 -42508
rect -73485 -42828 -73443 -42592
rect -73207 -42828 -73165 -42592
rect -73485 -42890 -73165 -42828
rect -72485 -42272 -72165 -42210
rect -72485 -42508 -72443 -42272
rect -72207 -42508 -72165 -42272
rect -72485 -42592 -72165 -42508
rect -72485 -42828 -72443 -42592
rect -72207 -42828 -72165 -42592
rect -72485 -42890 -72165 -42828
rect -71485 -42272 -71165 -42210
rect -71485 -42508 -71443 -42272
rect -71207 -42508 -71165 -42272
rect -71485 -42592 -71165 -42508
rect -71485 -42828 -71443 -42592
rect -71207 -42828 -71165 -42592
rect -71485 -42890 -71165 -42828
rect -70485 -42272 -70165 -42210
rect -70485 -42508 -70443 -42272
rect -70207 -42508 -70165 -42272
rect -70485 -42592 -70165 -42508
rect -70485 -42828 -70443 -42592
rect -70207 -42828 -70165 -42592
rect -70485 -42890 -70165 -42828
rect -69485 -42272 -69165 -42210
rect -69485 -42508 -69443 -42272
rect -69207 -42508 -69165 -42272
rect -69485 -42592 -69165 -42508
rect -69485 -42828 -69443 -42592
rect -69207 -42828 -69165 -42592
rect -69485 -42890 -69165 -42828
rect -68485 -42272 -68165 -42210
rect -68485 -42508 -68443 -42272
rect -68207 -42508 -68165 -42272
rect -68485 -42592 -68165 -42508
rect -68485 -42828 -68443 -42592
rect -68207 -42828 -68165 -42592
rect -68485 -42890 -68165 -42828
rect -67485 -42272 -67165 -42210
rect -67485 -42508 -67443 -42272
rect -67207 -42508 -67165 -42272
rect -67485 -42592 -67165 -42508
rect -67485 -42828 -67443 -42592
rect -67207 -42828 -67165 -42592
rect -67485 -42890 -67165 -42828
rect -66485 -42272 -66165 -42210
rect -66485 -42508 -66443 -42272
rect -66207 -42508 -66165 -42272
rect -66485 -42592 -66165 -42508
rect -66485 -42828 -66443 -42592
rect -66207 -42828 -66165 -42592
rect -66485 -42890 -66165 -42828
rect -65485 -42272 -65165 -42210
rect -65485 -42508 -65443 -42272
rect -65207 -42508 -65165 -42272
rect -65485 -42592 -65165 -42508
rect -65485 -42828 -65443 -42592
rect -65207 -42828 -65165 -42592
rect -65485 -42890 -65165 -42828
rect -64485 -42272 -64165 -42210
rect -64485 -42508 -64443 -42272
rect -64207 -42508 -64165 -42272
rect -64485 -42592 -64165 -42508
rect -64485 -42828 -64443 -42592
rect -64207 -42828 -64165 -42592
rect -64485 -42890 -64165 -42828
rect -63485 -42272 -63165 -42210
rect -63485 -42508 -63443 -42272
rect -63207 -42508 -63165 -42272
rect -63485 -42592 -63165 -42508
rect -63485 -42828 -63443 -42592
rect -63207 -42828 -63165 -42592
rect -63485 -42890 -63165 -42828
rect -62485 -42272 -62165 -42210
rect -62485 -42508 -62443 -42272
rect -62207 -42508 -62165 -42272
rect -62485 -42592 -62165 -42508
rect -62485 -42828 -62443 -42592
rect -62207 -42828 -62165 -42592
rect -62485 -42890 -62165 -42828
rect -61485 -42272 -61165 -42210
rect -61485 -42508 -61443 -42272
rect -61207 -42508 -61165 -42272
rect -61485 -42592 -61165 -42508
rect -61485 -42828 -61443 -42592
rect -61207 -42828 -61165 -42592
rect -61485 -42890 -61165 -42828
rect -60485 -42272 -60165 -42210
rect -60485 -42508 -60443 -42272
rect -60207 -42508 -60165 -42272
rect -60485 -42592 -60165 -42508
rect -60485 -42828 -60443 -42592
rect -60207 -42828 -60165 -42592
rect -60485 -42890 -60165 -42828
rect -59485 -42272 -59165 -42210
rect -59485 -42508 -59443 -42272
rect -59207 -42508 -59165 -42272
rect -59485 -42592 -59165 -42508
rect -59485 -42828 -59443 -42592
rect -59207 -42828 -59165 -42592
rect -59485 -42890 -59165 -42828
rect -58485 -42272 -58165 -42210
rect -58485 -42508 -58443 -42272
rect -58207 -42508 -58165 -42272
rect -58485 -42592 -58165 -42508
rect -58485 -42828 -58443 -42592
rect -58207 -42828 -58165 -42592
rect -58485 -42890 -58165 -42828
rect -57485 -42272 -57165 -42210
rect -57485 -42508 -57443 -42272
rect -57207 -42508 -57165 -42272
rect -57485 -42592 -57165 -42508
rect -57485 -42828 -57443 -42592
rect -57207 -42828 -57165 -42592
rect -57485 -42890 -57165 -42828
rect -56485 -42272 -56165 -42210
rect -56485 -42508 -56443 -42272
rect -56207 -42508 -56165 -42272
rect -56485 -42592 -56165 -42508
rect -56485 -42828 -56443 -42592
rect -56207 -42828 -56165 -42592
rect -56485 -42890 -56165 -42828
rect -55485 -42272 -55165 -42210
rect -55485 -42508 -55443 -42272
rect -55207 -42508 -55165 -42272
rect -55485 -42592 -55165 -42508
rect -55485 -42828 -55443 -42592
rect -55207 -42828 -55165 -42592
rect -55485 -42890 -55165 -42828
rect -54485 -42272 -54165 -42210
rect -54485 -42508 -54443 -42272
rect -54207 -42508 -54165 -42272
rect -54485 -42592 -54165 -42508
rect -54485 -42828 -54443 -42592
rect -54207 -42828 -54165 -42592
rect -54485 -42890 -54165 -42828
rect -53485 -42272 -53165 -42210
rect -53485 -42508 -53443 -42272
rect -53207 -42508 -53165 -42272
rect -53485 -42592 -53165 -42508
rect -53485 -42828 -53443 -42592
rect -53207 -42828 -53165 -42592
rect -53485 -42890 -53165 -42828
rect -52485 -42272 -52165 -42210
rect -52485 -42508 -52443 -42272
rect -52207 -42508 -52165 -42272
rect -52485 -42592 -52165 -42508
rect -52485 -42828 -52443 -42592
rect -52207 -42828 -52165 -42592
rect -52485 -42890 -52165 -42828
rect -51485 -42272 -51165 -42210
rect -51485 -42508 -51443 -42272
rect -51207 -42508 -51165 -42272
rect -51485 -42592 -51165 -42508
rect -51485 -42828 -51443 -42592
rect -51207 -42828 -51165 -42592
rect -51485 -42890 -51165 -42828
rect -50485 -42272 -50165 -42210
rect -50485 -42508 -50443 -42272
rect -50207 -42508 -50165 -42272
rect -50485 -42592 -50165 -42508
rect -50485 -42828 -50443 -42592
rect -50207 -42828 -50165 -42592
rect -50485 -42890 -50165 -42828
rect -49485 -42272 -49165 -42210
rect -49485 -42508 -49443 -42272
rect -49207 -42508 -49165 -42272
rect -49485 -42592 -49165 -42508
rect -49485 -42828 -49443 -42592
rect -49207 -42828 -49165 -42592
rect -49485 -42890 -49165 -42828
rect -74825 -42932 -48825 -42890
rect -74825 -43168 -74783 -42932
rect -74547 -43168 -74443 -42932
rect -74207 -43168 -74103 -42932
rect -73867 -43168 -73783 -42932
rect -73547 -43168 -73443 -42932
rect -73207 -43168 -73103 -42932
rect -72867 -43168 -72783 -42932
rect -72547 -43168 -72443 -42932
rect -72207 -43168 -72103 -42932
rect -71867 -43168 -71783 -42932
rect -71547 -43168 -71443 -42932
rect -71207 -43168 -71103 -42932
rect -70867 -43168 -70783 -42932
rect -70547 -43168 -70443 -42932
rect -70207 -43168 -70103 -42932
rect -69867 -43168 -69783 -42932
rect -69547 -43168 -69443 -42932
rect -69207 -43168 -69103 -42932
rect -68867 -43168 -68783 -42932
rect -68547 -43168 -68443 -42932
rect -68207 -43168 -68103 -42932
rect -67867 -43168 -67783 -42932
rect -67547 -43168 -67443 -42932
rect -67207 -43168 -67103 -42932
rect -66867 -43168 -66783 -42932
rect -66547 -43168 -66443 -42932
rect -66207 -43168 -66103 -42932
rect -65867 -43168 -65783 -42932
rect -65547 -43168 -65443 -42932
rect -65207 -43168 -65103 -42932
rect -64867 -43168 -64783 -42932
rect -64547 -43168 -64443 -42932
rect -64207 -43168 -64103 -42932
rect -63867 -43168 -63783 -42932
rect -63547 -43168 -63443 -42932
rect -63207 -43168 -63103 -42932
rect -62867 -43168 -62783 -42932
rect -62547 -43168 -62443 -42932
rect -62207 -43168 -62103 -42932
rect -61867 -43168 -61783 -42932
rect -61547 -43168 -61443 -42932
rect -61207 -43168 -61103 -42932
rect -60867 -43168 -60783 -42932
rect -60547 -43168 -60443 -42932
rect -60207 -43168 -60103 -42932
rect -59867 -43168 -59783 -42932
rect -59547 -43168 -59443 -42932
rect -59207 -43168 -59103 -42932
rect -58867 -43168 -58783 -42932
rect -58547 -43168 -58443 -42932
rect -58207 -43168 -58103 -42932
rect -57867 -43168 -57783 -42932
rect -57547 -43168 -57443 -42932
rect -57207 -43168 -57103 -42932
rect -56867 -43168 -56783 -42932
rect -56547 -43168 -56443 -42932
rect -56207 -43168 -56103 -42932
rect -55867 -43168 -55783 -42932
rect -55547 -43168 -55443 -42932
rect -55207 -43168 -55103 -42932
rect -54867 -43168 -54783 -42932
rect -54547 -43168 -54443 -42932
rect -54207 -43168 -54103 -42932
rect -53867 -43168 -53783 -42932
rect -53547 -43168 -53443 -42932
rect -53207 -43168 -53103 -42932
rect -52867 -43168 -52783 -42932
rect -52547 -43168 -52443 -42932
rect -52207 -43168 -52103 -42932
rect -51867 -43168 -51783 -42932
rect -51547 -43168 -51443 -42932
rect -51207 -43168 -51103 -42932
rect -50867 -43168 -50783 -42932
rect -50547 -43168 -50443 -42932
rect -50207 -43168 -50103 -42932
rect -49867 -43168 -49783 -42932
rect -49547 -43168 -49443 -42932
rect -49207 -43168 -49103 -42932
rect -48867 -43168 -48825 -42932
rect -74825 -43210 -48825 -43168
rect -74485 -43272 -74165 -43210
rect -74485 -43508 -74443 -43272
rect -74207 -43508 -74165 -43272
rect -74485 -43592 -74165 -43508
rect -74485 -43828 -74443 -43592
rect -74207 -43828 -74165 -43592
rect -74485 -43890 -74165 -43828
rect -73485 -43272 -73165 -43210
rect -73485 -43508 -73443 -43272
rect -73207 -43508 -73165 -43272
rect -73485 -43592 -73165 -43508
rect -73485 -43828 -73443 -43592
rect -73207 -43828 -73165 -43592
rect -73485 -43890 -73165 -43828
rect -72485 -43272 -72165 -43210
rect -72485 -43508 -72443 -43272
rect -72207 -43508 -72165 -43272
rect -72485 -43592 -72165 -43508
rect -72485 -43828 -72443 -43592
rect -72207 -43828 -72165 -43592
rect -72485 -43890 -72165 -43828
rect -71485 -43272 -71165 -43210
rect -71485 -43508 -71443 -43272
rect -71207 -43508 -71165 -43272
rect -71485 -43592 -71165 -43508
rect -71485 -43828 -71443 -43592
rect -71207 -43828 -71165 -43592
rect -71485 -43890 -71165 -43828
rect -70485 -43272 -70165 -43210
rect -70485 -43508 -70443 -43272
rect -70207 -43508 -70165 -43272
rect -70485 -43592 -70165 -43508
rect -70485 -43828 -70443 -43592
rect -70207 -43828 -70165 -43592
rect -70485 -43890 -70165 -43828
rect -69485 -43272 -69165 -43210
rect -69485 -43508 -69443 -43272
rect -69207 -43508 -69165 -43272
rect -69485 -43592 -69165 -43508
rect -69485 -43828 -69443 -43592
rect -69207 -43828 -69165 -43592
rect -69485 -43890 -69165 -43828
rect -68485 -43272 -68165 -43210
rect -68485 -43508 -68443 -43272
rect -68207 -43508 -68165 -43272
rect -68485 -43592 -68165 -43508
rect -68485 -43828 -68443 -43592
rect -68207 -43828 -68165 -43592
rect -68485 -43890 -68165 -43828
rect -67485 -43272 -67165 -43210
rect -67485 -43508 -67443 -43272
rect -67207 -43508 -67165 -43272
rect -67485 -43592 -67165 -43508
rect -67485 -43828 -67443 -43592
rect -67207 -43828 -67165 -43592
rect -67485 -43890 -67165 -43828
rect -66485 -43272 -66165 -43210
rect -66485 -43508 -66443 -43272
rect -66207 -43508 -66165 -43272
rect -66485 -43592 -66165 -43508
rect -66485 -43828 -66443 -43592
rect -66207 -43828 -66165 -43592
rect -66485 -43890 -66165 -43828
rect -65485 -43272 -65165 -43210
rect -65485 -43508 -65443 -43272
rect -65207 -43508 -65165 -43272
rect -65485 -43592 -65165 -43508
rect -65485 -43828 -65443 -43592
rect -65207 -43828 -65165 -43592
rect -65485 -43890 -65165 -43828
rect -64485 -43272 -64165 -43210
rect -64485 -43508 -64443 -43272
rect -64207 -43508 -64165 -43272
rect -64485 -43592 -64165 -43508
rect -64485 -43828 -64443 -43592
rect -64207 -43828 -64165 -43592
rect -64485 -43890 -64165 -43828
rect -63485 -43272 -63165 -43210
rect -63485 -43508 -63443 -43272
rect -63207 -43508 -63165 -43272
rect -63485 -43592 -63165 -43508
rect -63485 -43828 -63443 -43592
rect -63207 -43828 -63165 -43592
rect -63485 -43890 -63165 -43828
rect -62485 -43272 -62165 -43210
rect -62485 -43508 -62443 -43272
rect -62207 -43508 -62165 -43272
rect -62485 -43592 -62165 -43508
rect -62485 -43828 -62443 -43592
rect -62207 -43828 -62165 -43592
rect -62485 -43890 -62165 -43828
rect -61485 -43272 -61165 -43210
rect -61485 -43508 -61443 -43272
rect -61207 -43508 -61165 -43272
rect -61485 -43592 -61165 -43508
rect -61485 -43828 -61443 -43592
rect -61207 -43828 -61165 -43592
rect -61485 -43890 -61165 -43828
rect -60485 -43272 -60165 -43210
rect -60485 -43508 -60443 -43272
rect -60207 -43508 -60165 -43272
rect -60485 -43592 -60165 -43508
rect -60485 -43828 -60443 -43592
rect -60207 -43828 -60165 -43592
rect -60485 -43890 -60165 -43828
rect -59485 -43272 -59165 -43210
rect -59485 -43508 -59443 -43272
rect -59207 -43508 -59165 -43272
rect -59485 -43592 -59165 -43508
rect -59485 -43828 -59443 -43592
rect -59207 -43828 -59165 -43592
rect -59485 -43890 -59165 -43828
rect -58485 -43272 -58165 -43210
rect -58485 -43508 -58443 -43272
rect -58207 -43508 -58165 -43272
rect -58485 -43592 -58165 -43508
rect -58485 -43828 -58443 -43592
rect -58207 -43828 -58165 -43592
rect -58485 -43890 -58165 -43828
rect -57485 -43272 -57165 -43210
rect -57485 -43508 -57443 -43272
rect -57207 -43508 -57165 -43272
rect -57485 -43592 -57165 -43508
rect -57485 -43828 -57443 -43592
rect -57207 -43828 -57165 -43592
rect -57485 -43890 -57165 -43828
rect -56485 -43272 -56165 -43210
rect -56485 -43508 -56443 -43272
rect -56207 -43508 -56165 -43272
rect -56485 -43592 -56165 -43508
rect -56485 -43828 -56443 -43592
rect -56207 -43828 -56165 -43592
rect -56485 -43890 -56165 -43828
rect -55485 -43272 -55165 -43210
rect -55485 -43508 -55443 -43272
rect -55207 -43508 -55165 -43272
rect -55485 -43592 -55165 -43508
rect -55485 -43828 -55443 -43592
rect -55207 -43828 -55165 -43592
rect -55485 -43890 -55165 -43828
rect -54485 -43272 -54165 -43210
rect -54485 -43508 -54443 -43272
rect -54207 -43508 -54165 -43272
rect -54485 -43592 -54165 -43508
rect -54485 -43828 -54443 -43592
rect -54207 -43828 -54165 -43592
rect -54485 -43890 -54165 -43828
rect -53485 -43272 -53165 -43210
rect -53485 -43508 -53443 -43272
rect -53207 -43508 -53165 -43272
rect -53485 -43592 -53165 -43508
rect -53485 -43828 -53443 -43592
rect -53207 -43828 -53165 -43592
rect -53485 -43890 -53165 -43828
rect -52485 -43272 -52165 -43210
rect -52485 -43508 -52443 -43272
rect -52207 -43508 -52165 -43272
rect -52485 -43592 -52165 -43508
rect -52485 -43828 -52443 -43592
rect -52207 -43828 -52165 -43592
rect -52485 -43890 -52165 -43828
rect -51485 -43272 -51165 -43210
rect -51485 -43508 -51443 -43272
rect -51207 -43508 -51165 -43272
rect -51485 -43592 -51165 -43508
rect -51485 -43828 -51443 -43592
rect -51207 -43828 -51165 -43592
rect -51485 -43890 -51165 -43828
rect -50485 -43272 -50165 -43210
rect -50485 -43508 -50443 -43272
rect -50207 -43508 -50165 -43272
rect -50485 -43592 -50165 -43508
rect -50485 -43828 -50443 -43592
rect -50207 -43828 -50165 -43592
rect -50485 -43890 -50165 -43828
rect -49485 -43272 -49165 -43210
rect -49485 -43508 -49443 -43272
rect -49207 -43508 -49165 -43272
rect -49485 -43592 -49165 -43508
rect -49485 -43828 -49443 -43592
rect -49207 -43828 -49165 -43592
rect -49485 -43890 -49165 -43828
rect -74825 -43932 -48825 -43890
rect -74825 -44168 -74783 -43932
rect -74547 -44168 -74443 -43932
rect -74207 -44168 -74103 -43932
rect -73867 -44168 -73783 -43932
rect -73547 -44168 -73443 -43932
rect -73207 -44168 -73103 -43932
rect -72867 -44168 -72783 -43932
rect -72547 -44168 -72443 -43932
rect -72207 -44168 -72103 -43932
rect -71867 -44168 -71783 -43932
rect -71547 -44168 -71443 -43932
rect -71207 -44168 -71103 -43932
rect -70867 -44168 -70783 -43932
rect -70547 -44168 -70443 -43932
rect -70207 -44168 -70103 -43932
rect -69867 -44168 -69783 -43932
rect -69547 -44168 -69443 -43932
rect -69207 -44168 -69103 -43932
rect -68867 -44168 -68783 -43932
rect -68547 -44168 -68443 -43932
rect -68207 -44168 -68103 -43932
rect -67867 -44168 -67783 -43932
rect -67547 -44168 -67443 -43932
rect -67207 -44168 -67103 -43932
rect -66867 -44168 -66783 -43932
rect -66547 -44168 -66443 -43932
rect -66207 -44168 -66103 -43932
rect -65867 -44168 -65783 -43932
rect -65547 -44168 -65443 -43932
rect -65207 -44168 -65103 -43932
rect -64867 -44168 -64783 -43932
rect -64547 -44168 -64443 -43932
rect -64207 -44168 -64103 -43932
rect -63867 -44168 -63783 -43932
rect -63547 -44168 -63443 -43932
rect -63207 -44168 -63103 -43932
rect -62867 -44168 -62783 -43932
rect -62547 -44168 -62443 -43932
rect -62207 -44168 -62103 -43932
rect -61867 -44168 -61783 -43932
rect -61547 -44168 -61443 -43932
rect -61207 -44168 -61103 -43932
rect -60867 -44168 -60783 -43932
rect -60547 -44168 -60443 -43932
rect -60207 -44168 -60103 -43932
rect -59867 -44168 -59783 -43932
rect -59547 -44168 -59443 -43932
rect -59207 -44168 -59103 -43932
rect -58867 -44168 -58783 -43932
rect -58547 -44168 -58443 -43932
rect -58207 -44168 -58103 -43932
rect -57867 -44168 -57783 -43932
rect -57547 -44168 -57443 -43932
rect -57207 -44168 -57103 -43932
rect -56867 -44168 -56783 -43932
rect -56547 -44168 -56443 -43932
rect -56207 -44168 -56103 -43932
rect -55867 -44168 -55783 -43932
rect -55547 -44168 -55443 -43932
rect -55207 -44168 -55103 -43932
rect -54867 -44168 -54783 -43932
rect -54547 -44168 -54443 -43932
rect -54207 -44168 -54103 -43932
rect -53867 -44168 -53783 -43932
rect -53547 -44168 -53443 -43932
rect -53207 -44168 -53103 -43932
rect -52867 -44168 -52783 -43932
rect -52547 -44168 -52443 -43932
rect -52207 -44168 -52103 -43932
rect -51867 -44168 -51783 -43932
rect -51547 -44168 -51443 -43932
rect -51207 -44168 -51103 -43932
rect -50867 -44168 -50783 -43932
rect -50547 -44168 -50443 -43932
rect -50207 -44168 -50103 -43932
rect -49867 -44168 -49783 -43932
rect -49547 -44168 -49443 -43932
rect -49207 -44168 -49103 -43932
rect -48867 -44168 -48825 -43932
rect -74825 -44210 -48825 -44168
rect -74485 -44272 -74165 -44210
rect -74485 -44508 -74443 -44272
rect -74207 -44508 -74165 -44272
rect -74485 -44592 -74165 -44508
rect -74485 -44828 -74443 -44592
rect -74207 -44828 -74165 -44592
rect -74485 -44890 -74165 -44828
rect -73485 -44272 -73165 -44210
rect -73485 -44508 -73443 -44272
rect -73207 -44508 -73165 -44272
rect -73485 -44592 -73165 -44508
rect -73485 -44828 -73443 -44592
rect -73207 -44828 -73165 -44592
rect -73485 -44890 -73165 -44828
rect -72485 -44272 -72165 -44210
rect -72485 -44508 -72443 -44272
rect -72207 -44508 -72165 -44272
rect -72485 -44592 -72165 -44508
rect -72485 -44828 -72443 -44592
rect -72207 -44828 -72165 -44592
rect -72485 -44890 -72165 -44828
rect -71485 -44272 -71165 -44210
rect -71485 -44508 -71443 -44272
rect -71207 -44508 -71165 -44272
rect -71485 -44592 -71165 -44508
rect -71485 -44828 -71443 -44592
rect -71207 -44828 -71165 -44592
rect -71485 -44890 -71165 -44828
rect -70485 -44272 -70165 -44210
rect -70485 -44508 -70443 -44272
rect -70207 -44508 -70165 -44272
rect -70485 -44592 -70165 -44508
rect -70485 -44828 -70443 -44592
rect -70207 -44828 -70165 -44592
rect -70485 -44890 -70165 -44828
rect -69485 -44272 -69165 -44210
rect -69485 -44508 -69443 -44272
rect -69207 -44508 -69165 -44272
rect -69485 -44592 -69165 -44508
rect -69485 -44828 -69443 -44592
rect -69207 -44828 -69165 -44592
rect -69485 -44890 -69165 -44828
rect -68485 -44272 -68165 -44210
rect -68485 -44508 -68443 -44272
rect -68207 -44508 -68165 -44272
rect -68485 -44592 -68165 -44508
rect -68485 -44828 -68443 -44592
rect -68207 -44828 -68165 -44592
rect -68485 -44890 -68165 -44828
rect -67485 -44272 -67165 -44210
rect -67485 -44508 -67443 -44272
rect -67207 -44508 -67165 -44272
rect -67485 -44592 -67165 -44508
rect -67485 -44828 -67443 -44592
rect -67207 -44828 -67165 -44592
rect -67485 -44890 -67165 -44828
rect -66485 -44272 -66165 -44210
rect -66485 -44508 -66443 -44272
rect -66207 -44508 -66165 -44272
rect -66485 -44592 -66165 -44508
rect -66485 -44828 -66443 -44592
rect -66207 -44828 -66165 -44592
rect -66485 -44890 -66165 -44828
rect -65485 -44272 -65165 -44210
rect -65485 -44508 -65443 -44272
rect -65207 -44508 -65165 -44272
rect -65485 -44592 -65165 -44508
rect -65485 -44828 -65443 -44592
rect -65207 -44828 -65165 -44592
rect -65485 -44890 -65165 -44828
rect -64485 -44272 -64165 -44210
rect -64485 -44508 -64443 -44272
rect -64207 -44508 -64165 -44272
rect -64485 -44592 -64165 -44508
rect -64485 -44828 -64443 -44592
rect -64207 -44828 -64165 -44592
rect -64485 -44890 -64165 -44828
rect -63485 -44272 -63165 -44210
rect -63485 -44508 -63443 -44272
rect -63207 -44508 -63165 -44272
rect -63485 -44592 -63165 -44508
rect -63485 -44828 -63443 -44592
rect -63207 -44828 -63165 -44592
rect -63485 -44890 -63165 -44828
rect -62485 -44272 -62165 -44210
rect -62485 -44508 -62443 -44272
rect -62207 -44508 -62165 -44272
rect -62485 -44592 -62165 -44508
rect -62485 -44828 -62443 -44592
rect -62207 -44828 -62165 -44592
rect -62485 -44890 -62165 -44828
rect -61485 -44272 -61165 -44210
rect -61485 -44508 -61443 -44272
rect -61207 -44508 -61165 -44272
rect -61485 -44592 -61165 -44508
rect -61485 -44828 -61443 -44592
rect -61207 -44828 -61165 -44592
rect -61485 -44890 -61165 -44828
rect -60485 -44272 -60165 -44210
rect -60485 -44508 -60443 -44272
rect -60207 -44508 -60165 -44272
rect -60485 -44592 -60165 -44508
rect -60485 -44828 -60443 -44592
rect -60207 -44828 -60165 -44592
rect -60485 -44890 -60165 -44828
rect -59485 -44272 -59165 -44210
rect -59485 -44508 -59443 -44272
rect -59207 -44508 -59165 -44272
rect -59485 -44592 -59165 -44508
rect -59485 -44828 -59443 -44592
rect -59207 -44828 -59165 -44592
rect -59485 -44890 -59165 -44828
rect -58485 -44272 -58165 -44210
rect -58485 -44508 -58443 -44272
rect -58207 -44508 -58165 -44272
rect -58485 -44592 -58165 -44508
rect -58485 -44828 -58443 -44592
rect -58207 -44828 -58165 -44592
rect -58485 -44890 -58165 -44828
rect -57485 -44272 -57165 -44210
rect -57485 -44508 -57443 -44272
rect -57207 -44508 -57165 -44272
rect -57485 -44592 -57165 -44508
rect -57485 -44828 -57443 -44592
rect -57207 -44828 -57165 -44592
rect -57485 -44890 -57165 -44828
rect -56485 -44272 -56165 -44210
rect -56485 -44508 -56443 -44272
rect -56207 -44508 -56165 -44272
rect -56485 -44592 -56165 -44508
rect -56485 -44828 -56443 -44592
rect -56207 -44828 -56165 -44592
rect -56485 -44890 -56165 -44828
rect -55485 -44272 -55165 -44210
rect -55485 -44508 -55443 -44272
rect -55207 -44508 -55165 -44272
rect -55485 -44592 -55165 -44508
rect -55485 -44828 -55443 -44592
rect -55207 -44828 -55165 -44592
rect -55485 -44890 -55165 -44828
rect -54485 -44272 -54165 -44210
rect -54485 -44508 -54443 -44272
rect -54207 -44508 -54165 -44272
rect -54485 -44592 -54165 -44508
rect -54485 -44828 -54443 -44592
rect -54207 -44828 -54165 -44592
rect -54485 -44890 -54165 -44828
rect -53485 -44272 -53165 -44210
rect -53485 -44508 -53443 -44272
rect -53207 -44508 -53165 -44272
rect -53485 -44592 -53165 -44508
rect -53485 -44828 -53443 -44592
rect -53207 -44828 -53165 -44592
rect -53485 -44890 -53165 -44828
rect -52485 -44272 -52165 -44210
rect -52485 -44508 -52443 -44272
rect -52207 -44508 -52165 -44272
rect -52485 -44592 -52165 -44508
rect -52485 -44828 -52443 -44592
rect -52207 -44828 -52165 -44592
rect -52485 -44890 -52165 -44828
rect -51485 -44272 -51165 -44210
rect -51485 -44508 -51443 -44272
rect -51207 -44508 -51165 -44272
rect -51485 -44592 -51165 -44508
rect -51485 -44828 -51443 -44592
rect -51207 -44828 -51165 -44592
rect -51485 -44890 -51165 -44828
rect -50485 -44272 -50165 -44210
rect -50485 -44508 -50443 -44272
rect -50207 -44508 -50165 -44272
rect -50485 -44592 -50165 -44508
rect -50485 -44828 -50443 -44592
rect -50207 -44828 -50165 -44592
rect -50485 -44890 -50165 -44828
rect -49485 -44272 -49165 -44210
rect -49485 -44508 -49443 -44272
rect -49207 -44508 -49165 -44272
rect -49485 -44592 -49165 -44508
rect -46275 -44428 -46198 -32672
rect -36362 -44428 -36275 -32672
tri -36275 -32700 -36155 -32580 nw
tri -23025 -32700 -22905 -32580 se
rect -22905 -32700 -17645 -32580
tri -17645 -32700 -17525 -32580 sw
tri -4395 -32700 -4275 -32580 ne
rect -4275 -32672 5725 -32580
tri -23215 -32890 -23025 -32700 se
rect -23025 -32890 -17525 -32700
tri -23535 -33210 -23215 -32890 se
rect -23215 -33210 -17525 -32890
tri -24215 -33890 -23535 -33210 se
rect -23535 -33890 -17525 -33210
tri -24535 -34210 -24215 -33890 se
rect -24215 -34210 -17525 -33890
tri -24875 -34550 -24535 -34210 se
rect -24535 -34550 -17525 -34210
tri -17525 -34550 -15675 -32700 sw
rect -24875 -42550 -15675 -34550
tri -24875 -42890 -24535 -42550 ne
rect -24535 -42890 -17645 -42550
tri -24535 -43210 -24215 -42890 ne
rect -24215 -43210 -17645 -42890
tri -24215 -43890 -23535 -43210 ne
rect -23535 -43890 -17645 -43210
tri -23535 -44210 -23215 -43890 ne
rect -23215 -44210 -17645 -43890
rect -46275 -44550 -36275 -44428
tri -23215 -44520 -22905 -44210 ne
rect -22905 -44520 -17645 -44210
tri -17645 -44520 -15675 -42550 nw
rect -4275 -44428 -4198 -32672
rect 5638 -44428 5725 -32672
rect 8615 -32592 8935 -32508
rect 8615 -32828 8657 -32592
rect 8893 -32828 8935 -32592
rect 8615 -32890 8935 -32828
rect 9615 -32272 9935 -32210
rect 9615 -32508 9657 -32272
rect 9893 -32508 9935 -32272
rect 9615 -32592 9935 -32508
rect 9615 -32828 9657 -32592
rect 9893 -32828 9935 -32592
rect 9615 -32890 9935 -32828
rect 10615 -32272 10935 -32210
rect 10615 -32508 10657 -32272
rect 10893 -32508 10935 -32272
rect 10615 -32592 10935 -32508
rect 10615 -32828 10657 -32592
rect 10893 -32828 10935 -32592
rect 10615 -32890 10935 -32828
rect 11615 -32272 11935 -32210
rect 11615 -32508 11657 -32272
rect 11893 -32508 11935 -32272
rect 11615 -32592 11935 -32508
rect 11615 -32828 11657 -32592
rect 11893 -32828 11935 -32592
rect 11615 -32890 11935 -32828
rect 12615 -32272 12935 -32210
rect 12615 -32508 12657 -32272
rect 12893 -32508 12935 -32272
rect 12615 -32592 12935 -32508
rect 12615 -32828 12657 -32592
rect 12893 -32828 12935 -32592
rect 12615 -32890 12935 -32828
rect 13615 -32272 13935 -32210
rect 13615 -32508 13657 -32272
rect 13893 -32508 13935 -32272
rect 13615 -32592 13935 -32508
rect 13615 -32828 13657 -32592
rect 13893 -32828 13935 -32592
rect 13615 -32890 13935 -32828
rect 14615 -32272 14935 -32210
rect 14615 -32508 14657 -32272
rect 14893 -32508 14935 -32272
rect 14615 -32592 14935 -32508
rect 14615 -32828 14657 -32592
rect 14893 -32828 14935 -32592
rect 14615 -32890 14935 -32828
rect 15615 -32272 15935 -32210
rect 15615 -32508 15657 -32272
rect 15893 -32508 15935 -32272
rect 15615 -32592 15935 -32508
rect 15615 -32828 15657 -32592
rect 15893 -32828 15935 -32592
rect 15615 -32890 15935 -32828
rect 16615 -32272 16935 -32210
rect 16615 -32508 16657 -32272
rect 16893 -32508 16935 -32272
rect 16615 -32592 16935 -32508
rect 16615 -32828 16657 -32592
rect 16893 -32828 16935 -32592
rect 16615 -32890 16935 -32828
rect 17615 -32272 17935 -32210
rect 17615 -32508 17657 -32272
rect 17893 -32508 17935 -32272
rect 17615 -32592 17935 -32508
rect 17615 -32828 17657 -32592
rect 17893 -32828 17935 -32592
rect 17615 -32890 17935 -32828
rect 18615 -32272 18935 -32210
rect 18615 -32508 18657 -32272
rect 18893 -32508 18935 -32272
rect 18615 -32592 18935 -32508
rect 18615 -32828 18657 -32592
rect 18893 -32828 18935 -32592
rect 18615 -32890 18935 -32828
rect 19615 -32272 19935 -32210
rect 19615 -32508 19657 -32272
rect 19893 -32508 19935 -32272
rect 19615 -32592 19935 -32508
rect 19615 -32828 19657 -32592
rect 19893 -32828 19935 -32592
rect 19615 -32890 19935 -32828
rect 20615 -32272 20935 -32210
rect 20615 -32508 20657 -32272
rect 20893 -32508 20935 -32272
rect 20615 -32592 20935 -32508
rect 20615 -32828 20657 -32592
rect 20893 -32828 20935 -32592
rect 20615 -32890 20935 -32828
rect 21615 -32272 21935 -32210
rect 21615 -32508 21657 -32272
rect 21893 -32508 21935 -32272
rect 21615 -32592 21935 -32508
rect 21615 -32828 21657 -32592
rect 21893 -32828 21935 -32592
rect 21615 -32890 21935 -32828
rect 22615 -32272 22935 -32210
rect 22615 -32508 22657 -32272
rect 22893 -32508 22935 -32272
rect 22615 -32592 22935 -32508
rect 22615 -32828 22657 -32592
rect 22893 -32828 22935 -32592
rect 22615 -32890 22935 -32828
rect 23615 -32272 23935 -32210
rect 23615 -32508 23657 -32272
rect 23893 -32508 23935 -32272
rect 23615 -32592 23935 -32508
rect 23615 -32828 23657 -32592
rect 23893 -32828 23935 -32592
rect 23615 -32890 23935 -32828
rect 24615 -32272 24935 -32210
rect 24615 -32508 24657 -32272
rect 24893 -32508 24935 -32272
rect 24615 -32592 24935 -32508
rect 24615 -32828 24657 -32592
rect 24893 -32828 24935 -32592
rect 24615 -32890 24935 -32828
rect 25615 -32272 25935 -32210
rect 25615 -32508 25657 -32272
rect 25893 -32508 25935 -32272
rect 25615 -32592 25935 -32508
rect 25615 -32828 25657 -32592
rect 25893 -32828 25935 -32592
rect 25615 -32890 25935 -32828
rect 26615 -32272 26935 -32210
rect 26615 -32508 26657 -32272
rect 26893 -32508 26935 -32272
rect 26615 -32592 26935 -32508
rect 26615 -32828 26657 -32592
rect 26893 -32828 26935 -32592
rect 26615 -32890 26935 -32828
rect 27615 -32272 27935 -32210
rect 27615 -32508 27657 -32272
rect 27893 -32508 27935 -32272
rect 27615 -32592 27935 -32508
rect 27615 -32828 27657 -32592
rect 27893 -32828 27935 -32592
rect 27615 -32890 27935 -32828
rect 28615 -32272 28935 -32210
rect 28615 -32508 28657 -32272
rect 28893 -32508 28935 -32272
rect 28615 -32592 28935 -32508
rect 28615 -32828 28657 -32592
rect 28893 -32828 28935 -32592
rect 28615 -32890 28935 -32828
rect 29615 -32272 29935 -32210
rect 29615 -32508 29657 -32272
rect 29893 -32508 29935 -32272
rect 29615 -32592 29935 -32508
rect 29615 -32828 29657 -32592
rect 29893 -32828 29935 -32592
rect 29615 -32890 29935 -32828
rect 30615 -32272 30935 -32210
rect 30615 -32508 30657 -32272
rect 30893 -32508 30935 -32272
rect 30615 -32592 30935 -32508
rect 30615 -32828 30657 -32592
rect 30893 -32828 30935 -32592
rect 30615 -32890 30935 -32828
rect 31615 -32272 31935 -32210
rect 31615 -32508 31657 -32272
rect 31893 -32508 31935 -32272
rect 31615 -32592 31935 -32508
rect 31615 -32828 31657 -32592
rect 31893 -32828 31935 -32592
rect 31615 -32890 31935 -32828
rect 32615 -32272 32935 -32210
rect 32615 -32508 32657 -32272
rect 32893 -32508 32935 -32272
rect 32615 -32592 32935 -32508
rect 32615 -32828 32657 -32592
rect 32893 -32828 32935 -32592
rect 32615 -32890 32935 -32828
rect 33615 -32272 33935 -32210
rect 33615 -32508 33657 -32272
rect 33893 -32508 33935 -32272
rect 33615 -32592 33935 -32508
rect 33615 -32828 33657 -32592
rect 33893 -32828 33935 -32592
rect 33615 -32890 33935 -32828
rect 8275 -32932 34275 -32890
rect 8275 -33168 8317 -32932
rect 8553 -33168 8657 -32932
rect 8893 -33168 8997 -32932
rect 9233 -33168 9317 -32932
rect 9553 -33168 9657 -32932
rect 9893 -33168 9997 -32932
rect 10233 -33168 10317 -32932
rect 10553 -33168 10657 -32932
rect 10893 -33168 10997 -32932
rect 11233 -33168 11317 -32932
rect 11553 -33168 11657 -32932
rect 11893 -33168 11997 -32932
rect 12233 -33168 12317 -32932
rect 12553 -33168 12657 -32932
rect 12893 -33168 12997 -32932
rect 13233 -33168 13317 -32932
rect 13553 -33168 13657 -32932
rect 13893 -33168 13997 -32932
rect 14233 -33168 14317 -32932
rect 14553 -33168 14657 -32932
rect 14893 -33168 14997 -32932
rect 15233 -33168 15317 -32932
rect 15553 -33168 15657 -32932
rect 15893 -33168 15997 -32932
rect 16233 -33168 16317 -32932
rect 16553 -33168 16657 -32932
rect 16893 -33168 16997 -32932
rect 17233 -33168 17317 -32932
rect 17553 -33168 17657 -32932
rect 17893 -33168 17997 -32932
rect 18233 -33168 18317 -32932
rect 18553 -33168 18657 -32932
rect 18893 -33168 18997 -32932
rect 19233 -33168 19317 -32932
rect 19553 -33168 19657 -32932
rect 19893 -33168 19997 -32932
rect 20233 -33168 20317 -32932
rect 20553 -33168 20657 -32932
rect 20893 -33168 20997 -32932
rect 21233 -33168 21317 -32932
rect 21553 -33168 21657 -32932
rect 21893 -33168 21997 -32932
rect 22233 -33168 22317 -32932
rect 22553 -33168 22657 -32932
rect 22893 -33168 22997 -32932
rect 23233 -33168 23317 -32932
rect 23553 -33168 23657 -32932
rect 23893 -33168 23997 -32932
rect 24233 -33168 24317 -32932
rect 24553 -33168 24657 -32932
rect 24893 -33168 24997 -32932
rect 25233 -33168 25317 -32932
rect 25553 -33168 25657 -32932
rect 25893 -33168 25997 -32932
rect 26233 -33168 26317 -32932
rect 26553 -33168 26657 -32932
rect 26893 -33168 26997 -32932
rect 27233 -33168 27317 -32932
rect 27553 -33168 27657 -32932
rect 27893 -33168 27997 -32932
rect 28233 -33168 28317 -32932
rect 28553 -33168 28657 -32932
rect 28893 -33168 28997 -32932
rect 29233 -33168 29317 -32932
rect 29553 -33168 29657 -32932
rect 29893 -33168 29997 -32932
rect 30233 -33168 30317 -32932
rect 30553 -33168 30657 -32932
rect 30893 -33168 30997 -32932
rect 31233 -33168 31317 -32932
rect 31553 -33168 31657 -32932
rect 31893 -33168 31997 -32932
rect 32233 -33168 32317 -32932
rect 32553 -33168 32657 -32932
rect 32893 -33168 32997 -32932
rect 33233 -33168 33317 -32932
rect 33553 -33168 33657 -32932
rect 33893 -33168 33997 -32932
rect 34233 -33168 34275 -32932
rect 8275 -33210 34275 -33168
rect 8615 -33272 8935 -33210
rect 8615 -33508 8657 -33272
rect 8893 -33508 8935 -33272
rect 8615 -33592 8935 -33508
rect 8615 -33828 8657 -33592
rect 8893 -33828 8935 -33592
rect 8615 -33890 8935 -33828
rect 9615 -33272 9935 -33210
rect 9615 -33508 9657 -33272
rect 9893 -33508 9935 -33272
rect 9615 -33592 9935 -33508
rect 9615 -33828 9657 -33592
rect 9893 -33828 9935 -33592
rect 9615 -33890 9935 -33828
rect 10615 -33272 10935 -33210
rect 10615 -33508 10657 -33272
rect 10893 -33508 10935 -33272
rect 10615 -33592 10935 -33508
rect 10615 -33828 10657 -33592
rect 10893 -33828 10935 -33592
rect 10615 -33890 10935 -33828
rect 11615 -33272 11935 -33210
rect 11615 -33508 11657 -33272
rect 11893 -33508 11935 -33272
rect 11615 -33592 11935 -33508
rect 11615 -33828 11657 -33592
rect 11893 -33828 11935 -33592
rect 11615 -33890 11935 -33828
rect 12615 -33272 12935 -33210
rect 12615 -33508 12657 -33272
rect 12893 -33508 12935 -33272
rect 12615 -33592 12935 -33508
rect 12615 -33828 12657 -33592
rect 12893 -33828 12935 -33592
rect 12615 -33890 12935 -33828
rect 13615 -33272 13935 -33210
rect 13615 -33508 13657 -33272
rect 13893 -33508 13935 -33272
rect 13615 -33592 13935 -33508
rect 13615 -33828 13657 -33592
rect 13893 -33828 13935 -33592
rect 13615 -33890 13935 -33828
rect 14615 -33272 14935 -33210
rect 14615 -33508 14657 -33272
rect 14893 -33508 14935 -33272
rect 14615 -33592 14935 -33508
rect 14615 -33828 14657 -33592
rect 14893 -33828 14935 -33592
rect 14615 -33890 14935 -33828
rect 15615 -33272 15935 -33210
rect 15615 -33508 15657 -33272
rect 15893 -33508 15935 -33272
rect 15615 -33592 15935 -33508
rect 15615 -33828 15657 -33592
rect 15893 -33828 15935 -33592
rect 15615 -33890 15935 -33828
rect 16615 -33272 16935 -33210
rect 16615 -33508 16657 -33272
rect 16893 -33508 16935 -33272
rect 16615 -33592 16935 -33508
rect 16615 -33828 16657 -33592
rect 16893 -33828 16935 -33592
rect 16615 -33890 16935 -33828
rect 17615 -33272 17935 -33210
rect 17615 -33508 17657 -33272
rect 17893 -33508 17935 -33272
rect 17615 -33592 17935 -33508
rect 17615 -33828 17657 -33592
rect 17893 -33828 17935 -33592
rect 17615 -33890 17935 -33828
rect 18615 -33272 18935 -33210
rect 18615 -33508 18657 -33272
rect 18893 -33508 18935 -33272
rect 18615 -33592 18935 -33508
rect 18615 -33828 18657 -33592
rect 18893 -33828 18935 -33592
rect 18615 -33890 18935 -33828
rect 19615 -33272 19935 -33210
rect 19615 -33508 19657 -33272
rect 19893 -33508 19935 -33272
rect 19615 -33592 19935 -33508
rect 19615 -33828 19657 -33592
rect 19893 -33828 19935 -33592
rect 19615 -33890 19935 -33828
rect 20615 -33272 20935 -33210
rect 20615 -33508 20657 -33272
rect 20893 -33508 20935 -33272
rect 20615 -33592 20935 -33508
rect 20615 -33828 20657 -33592
rect 20893 -33828 20935 -33592
rect 20615 -33890 20935 -33828
rect 21615 -33272 21935 -33210
rect 21615 -33508 21657 -33272
rect 21893 -33508 21935 -33272
rect 21615 -33592 21935 -33508
rect 21615 -33828 21657 -33592
rect 21893 -33828 21935 -33592
rect 21615 -33890 21935 -33828
rect 22615 -33272 22935 -33210
rect 22615 -33508 22657 -33272
rect 22893 -33508 22935 -33272
rect 22615 -33592 22935 -33508
rect 22615 -33828 22657 -33592
rect 22893 -33828 22935 -33592
rect 22615 -33890 22935 -33828
rect 23615 -33272 23935 -33210
rect 23615 -33508 23657 -33272
rect 23893 -33508 23935 -33272
rect 23615 -33592 23935 -33508
rect 23615 -33828 23657 -33592
rect 23893 -33828 23935 -33592
rect 23615 -33890 23935 -33828
rect 24615 -33272 24935 -33210
rect 24615 -33508 24657 -33272
rect 24893 -33508 24935 -33272
rect 24615 -33592 24935 -33508
rect 24615 -33828 24657 -33592
rect 24893 -33828 24935 -33592
rect 24615 -33890 24935 -33828
rect 25615 -33272 25935 -33210
rect 25615 -33508 25657 -33272
rect 25893 -33508 25935 -33272
rect 25615 -33592 25935 -33508
rect 25615 -33828 25657 -33592
rect 25893 -33828 25935 -33592
rect 25615 -33890 25935 -33828
rect 26615 -33272 26935 -33210
rect 26615 -33508 26657 -33272
rect 26893 -33508 26935 -33272
rect 26615 -33592 26935 -33508
rect 26615 -33828 26657 -33592
rect 26893 -33828 26935 -33592
rect 26615 -33890 26935 -33828
rect 27615 -33272 27935 -33210
rect 27615 -33508 27657 -33272
rect 27893 -33508 27935 -33272
rect 27615 -33592 27935 -33508
rect 27615 -33828 27657 -33592
rect 27893 -33828 27935 -33592
rect 27615 -33890 27935 -33828
rect 28615 -33272 28935 -33210
rect 28615 -33508 28657 -33272
rect 28893 -33508 28935 -33272
rect 28615 -33592 28935 -33508
rect 28615 -33828 28657 -33592
rect 28893 -33828 28935 -33592
rect 28615 -33890 28935 -33828
rect 29615 -33272 29935 -33210
rect 29615 -33508 29657 -33272
rect 29893 -33508 29935 -33272
rect 29615 -33592 29935 -33508
rect 29615 -33828 29657 -33592
rect 29893 -33828 29935 -33592
rect 29615 -33890 29935 -33828
rect 30615 -33272 30935 -33210
rect 30615 -33508 30657 -33272
rect 30893 -33508 30935 -33272
rect 30615 -33592 30935 -33508
rect 30615 -33828 30657 -33592
rect 30893 -33828 30935 -33592
rect 30615 -33890 30935 -33828
rect 31615 -33272 31935 -33210
rect 31615 -33508 31657 -33272
rect 31893 -33508 31935 -33272
rect 31615 -33592 31935 -33508
rect 31615 -33828 31657 -33592
rect 31893 -33828 31935 -33592
rect 31615 -33890 31935 -33828
rect 32615 -33272 32935 -33210
rect 32615 -33508 32657 -33272
rect 32893 -33508 32935 -33272
rect 32615 -33592 32935 -33508
rect 32615 -33828 32657 -33592
rect 32893 -33828 32935 -33592
rect 32615 -33890 32935 -33828
rect 33615 -33272 33935 -33210
rect 33615 -33508 33657 -33272
rect 33893 -33508 33935 -33272
rect 33615 -33592 33935 -33508
rect 33615 -33828 33657 -33592
rect 33893 -33828 33935 -33592
rect 33615 -33890 33935 -33828
rect 8275 -33932 34275 -33890
rect 8275 -34168 8317 -33932
rect 8553 -34168 8657 -33932
rect 8893 -34168 8997 -33932
rect 9233 -34168 9317 -33932
rect 9553 -34168 9657 -33932
rect 9893 -34168 9997 -33932
rect 10233 -34168 10317 -33932
rect 10553 -34168 10657 -33932
rect 10893 -34168 10997 -33932
rect 11233 -34168 11317 -33932
rect 11553 -34168 11657 -33932
rect 11893 -34168 11997 -33932
rect 12233 -34168 12317 -33932
rect 12553 -34168 12657 -33932
rect 12893 -34168 12997 -33932
rect 13233 -34168 13317 -33932
rect 13553 -34168 13657 -33932
rect 13893 -34168 13997 -33932
rect 14233 -34168 14317 -33932
rect 14553 -34168 14657 -33932
rect 14893 -34168 14997 -33932
rect 15233 -34168 15317 -33932
rect 15553 -34168 15657 -33932
rect 15893 -34168 15997 -33932
rect 16233 -34168 16317 -33932
rect 16553 -34168 16657 -33932
rect 16893 -34168 16997 -33932
rect 17233 -34168 17317 -33932
rect 17553 -34168 17657 -33932
rect 17893 -34168 17997 -33932
rect 18233 -34168 18317 -33932
rect 18553 -34168 18657 -33932
rect 18893 -34168 18997 -33932
rect 19233 -34168 19317 -33932
rect 19553 -34168 19657 -33932
rect 19893 -34168 19997 -33932
rect 20233 -34168 20317 -33932
rect 20553 -34168 20657 -33932
rect 20893 -34168 20997 -33932
rect 21233 -34168 21317 -33932
rect 21553 -34168 21657 -33932
rect 21893 -34168 21997 -33932
rect 22233 -34168 22317 -33932
rect 22553 -34168 22657 -33932
rect 22893 -34168 22997 -33932
rect 23233 -34168 23317 -33932
rect 23553 -34168 23657 -33932
rect 23893 -34168 23997 -33932
rect 24233 -34168 24317 -33932
rect 24553 -34168 24657 -33932
rect 24893 -34168 24997 -33932
rect 25233 -34168 25317 -33932
rect 25553 -34168 25657 -33932
rect 25893 -34168 25997 -33932
rect 26233 -34168 26317 -33932
rect 26553 -34168 26657 -33932
rect 26893 -34168 26997 -33932
rect 27233 -34168 27317 -33932
rect 27553 -34168 27657 -33932
rect 27893 -34168 27997 -33932
rect 28233 -34168 28317 -33932
rect 28553 -34168 28657 -33932
rect 28893 -34168 28997 -33932
rect 29233 -34168 29317 -33932
rect 29553 -34168 29657 -33932
rect 29893 -34168 29997 -33932
rect 30233 -34168 30317 -33932
rect 30553 -34168 30657 -33932
rect 30893 -34168 30997 -33932
rect 31233 -34168 31317 -33932
rect 31553 -34168 31657 -33932
rect 31893 -34168 31997 -33932
rect 32233 -34168 32317 -33932
rect 32553 -34168 32657 -33932
rect 32893 -34168 32997 -33932
rect 33233 -34168 33317 -33932
rect 33553 -34168 33657 -33932
rect 33893 -34168 33997 -33932
rect 34233 -34168 34275 -33932
rect 8275 -34210 34275 -34168
rect 8615 -34272 8935 -34210
rect 8615 -34508 8657 -34272
rect 8893 -34508 8935 -34272
rect 8615 -34592 8935 -34508
rect 8615 -34828 8657 -34592
rect 8893 -34828 8935 -34592
rect 8615 -34890 8935 -34828
rect 9615 -34272 9935 -34210
rect 9615 -34508 9657 -34272
rect 9893 -34508 9935 -34272
rect 9615 -34592 9935 -34508
rect 9615 -34828 9657 -34592
rect 9893 -34828 9935 -34592
rect 9615 -34890 9935 -34828
rect 10615 -34272 10935 -34210
rect 10615 -34508 10657 -34272
rect 10893 -34508 10935 -34272
rect 10615 -34592 10935 -34508
rect 10615 -34828 10657 -34592
rect 10893 -34828 10935 -34592
rect 10615 -34890 10935 -34828
rect 11615 -34272 11935 -34210
rect 11615 -34508 11657 -34272
rect 11893 -34508 11935 -34272
rect 11615 -34592 11935 -34508
rect 11615 -34828 11657 -34592
rect 11893 -34828 11935 -34592
rect 11615 -34890 11935 -34828
rect 12615 -34272 12935 -34210
rect 12615 -34508 12657 -34272
rect 12893 -34508 12935 -34272
rect 12615 -34592 12935 -34508
rect 12615 -34828 12657 -34592
rect 12893 -34828 12935 -34592
rect 12615 -34890 12935 -34828
rect 13615 -34272 13935 -34210
rect 13615 -34508 13657 -34272
rect 13893 -34508 13935 -34272
rect 13615 -34592 13935 -34508
rect 13615 -34828 13657 -34592
rect 13893 -34828 13935 -34592
rect 13615 -34890 13935 -34828
rect 14615 -34272 14935 -34210
rect 14615 -34508 14657 -34272
rect 14893 -34508 14935 -34272
rect 14615 -34592 14935 -34508
rect 14615 -34828 14657 -34592
rect 14893 -34828 14935 -34592
rect 14615 -34890 14935 -34828
rect 15615 -34272 15935 -34210
rect 15615 -34508 15657 -34272
rect 15893 -34508 15935 -34272
rect 15615 -34592 15935 -34508
rect 15615 -34828 15657 -34592
rect 15893 -34828 15935 -34592
rect 15615 -34890 15935 -34828
rect 16615 -34272 16935 -34210
rect 16615 -34508 16657 -34272
rect 16893 -34508 16935 -34272
rect 16615 -34592 16935 -34508
rect 16615 -34828 16657 -34592
rect 16893 -34828 16935 -34592
rect 16615 -34890 16935 -34828
rect 17615 -34272 17935 -34210
rect 17615 -34508 17657 -34272
rect 17893 -34508 17935 -34272
rect 17615 -34592 17935 -34508
rect 17615 -34828 17657 -34592
rect 17893 -34828 17935 -34592
rect 17615 -34890 17935 -34828
rect 18615 -34272 18935 -34210
rect 18615 -34508 18657 -34272
rect 18893 -34508 18935 -34272
rect 18615 -34592 18935 -34508
rect 18615 -34828 18657 -34592
rect 18893 -34828 18935 -34592
rect 18615 -34890 18935 -34828
rect 19615 -34272 19935 -34210
rect 19615 -34508 19657 -34272
rect 19893 -34508 19935 -34272
rect 19615 -34592 19935 -34508
rect 19615 -34828 19657 -34592
rect 19893 -34828 19935 -34592
rect 19615 -34890 19935 -34828
rect 20615 -34272 20935 -34210
rect 20615 -34508 20657 -34272
rect 20893 -34508 20935 -34272
rect 20615 -34592 20935 -34508
rect 20615 -34828 20657 -34592
rect 20893 -34828 20935 -34592
rect 20615 -34890 20935 -34828
rect 21615 -34272 21935 -34210
rect 21615 -34508 21657 -34272
rect 21893 -34508 21935 -34272
rect 21615 -34592 21935 -34508
rect 21615 -34828 21657 -34592
rect 21893 -34828 21935 -34592
rect 21615 -34890 21935 -34828
rect 22615 -34272 22935 -34210
rect 22615 -34508 22657 -34272
rect 22893 -34508 22935 -34272
rect 22615 -34592 22935 -34508
rect 22615 -34828 22657 -34592
rect 22893 -34828 22935 -34592
rect 22615 -34890 22935 -34828
rect 23615 -34272 23935 -34210
rect 23615 -34508 23657 -34272
rect 23893 -34508 23935 -34272
rect 23615 -34592 23935 -34508
rect 23615 -34828 23657 -34592
rect 23893 -34828 23935 -34592
rect 23615 -34890 23935 -34828
rect 24615 -34272 24935 -34210
rect 24615 -34508 24657 -34272
rect 24893 -34508 24935 -34272
rect 24615 -34592 24935 -34508
rect 24615 -34828 24657 -34592
rect 24893 -34828 24935 -34592
rect 24615 -34890 24935 -34828
rect 25615 -34272 25935 -34210
rect 25615 -34508 25657 -34272
rect 25893 -34508 25935 -34272
rect 25615 -34592 25935 -34508
rect 25615 -34828 25657 -34592
rect 25893 -34828 25935 -34592
rect 25615 -34890 25935 -34828
rect 26615 -34272 26935 -34210
rect 26615 -34508 26657 -34272
rect 26893 -34508 26935 -34272
rect 26615 -34592 26935 -34508
rect 26615 -34828 26657 -34592
rect 26893 -34828 26935 -34592
rect 26615 -34890 26935 -34828
rect 27615 -34272 27935 -34210
rect 27615 -34508 27657 -34272
rect 27893 -34508 27935 -34272
rect 27615 -34592 27935 -34508
rect 27615 -34828 27657 -34592
rect 27893 -34828 27935 -34592
rect 27615 -34890 27935 -34828
rect 28615 -34272 28935 -34210
rect 28615 -34508 28657 -34272
rect 28893 -34508 28935 -34272
rect 28615 -34592 28935 -34508
rect 28615 -34828 28657 -34592
rect 28893 -34828 28935 -34592
rect 28615 -34890 28935 -34828
rect 29615 -34272 29935 -34210
rect 29615 -34508 29657 -34272
rect 29893 -34508 29935 -34272
rect 29615 -34592 29935 -34508
rect 29615 -34828 29657 -34592
rect 29893 -34828 29935 -34592
rect 29615 -34890 29935 -34828
rect 30615 -34272 30935 -34210
rect 30615 -34508 30657 -34272
rect 30893 -34508 30935 -34272
rect 30615 -34592 30935 -34508
rect 30615 -34828 30657 -34592
rect 30893 -34828 30935 -34592
rect 30615 -34890 30935 -34828
rect 31615 -34272 31935 -34210
rect 31615 -34508 31657 -34272
rect 31893 -34508 31935 -34272
rect 31615 -34592 31935 -34508
rect 31615 -34828 31657 -34592
rect 31893 -34828 31935 -34592
rect 31615 -34890 31935 -34828
rect 32615 -34272 32935 -34210
rect 32615 -34508 32657 -34272
rect 32893 -34508 32935 -34272
rect 32615 -34592 32935 -34508
rect 32615 -34828 32657 -34592
rect 32893 -34828 32935 -34592
rect 32615 -34890 32935 -34828
rect 33615 -34272 33935 -34210
rect 33615 -34508 33657 -34272
rect 33893 -34508 33935 -34272
rect 33615 -34592 33935 -34508
rect 33615 -34828 33657 -34592
rect 33893 -34828 33935 -34592
rect 33615 -34890 33935 -34828
rect 8275 -34932 34275 -34890
rect 8275 -35168 8317 -34932
rect 8553 -35168 8657 -34932
rect 8893 -35168 8997 -34932
rect 9233 -35168 9317 -34932
rect 9553 -35168 9657 -34932
rect 9893 -35168 9997 -34932
rect 10233 -35168 10317 -34932
rect 10553 -35168 10657 -34932
rect 10893 -35168 10997 -34932
rect 11233 -35168 11317 -34932
rect 11553 -35168 11657 -34932
rect 11893 -35168 11997 -34932
rect 12233 -35168 12317 -34932
rect 12553 -35168 12657 -34932
rect 12893 -35168 12997 -34932
rect 13233 -35168 13317 -34932
rect 13553 -35168 13657 -34932
rect 13893 -35168 13997 -34932
rect 14233 -35168 14317 -34932
rect 14553 -35168 14657 -34932
rect 14893 -35168 14997 -34932
rect 15233 -35168 15317 -34932
rect 15553 -35168 15657 -34932
rect 15893 -35168 15997 -34932
rect 16233 -35168 16317 -34932
rect 16553 -35168 16657 -34932
rect 16893 -35168 16997 -34932
rect 17233 -35168 17317 -34932
rect 17553 -35168 17657 -34932
rect 17893 -35168 17997 -34932
rect 18233 -35168 18317 -34932
rect 18553 -35168 18657 -34932
rect 18893 -35168 18997 -34932
rect 19233 -35168 19317 -34932
rect 19553 -35168 19657 -34932
rect 19893 -35168 19997 -34932
rect 20233 -35168 20317 -34932
rect 20553 -35168 20657 -34932
rect 20893 -35168 20997 -34932
rect 21233 -35168 21317 -34932
rect 21553 -35168 21657 -34932
rect 21893 -35168 21997 -34932
rect 22233 -35168 22317 -34932
rect 22553 -35168 22657 -34932
rect 22893 -35168 22997 -34932
rect 23233 -35168 23317 -34932
rect 23553 -35168 23657 -34932
rect 23893 -35168 23997 -34932
rect 24233 -35168 24317 -34932
rect 24553 -35168 24657 -34932
rect 24893 -35168 24997 -34932
rect 25233 -35168 25317 -34932
rect 25553 -35168 25657 -34932
rect 25893 -35168 25997 -34932
rect 26233 -35168 26317 -34932
rect 26553 -35168 26657 -34932
rect 26893 -35168 26997 -34932
rect 27233 -35168 27317 -34932
rect 27553 -35168 27657 -34932
rect 27893 -35168 27997 -34932
rect 28233 -35168 28317 -34932
rect 28553 -35168 28657 -34932
rect 28893 -35168 28997 -34932
rect 29233 -35168 29317 -34932
rect 29553 -35168 29657 -34932
rect 29893 -35168 29997 -34932
rect 30233 -35168 30317 -34932
rect 30553 -35168 30657 -34932
rect 30893 -35168 30997 -34932
rect 31233 -35168 31317 -34932
rect 31553 -35168 31657 -34932
rect 31893 -35168 31997 -34932
rect 32233 -35168 32317 -34932
rect 32553 -35168 32657 -34932
rect 32893 -35168 32997 -34932
rect 33233 -35168 33317 -34932
rect 33553 -35168 33657 -34932
rect 33893 -35168 33997 -34932
rect 34233 -35168 34275 -34932
rect 8275 -35210 34275 -35168
rect 8615 -35272 8935 -35210
rect 8615 -35508 8657 -35272
rect 8893 -35508 8935 -35272
rect 8615 -35592 8935 -35508
rect 8615 -35828 8657 -35592
rect 8893 -35828 8935 -35592
rect 8615 -35890 8935 -35828
rect 9615 -35272 9935 -35210
rect 9615 -35508 9657 -35272
rect 9893 -35508 9935 -35272
rect 9615 -35592 9935 -35508
rect 9615 -35828 9657 -35592
rect 9893 -35828 9935 -35592
rect 9615 -35890 9935 -35828
rect 10615 -35272 10935 -35210
rect 10615 -35508 10657 -35272
rect 10893 -35508 10935 -35272
rect 10615 -35592 10935 -35508
rect 10615 -35828 10657 -35592
rect 10893 -35828 10935 -35592
rect 10615 -35890 10935 -35828
rect 11615 -35272 11935 -35210
rect 11615 -35508 11657 -35272
rect 11893 -35508 11935 -35272
rect 11615 -35592 11935 -35508
rect 11615 -35828 11657 -35592
rect 11893 -35828 11935 -35592
rect 11615 -35890 11935 -35828
rect 12615 -35272 12935 -35210
rect 12615 -35508 12657 -35272
rect 12893 -35508 12935 -35272
rect 12615 -35592 12935 -35508
rect 12615 -35828 12657 -35592
rect 12893 -35828 12935 -35592
rect 12615 -35890 12935 -35828
rect 13615 -35272 13935 -35210
rect 13615 -35508 13657 -35272
rect 13893 -35508 13935 -35272
rect 13615 -35592 13935 -35508
rect 13615 -35828 13657 -35592
rect 13893 -35828 13935 -35592
rect 13615 -35890 13935 -35828
rect 14615 -35272 14935 -35210
rect 14615 -35508 14657 -35272
rect 14893 -35508 14935 -35272
rect 14615 -35592 14935 -35508
rect 14615 -35828 14657 -35592
rect 14893 -35828 14935 -35592
rect 14615 -35890 14935 -35828
rect 15615 -35272 15935 -35210
rect 15615 -35508 15657 -35272
rect 15893 -35508 15935 -35272
rect 15615 -35592 15935 -35508
rect 15615 -35828 15657 -35592
rect 15893 -35828 15935 -35592
rect 15615 -35890 15935 -35828
rect 16615 -35272 16935 -35210
rect 16615 -35508 16657 -35272
rect 16893 -35508 16935 -35272
rect 16615 -35592 16935 -35508
rect 16615 -35828 16657 -35592
rect 16893 -35828 16935 -35592
rect 16615 -35890 16935 -35828
rect 17615 -35272 17935 -35210
rect 17615 -35508 17657 -35272
rect 17893 -35508 17935 -35272
rect 17615 -35592 17935 -35508
rect 17615 -35828 17657 -35592
rect 17893 -35828 17935 -35592
rect 17615 -35890 17935 -35828
rect 18615 -35272 18935 -35210
rect 18615 -35508 18657 -35272
rect 18893 -35508 18935 -35272
rect 18615 -35592 18935 -35508
rect 18615 -35828 18657 -35592
rect 18893 -35828 18935 -35592
rect 18615 -35890 18935 -35828
rect 19615 -35272 19935 -35210
rect 19615 -35508 19657 -35272
rect 19893 -35508 19935 -35272
rect 19615 -35592 19935 -35508
rect 19615 -35828 19657 -35592
rect 19893 -35828 19935 -35592
rect 19615 -35890 19935 -35828
rect 20615 -35272 20935 -35210
rect 20615 -35508 20657 -35272
rect 20893 -35508 20935 -35272
rect 20615 -35592 20935 -35508
rect 20615 -35828 20657 -35592
rect 20893 -35828 20935 -35592
rect 20615 -35890 20935 -35828
rect 21615 -35272 21935 -35210
rect 21615 -35508 21657 -35272
rect 21893 -35508 21935 -35272
rect 21615 -35592 21935 -35508
rect 21615 -35828 21657 -35592
rect 21893 -35828 21935 -35592
rect 21615 -35890 21935 -35828
rect 22615 -35272 22935 -35210
rect 22615 -35508 22657 -35272
rect 22893 -35508 22935 -35272
rect 22615 -35592 22935 -35508
rect 22615 -35828 22657 -35592
rect 22893 -35828 22935 -35592
rect 22615 -35890 22935 -35828
rect 23615 -35272 23935 -35210
rect 23615 -35508 23657 -35272
rect 23893 -35508 23935 -35272
rect 23615 -35592 23935 -35508
rect 23615 -35828 23657 -35592
rect 23893 -35828 23935 -35592
rect 23615 -35890 23935 -35828
rect 24615 -35272 24935 -35210
rect 24615 -35508 24657 -35272
rect 24893 -35508 24935 -35272
rect 24615 -35592 24935 -35508
rect 24615 -35828 24657 -35592
rect 24893 -35828 24935 -35592
rect 24615 -35890 24935 -35828
rect 25615 -35272 25935 -35210
rect 25615 -35508 25657 -35272
rect 25893 -35508 25935 -35272
rect 25615 -35592 25935 -35508
rect 25615 -35828 25657 -35592
rect 25893 -35828 25935 -35592
rect 25615 -35890 25935 -35828
rect 26615 -35272 26935 -35210
rect 26615 -35508 26657 -35272
rect 26893 -35508 26935 -35272
rect 26615 -35592 26935 -35508
rect 26615 -35828 26657 -35592
rect 26893 -35828 26935 -35592
rect 26615 -35890 26935 -35828
rect 27615 -35272 27935 -35210
rect 27615 -35508 27657 -35272
rect 27893 -35508 27935 -35272
rect 27615 -35592 27935 -35508
rect 27615 -35828 27657 -35592
rect 27893 -35828 27935 -35592
rect 27615 -35890 27935 -35828
rect 28615 -35272 28935 -35210
rect 28615 -35508 28657 -35272
rect 28893 -35508 28935 -35272
rect 28615 -35592 28935 -35508
rect 28615 -35828 28657 -35592
rect 28893 -35828 28935 -35592
rect 28615 -35890 28935 -35828
rect 29615 -35272 29935 -35210
rect 29615 -35508 29657 -35272
rect 29893 -35508 29935 -35272
rect 29615 -35592 29935 -35508
rect 29615 -35828 29657 -35592
rect 29893 -35828 29935 -35592
rect 29615 -35890 29935 -35828
rect 30615 -35272 30935 -35210
rect 30615 -35508 30657 -35272
rect 30893 -35508 30935 -35272
rect 30615 -35592 30935 -35508
rect 30615 -35828 30657 -35592
rect 30893 -35828 30935 -35592
rect 30615 -35890 30935 -35828
rect 31615 -35272 31935 -35210
rect 31615 -35508 31657 -35272
rect 31893 -35508 31935 -35272
rect 31615 -35592 31935 -35508
rect 31615 -35828 31657 -35592
rect 31893 -35828 31935 -35592
rect 31615 -35890 31935 -35828
rect 32615 -35272 32935 -35210
rect 32615 -35508 32657 -35272
rect 32893 -35508 32935 -35272
rect 32615 -35592 32935 -35508
rect 32615 -35828 32657 -35592
rect 32893 -35828 32935 -35592
rect 32615 -35890 32935 -35828
rect 33615 -35272 33935 -35210
rect 33615 -35508 33657 -35272
rect 33893 -35508 33935 -35272
rect 33615 -35592 33935 -35508
rect 33615 -35828 33657 -35592
rect 33893 -35828 33935 -35592
rect 33615 -35890 33935 -35828
rect 8275 -35932 34275 -35890
rect 8275 -36168 8317 -35932
rect 8553 -36168 8657 -35932
rect 8893 -36168 8997 -35932
rect 9233 -36168 9317 -35932
rect 9553 -36168 9657 -35932
rect 9893 -36168 9997 -35932
rect 10233 -36168 10317 -35932
rect 10553 -36168 10657 -35932
rect 10893 -36168 10997 -35932
rect 11233 -36168 11317 -35932
rect 11553 -36168 11657 -35932
rect 11893 -36168 11997 -35932
rect 12233 -36168 12317 -35932
rect 12553 -36168 12657 -35932
rect 12893 -36168 12997 -35932
rect 13233 -36168 13317 -35932
rect 13553 -36168 13657 -35932
rect 13893 -36168 13997 -35932
rect 14233 -36168 14317 -35932
rect 14553 -36168 14657 -35932
rect 14893 -36168 14997 -35932
rect 15233 -36168 15317 -35932
rect 15553 -36168 15657 -35932
rect 15893 -36168 15997 -35932
rect 16233 -36168 16317 -35932
rect 16553 -36168 16657 -35932
rect 16893 -36168 16997 -35932
rect 17233 -36168 17317 -35932
rect 17553 -36168 17657 -35932
rect 17893 -36168 17997 -35932
rect 18233 -36168 18317 -35932
rect 18553 -36168 18657 -35932
rect 18893 -36168 18997 -35932
rect 19233 -36168 19317 -35932
rect 19553 -36168 19657 -35932
rect 19893 -36168 19997 -35932
rect 20233 -36168 20317 -35932
rect 20553 -36168 20657 -35932
rect 20893 -36168 20997 -35932
rect 21233 -36168 21317 -35932
rect 21553 -36168 21657 -35932
rect 21893 -36168 21997 -35932
rect 22233 -36168 22317 -35932
rect 22553 -36168 22657 -35932
rect 22893 -36168 22997 -35932
rect 23233 -36168 23317 -35932
rect 23553 -36168 23657 -35932
rect 23893 -36168 23997 -35932
rect 24233 -36168 24317 -35932
rect 24553 -36168 24657 -35932
rect 24893 -36168 24997 -35932
rect 25233 -36168 25317 -35932
rect 25553 -36168 25657 -35932
rect 25893 -36168 25997 -35932
rect 26233 -36168 26317 -35932
rect 26553 -36168 26657 -35932
rect 26893 -36168 26997 -35932
rect 27233 -36168 27317 -35932
rect 27553 -36168 27657 -35932
rect 27893 -36168 27997 -35932
rect 28233 -36168 28317 -35932
rect 28553 -36168 28657 -35932
rect 28893 -36168 28997 -35932
rect 29233 -36168 29317 -35932
rect 29553 -36168 29657 -35932
rect 29893 -36168 29997 -35932
rect 30233 -36168 30317 -35932
rect 30553 -36168 30657 -35932
rect 30893 -36168 30997 -35932
rect 31233 -36168 31317 -35932
rect 31553 -36168 31657 -35932
rect 31893 -36168 31997 -35932
rect 32233 -36168 32317 -35932
rect 32553 -36168 32657 -35932
rect 32893 -36168 32997 -35932
rect 33233 -36168 33317 -35932
rect 33553 -36168 33657 -35932
rect 33893 -36168 33997 -35932
rect 34233 -36168 34275 -35932
rect 8275 -36210 34275 -36168
rect 8615 -36272 8935 -36210
rect 8615 -36508 8657 -36272
rect 8893 -36508 8935 -36272
rect 8615 -36592 8935 -36508
rect 8615 -36828 8657 -36592
rect 8893 -36828 8935 -36592
rect 8615 -36890 8935 -36828
rect 9615 -36272 9935 -36210
rect 9615 -36508 9657 -36272
rect 9893 -36508 9935 -36272
rect 9615 -36592 9935 -36508
rect 9615 -36828 9657 -36592
rect 9893 -36828 9935 -36592
rect 9615 -36890 9935 -36828
rect 10615 -36272 10935 -36210
rect 10615 -36508 10657 -36272
rect 10893 -36508 10935 -36272
rect 10615 -36592 10935 -36508
rect 10615 -36828 10657 -36592
rect 10893 -36828 10935 -36592
rect 10615 -36890 10935 -36828
rect 11615 -36272 11935 -36210
rect 11615 -36508 11657 -36272
rect 11893 -36508 11935 -36272
rect 11615 -36592 11935 -36508
rect 11615 -36828 11657 -36592
rect 11893 -36828 11935 -36592
rect 11615 -36890 11935 -36828
rect 12615 -36272 12935 -36210
rect 12615 -36508 12657 -36272
rect 12893 -36508 12935 -36272
rect 12615 -36592 12935 -36508
rect 12615 -36828 12657 -36592
rect 12893 -36828 12935 -36592
rect 12615 -36890 12935 -36828
rect 13615 -36272 13935 -36210
rect 13615 -36508 13657 -36272
rect 13893 -36508 13935 -36272
rect 13615 -36592 13935 -36508
rect 13615 -36828 13657 -36592
rect 13893 -36828 13935 -36592
rect 13615 -36890 13935 -36828
rect 14615 -36272 14935 -36210
rect 14615 -36508 14657 -36272
rect 14893 -36508 14935 -36272
rect 14615 -36592 14935 -36508
rect 14615 -36828 14657 -36592
rect 14893 -36828 14935 -36592
rect 14615 -36890 14935 -36828
rect 15615 -36272 15935 -36210
rect 15615 -36508 15657 -36272
rect 15893 -36508 15935 -36272
rect 15615 -36592 15935 -36508
rect 15615 -36828 15657 -36592
rect 15893 -36828 15935 -36592
rect 15615 -36890 15935 -36828
rect 16615 -36272 16935 -36210
rect 16615 -36508 16657 -36272
rect 16893 -36508 16935 -36272
rect 16615 -36592 16935 -36508
rect 16615 -36828 16657 -36592
rect 16893 -36828 16935 -36592
rect 16615 -36890 16935 -36828
rect 17615 -36272 17935 -36210
rect 17615 -36508 17657 -36272
rect 17893 -36508 17935 -36272
rect 17615 -36592 17935 -36508
rect 17615 -36828 17657 -36592
rect 17893 -36828 17935 -36592
rect 17615 -36890 17935 -36828
rect 18615 -36272 18935 -36210
rect 18615 -36508 18657 -36272
rect 18893 -36508 18935 -36272
rect 18615 -36592 18935 -36508
rect 18615 -36828 18657 -36592
rect 18893 -36828 18935 -36592
rect 18615 -36890 18935 -36828
rect 19615 -36272 19935 -36210
rect 19615 -36508 19657 -36272
rect 19893 -36508 19935 -36272
rect 19615 -36592 19935 -36508
rect 19615 -36828 19657 -36592
rect 19893 -36828 19935 -36592
rect 19615 -36890 19935 -36828
rect 20615 -36272 20935 -36210
rect 20615 -36508 20657 -36272
rect 20893 -36508 20935 -36272
rect 20615 -36592 20935 -36508
rect 20615 -36828 20657 -36592
rect 20893 -36828 20935 -36592
rect 20615 -36890 20935 -36828
rect 21615 -36272 21935 -36210
rect 21615 -36508 21657 -36272
rect 21893 -36508 21935 -36272
rect 21615 -36592 21935 -36508
rect 21615 -36828 21657 -36592
rect 21893 -36828 21935 -36592
rect 21615 -36890 21935 -36828
rect 22615 -36272 22935 -36210
rect 22615 -36508 22657 -36272
rect 22893 -36508 22935 -36272
rect 22615 -36592 22935 -36508
rect 22615 -36828 22657 -36592
rect 22893 -36828 22935 -36592
rect 22615 -36890 22935 -36828
rect 23615 -36272 23935 -36210
rect 23615 -36508 23657 -36272
rect 23893 -36508 23935 -36272
rect 23615 -36592 23935 -36508
rect 23615 -36828 23657 -36592
rect 23893 -36828 23935 -36592
rect 23615 -36890 23935 -36828
rect 24615 -36272 24935 -36210
rect 24615 -36508 24657 -36272
rect 24893 -36508 24935 -36272
rect 24615 -36592 24935 -36508
rect 24615 -36828 24657 -36592
rect 24893 -36828 24935 -36592
rect 24615 -36890 24935 -36828
rect 25615 -36272 25935 -36210
rect 25615 -36508 25657 -36272
rect 25893 -36508 25935 -36272
rect 25615 -36592 25935 -36508
rect 25615 -36828 25657 -36592
rect 25893 -36828 25935 -36592
rect 25615 -36890 25935 -36828
rect 26615 -36272 26935 -36210
rect 26615 -36508 26657 -36272
rect 26893 -36508 26935 -36272
rect 26615 -36592 26935 -36508
rect 26615 -36828 26657 -36592
rect 26893 -36828 26935 -36592
rect 26615 -36890 26935 -36828
rect 27615 -36272 27935 -36210
rect 27615 -36508 27657 -36272
rect 27893 -36508 27935 -36272
rect 27615 -36592 27935 -36508
rect 27615 -36828 27657 -36592
rect 27893 -36828 27935 -36592
rect 27615 -36890 27935 -36828
rect 28615 -36272 28935 -36210
rect 28615 -36508 28657 -36272
rect 28893 -36508 28935 -36272
rect 28615 -36592 28935 -36508
rect 28615 -36828 28657 -36592
rect 28893 -36828 28935 -36592
rect 28615 -36890 28935 -36828
rect 29615 -36272 29935 -36210
rect 29615 -36508 29657 -36272
rect 29893 -36508 29935 -36272
rect 29615 -36592 29935 -36508
rect 29615 -36828 29657 -36592
rect 29893 -36828 29935 -36592
rect 29615 -36890 29935 -36828
rect 30615 -36272 30935 -36210
rect 30615 -36508 30657 -36272
rect 30893 -36508 30935 -36272
rect 30615 -36592 30935 -36508
rect 30615 -36828 30657 -36592
rect 30893 -36828 30935 -36592
rect 30615 -36890 30935 -36828
rect 31615 -36272 31935 -36210
rect 31615 -36508 31657 -36272
rect 31893 -36508 31935 -36272
rect 31615 -36592 31935 -36508
rect 31615 -36828 31657 -36592
rect 31893 -36828 31935 -36592
rect 31615 -36890 31935 -36828
rect 32615 -36272 32935 -36210
rect 32615 -36508 32657 -36272
rect 32893 -36508 32935 -36272
rect 32615 -36592 32935 -36508
rect 32615 -36828 32657 -36592
rect 32893 -36828 32935 -36592
rect 32615 -36890 32935 -36828
rect 33615 -36272 33935 -36210
rect 33615 -36508 33657 -36272
rect 33893 -36508 33935 -36272
rect 33615 -36592 33935 -36508
rect 33615 -36828 33657 -36592
rect 33893 -36828 33935 -36592
rect 33615 -36890 33935 -36828
rect 8275 -36932 34275 -36890
rect 8275 -37168 8317 -36932
rect 8553 -37168 8657 -36932
rect 8893 -37168 8997 -36932
rect 9233 -37168 9317 -36932
rect 9553 -37168 9657 -36932
rect 9893 -37168 9997 -36932
rect 10233 -37168 10317 -36932
rect 10553 -37168 10657 -36932
rect 10893 -37168 10997 -36932
rect 11233 -37168 11317 -36932
rect 11553 -37168 11657 -36932
rect 11893 -37168 11997 -36932
rect 12233 -37168 12317 -36932
rect 12553 -37168 12657 -36932
rect 12893 -37168 12997 -36932
rect 13233 -37168 13317 -36932
rect 13553 -37168 13657 -36932
rect 13893 -37168 13997 -36932
rect 14233 -37168 14317 -36932
rect 14553 -37168 14657 -36932
rect 14893 -37168 14997 -36932
rect 15233 -37168 15317 -36932
rect 15553 -37168 15657 -36932
rect 15893 -37168 15997 -36932
rect 16233 -37168 16317 -36932
rect 16553 -37168 16657 -36932
rect 16893 -37168 16997 -36932
rect 17233 -37168 17317 -36932
rect 17553 -37168 17657 -36932
rect 17893 -37168 17997 -36932
rect 18233 -37168 18317 -36932
rect 18553 -37168 18657 -36932
rect 18893 -37168 18997 -36932
rect 19233 -37168 19317 -36932
rect 19553 -37168 19657 -36932
rect 19893 -37168 19997 -36932
rect 20233 -37168 20317 -36932
rect 20553 -37168 20657 -36932
rect 20893 -37168 20997 -36932
rect 21233 -37168 21317 -36932
rect 21553 -37168 21657 -36932
rect 21893 -37168 21997 -36932
rect 22233 -37168 22317 -36932
rect 22553 -37168 22657 -36932
rect 22893 -37168 22997 -36932
rect 23233 -37168 23317 -36932
rect 23553 -37168 23657 -36932
rect 23893 -37168 23997 -36932
rect 24233 -37168 24317 -36932
rect 24553 -37168 24657 -36932
rect 24893 -37168 24997 -36932
rect 25233 -37168 25317 -36932
rect 25553 -37168 25657 -36932
rect 25893 -37168 25997 -36932
rect 26233 -37168 26317 -36932
rect 26553 -37168 26657 -36932
rect 26893 -37168 26997 -36932
rect 27233 -37168 27317 -36932
rect 27553 -37168 27657 -36932
rect 27893 -37168 27997 -36932
rect 28233 -37168 28317 -36932
rect 28553 -37168 28657 -36932
rect 28893 -37168 28997 -36932
rect 29233 -37168 29317 -36932
rect 29553 -37168 29657 -36932
rect 29893 -37168 29997 -36932
rect 30233 -37168 30317 -36932
rect 30553 -37168 30657 -36932
rect 30893 -37168 30997 -36932
rect 31233 -37168 31317 -36932
rect 31553 -37168 31657 -36932
rect 31893 -37168 31997 -36932
rect 32233 -37168 32317 -36932
rect 32553 -37168 32657 -36932
rect 32893 -37168 32997 -36932
rect 33233 -37168 33317 -36932
rect 33553 -37168 33657 -36932
rect 33893 -37168 33997 -36932
rect 34233 -37168 34275 -36932
rect 8275 -37210 34275 -37168
rect 8615 -37272 8935 -37210
rect 8615 -37508 8657 -37272
rect 8893 -37508 8935 -37272
rect 8615 -37592 8935 -37508
rect 8615 -37828 8657 -37592
rect 8893 -37828 8935 -37592
rect 8615 -37890 8935 -37828
rect 9615 -37272 9935 -37210
rect 9615 -37508 9657 -37272
rect 9893 -37508 9935 -37272
rect 9615 -37592 9935 -37508
rect 9615 -37828 9657 -37592
rect 9893 -37828 9935 -37592
rect 9615 -37890 9935 -37828
rect 10615 -37272 10935 -37210
rect 10615 -37508 10657 -37272
rect 10893 -37508 10935 -37272
rect 10615 -37592 10935 -37508
rect 10615 -37828 10657 -37592
rect 10893 -37828 10935 -37592
rect 10615 -37890 10935 -37828
rect 11615 -37272 11935 -37210
rect 11615 -37508 11657 -37272
rect 11893 -37508 11935 -37272
rect 11615 -37592 11935 -37508
rect 11615 -37828 11657 -37592
rect 11893 -37828 11935 -37592
rect 11615 -37890 11935 -37828
rect 12615 -37272 12935 -37210
rect 12615 -37508 12657 -37272
rect 12893 -37508 12935 -37272
rect 12615 -37592 12935 -37508
rect 12615 -37828 12657 -37592
rect 12893 -37828 12935 -37592
rect 12615 -37890 12935 -37828
rect 13615 -37272 13935 -37210
rect 13615 -37508 13657 -37272
rect 13893 -37508 13935 -37272
rect 13615 -37592 13935 -37508
rect 13615 -37828 13657 -37592
rect 13893 -37828 13935 -37592
rect 13615 -37890 13935 -37828
rect 14615 -37272 14935 -37210
rect 14615 -37508 14657 -37272
rect 14893 -37508 14935 -37272
rect 14615 -37592 14935 -37508
rect 14615 -37828 14657 -37592
rect 14893 -37828 14935 -37592
rect 14615 -37890 14935 -37828
rect 15615 -37272 15935 -37210
rect 15615 -37508 15657 -37272
rect 15893 -37508 15935 -37272
rect 15615 -37592 15935 -37508
rect 15615 -37828 15657 -37592
rect 15893 -37828 15935 -37592
rect 15615 -37890 15935 -37828
rect 16615 -37272 16935 -37210
rect 16615 -37508 16657 -37272
rect 16893 -37508 16935 -37272
rect 16615 -37592 16935 -37508
rect 16615 -37828 16657 -37592
rect 16893 -37828 16935 -37592
rect 16615 -37890 16935 -37828
rect 17615 -37272 17935 -37210
rect 17615 -37508 17657 -37272
rect 17893 -37508 17935 -37272
rect 17615 -37592 17935 -37508
rect 17615 -37828 17657 -37592
rect 17893 -37828 17935 -37592
rect 17615 -37890 17935 -37828
rect 18615 -37272 18935 -37210
rect 18615 -37508 18657 -37272
rect 18893 -37508 18935 -37272
rect 18615 -37592 18935 -37508
rect 18615 -37828 18657 -37592
rect 18893 -37828 18935 -37592
rect 18615 -37890 18935 -37828
rect 19615 -37272 19935 -37210
rect 19615 -37508 19657 -37272
rect 19893 -37508 19935 -37272
rect 19615 -37592 19935 -37508
rect 19615 -37828 19657 -37592
rect 19893 -37828 19935 -37592
rect 19615 -37890 19935 -37828
rect 20615 -37272 20935 -37210
rect 20615 -37508 20657 -37272
rect 20893 -37508 20935 -37272
rect 20615 -37592 20935 -37508
rect 20615 -37828 20657 -37592
rect 20893 -37828 20935 -37592
rect 20615 -37890 20935 -37828
rect 21615 -37272 21935 -37210
rect 21615 -37508 21657 -37272
rect 21893 -37508 21935 -37272
rect 21615 -37592 21935 -37508
rect 21615 -37828 21657 -37592
rect 21893 -37828 21935 -37592
rect 21615 -37890 21935 -37828
rect 22615 -37272 22935 -37210
rect 22615 -37508 22657 -37272
rect 22893 -37508 22935 -37272
rect 22615 -37592 22935 -37508
rect 22615 -37828 22657 -37592
rect 22893 -37828 22935 -37592
rect 22615 -37890 22935 -37828
rect 23615 -37272 23935 -37210
rect 23615 -37508 23657 -37272
rect 23893 -37508 23935 -37272
rect 23615 -37592 23935 -37508
rect 23615 -37828 23657 -37592
rect 23893 -37828 23935 -37592
rect 23615 -37890 23935 -37828
rect 24615 -37272 24935 -37210
rect 24615 -37508 24657 -37272
rect 24893 -37508 24935 -37272
rect 24615 -37592 24935 -37508
rect 24615 -37828 24657 -37592
rect 24893 -37828 24935 -37592
rect 24615 -37890 24935 -37828
rect 25615 -37272 25935 -37210
rect 25615 -37508 25657 -37272
rect 25893 -37508 25935 -37272
rect 25615 -37592 25935 -37508
rect 25615 -37828 25657 -37592
rect 25893 -37828 25935 -37592
rect 25615 -37890 25935 -37828
rect 26615 -37272 26935 -37210
rect 26615 -37508 26657 -37272
rect 26893 -37508 26935 -37272
rect 26615 -37592 26935 -37508
rect 26615 -37828 26657 -37592
rect 26893 -37828 26935 -37592
rect 26615 -37890 26935 -37828
rect 27615 -37272 27935 -37210
rect 27615 -37508 27657 -37272
rect 27893 -37508 27935 -37272
rect 27615 -37592 27935 -37508
rect 27615 -37828 27657 -37592
rect 27893 -37828 27935 -37592
rect 27615 -37890 27935 -37828
rect 28615 -37272 28935 -37210
rect 28615 -37508 28657 -37272
rect 28893 -37508 28935 -37272
rect 28615 -37592 28935 -37508
rect 28615 -37828 28657 -37592
rect 28893 -37828 28935 -37592
rect 28615 -37890 28935 -37828
rect 29615 -37272 29935 -37210
rect 29615 -37508 29657 -37272
rect 29893 -37508 29935 -37272
rect 29615 -37592 29935 -37508
rect 29615 -37828 29657 -37592
rect 29893 -37828 29935 -37592
rect 29615 -37890 29935 -37828
rect 30615 -37272 30935 -37210
rect 30615 -37508 30657 -37272
rect 30893 -37508 30935 -37272
rect 30615 -37592 30935 -37508
rect 30615 -37828 30657 -37592
rect 30893 -37828 30935 -37592
rect 30615 -37890 30935 -37828
rect 31615 -37272 31935 -37210
rect 31615 -37508 31657 -37272
rect 31893 -37508 31935 -37272
rect 31615 -37592 31935 -37508
rect 31615 -37828 31657 -37592
rect 31893 -37828 31935 -37592
rect 31615 -37890 31935 -37828
rect 32615 -37272 32935 -37210
rect 32615 -37508 32657 -37272
rect 32893 -37508 32935 -37272
rect 32615 -37592 32935 -37508
rect 32615 -37828 32657 -37592
rect 32893 -37828 32935 -37592
rect 32615 -37890 32935 -37828
rect 33615 -37272 33935 -37210
rect 33615 -37508 33657 -37272
rect 33893 -37508 33935 -37272
rect 33615 -37592 33935 -37508
rect 33615 -37828 33657 -37592
rect 33893 -37828 33935 -37592
rect 33615 -37890 33935 -37828
rect 8275 -37932 34275 -37890
rect 8275 -38168 8317 -37932
rect 8553 -38168 8657 -37932
rect 8893 -38168 8997 -37932
rect 9233 -38168 9317 -37932
rect 9553 -38168 9657 -37932
rect 9893 -38168 9997 -37932
rect 10233 -38168 10317 -37932
rect 10553 -38168 10657 -37932
rect 10893 -38168 10997 -37932
rect 11233 -38168 11317 -37932
rect 11553 -38168 11657 -37932
rect 11893 -38168 11997 -37932
rect 12233 -38168 12317 -37932
rect 12553 -38168 12657 -37932
rect 12893 -38168 12997 -37932
rect 13233 -38168 13317 -37932
rect 13553 -38168 13657 -37932
rect 13893 -38168 13997 -37932
rect 14233 -38168 14317 -37932
rect 14553 -38168 14657 -37932
rect 14893 -38168 14997 -37932
rect 15233 -38168 15317 -37932
rect 15553 -38168 15657 -37932
rect 15893 -38168 15997 -37932
rect 16233 -38168 16317 -37932
rect 16553 -38168 16657 -37932
rect 16893 -38168 16997 -37932
rect 17233 -38168 17317 -37932
rect 17553 -38168 17657 -37932
rect 17893 -38168 17997 -37932
rect 18233 -38168 18317 -37932
rect 18553 -38168 18657 -37932
rect 18893 -38168 18997 -37932
rect 19233 -38168 19317 -37932
rect 19553 -38168 19657 -37932
rect 19893 -38168 19997 -37932
rect 20233 -38168 20317 -37932
rect 20553 -38168 20657 -37932
rect 20893 -38168 20997 -37932
rect 21233 -38168 21317 -37932
rect 21553 -38168 21657 -37932
rect 21893 -38168 21997 -37932
rect 22233 -38168 22317 -37932
rect 22553 -38168 22657 -37932
rect 22893 -38168 22997 -37932
rect 23233 -38168 23317 -37932
rect 23553 -38168 23657 -37932
rect 23893 -38168 23997 -37932
rect 24233 -38168 24317 -37932
rect 24553 -38168 24657 -37932
rect 24893 -38168 24997 -37932
rect 25233 -38168 25317 -37932
rect 25553 -38168 25657 -37932
rect 25893 -38168 25997 -37932
rect 26233 -38168 26317 -37932
rect 26553 -38168 26657 -37932
rect 26893 -38168 26997 -37932
rect 27233 -38168 27317 -37932
rect 27553 -38168 27657 -37932
rect 27893 -38168 27997 -37932
rect 28233 -38168 28317 -37932
rect 28553 -38168 28657 -37932
rect 28893 -38168 28997 -37932
rect 29233 -38168 29317 -37932
rect 29553 -38168 29657 -37932
rect 29893 -38168 29997 -37932
rect 30233 -38168 30317 -37932
rect 30553 -38168 30657 -37932
rect 30893 -38168 30997 -37932
rect 31233 -38168 31317 -37932
rect 31553 -38168 31657 -37932
rect 31893 -38168 31997 -37932
rect 32233 -38168 32317 -37932
rect 32553 -38168 32657 -37932
rect 32893 -38168 32997 -37932
rect 33233 -38168 33317 -37932
rect 33553 -38168 33657 -37932
rect 33893 -38168 33997 -37932
rect 34233 -38168 34275 -37932
rect 8275 -38210 34275 -38168
rect 8615 -38272 8935 -38210
rect 8615 -38508 8657 -38272
rect 8893 -38508 8935 -38272
rect 8615 -38592 8935 -38508
rect 8615 -38828 8657 -38592
rect 8893 -38828 8935 -38592
rect 8615 -38890 8935 -38828
rect 9615 -38272 9935 -38210
rect 9615 -38508 9657 -38272
rect 9893 -38508 9935 -38272
rect 9615 -38592 9935 -38508
rect 9615 -38828 9657 -38592
rect 9893 -38828 9935 -38592
rect 9615 -38890 9935 -38828
rect 10615 -38272 10935 -38210
rect 10615 -38508 10657 -38272
rect 10893 -38508 10935 -38272
rect 10615 -38592 10935 -38508
rect 10615 -38828 10657 -38592
rect 10893 -38828 10935 -38592
rect 10615 -38890 10935 -38828
rect 11615 -38272 11935 -38210
rect 11615 -38508 11657 -38272
rect 11893 -38508 11935 -38272
rect 11615 -38592 11935 -38508
rect 11615 -38828 11657 -38592
rect 11893 -38828 11935 -38592
rect 11615 -38890 11935 -38828
rect 12615 -38272 12935 -38210
rect 12615 -38508 12657 -38272
rect 12893 -38508 12935 -38272
rect 12615 -38592 12935 -38508
rect 12615 -38828 12657 -38592
rect 12893 -38828 12935 -38592
rect 12615 -38890 12935 -38828
rect 13615 -38272 13935 -38210
rect 13615 -38508 13657 -38272
rect 13893 -38508 13935 -38272
rect 13615 -38592 13935 -38508
rect 13615 -38828 13657 -38592
rect 13893 -38828 13935 -38592
rect 13615 -38890 13935 -38828
rect 14615 -38272 14935 -38210
rect 14615 -38508 14657 -38272
rect 14893 -38508 14935 -38272
rect 14615 -38592 14935 -38508
rect 14615 -38828 14657 -38592
rect 14893 -38828 14935 -38592
rect 14615 -38890 14935 -38828
rect 15615 -38272 15935 -38210
rect 15615 -38508 15657 -38272
rect 15893 -38508 15935 -38272
rect 15615 -38592 15935 -38508
rect 15615 -38828 15657 -38592
rect 15893 -38828 15935 -38592
rect 15615 -38890 15935 -38828
rect 16615 -38272 16935 -38210
rect 16615 -38508 16657 -38272
rect 16893 -38508 16935 -38272
rect 16615 -38592 16935 -38508
rect 16615 -38828 16657 -38592
rect 16893 -38828 16935 -38592
rect 16615 -38890 16935 -38828
rect 17615 -38272 17935 -38210
rect 17615 -38508 17657 -38272
rect 17893 -38508 17935 -38272
rect 17615 -38592 17935 -38508
rect 17615 -38828 17657 -38592
rect 17893 -38828 17935 -38592
rect 17615 -38890 17935 -38828
rect 18615 -38272 18935 -38210
rect 18615 -38508 18657 -38272
rect 18893 -38508 18935 -38272
rect 18615 -38592 18935 -38508
rect 18615 -38828 18657 -38592
rect 18893 -38828 18935 -38592
rect 18615 -38890 18935 -38828
rect 19615 -38272 19935 -38210
rect 19615 -38508 19657 -38272
rect 19893 -38508 19935 -38272
rect 19615 -38592 19935 -38508
rect 19615 -38828 19657 -38592
rect 19893 -38828 19935 -38592
rect 19615 -38890 19935 -38828
rect 20615 -38272 20935 -38210
rect 20615 -38508 20657 -38272
rect 20893 -38508 20935 -38272
rect 20615 -38592 20935 -38508
rect 20615 -38828 20657 -38592
rect 20893 -38828 20935 -38592
rect 20615 -38890 20935 -38828
rect 21615 -38272 21935 -38210
rect 21615 -38508 21657 -38272
rect 21893 -38508 21935 -38272
rect 21615 -38592 21935 -38508
rect 21615 -38828 21657 -38592
rect 21893 -38828 21935 -38592
rect 21615 -38890 21935 -38828
rect 22615 -38272 22935 -38210
rect 22615 -38508 22657 -38272
rect 22893 -38508 22935 -38272
rect 22615 -38592 22935 -38508
rect 22615 -38828 22657 -38592
rect 22893 -38828 22935 -38592
rect 22615 -38890 22935 -38828
rect 23615 -38272 23935 -38210
rect 23615 -38508 23657 -38272
rect 23893 -38508 23935 -38272
rect 23615 -38592 23935 -38508
rect 23615 -38828 23657 -38592
rect 23893 -38828 23935 -38592
rect 23615 -38890 23935 -38828
rect 24615 -38272 24935 -38210
rect 24615 -38508 24657 -38272
rect 24893 -38508 24935 -38272
rect 24615 -38592 24935 -38508
rect 24615 -38828 24657 -38592
rect 24893 -38828 24935 -38592
rect 24615 -38890 24935 -38828
rect 25615 -38272 25935 -38210
rect 25615 -38508 25657 -38272
rect 25893 -38508 25935 -38272
rect 25615 -38592 25935 -38508
rect 25615 -38828 25657 -38592
rect 25893 -38828 25935 -38592
rect 25615 -38890 25935 -38828
rect 26615 -38272 26935 -38210
rect 26615 -38508 26657 -38272
rect 26893 -38508 26935 -38272
rect 26615 -38592 26935 -38508
rect 26615 -38828 26657 -38592
rect 26893 -38828 26935 -38592
rect 26615 -38890 26935 -38828
rect 27615 -38272 27935 -38210
rect 27615 -38508 27657 -38272
rect 27893 -38508 27935 -38272
rect 27615 -38592 27935 -38508
rect 27615 -38828 27657 -38592
rect 27893 -38828 27935 -38592
rect 27615 -38890 27935 -38828
rect 28615 -38272 28935 -38210
rect 28615 -38508 28657 -38272
rect 28893 -38508 28935 -38272
rect 28615 -38592 28935 -38508
rect 28615 -38828 28657 -38592
rect 28893 -38828 28935 -38592
rect 28615 -38890 28935 -38828
rect 29615 -38272 29935 -38210
rect 29615 -38508 29657 -38272
rect 29893 -38508 29935 -38272
rect 29615 -38592 29935 -38508
rect 29615 -38828 29657 -38592
rect 29893 -38828 29935 -38592
rect 29615 -38890 29935 -38828
rect 30615 -38272 30935 -38210
rect 30615 -38508 30657 -38272
rect 30893 -38508 30935 -38272
rect 30615 -38592 30935 -38508
rect 30615 -38828 30657 -38592
rect 30893 -38828 30935 -38592
rect 30615 -38890 30935 -38828
rect 31615 -38272 31935 -38210
rect 31615 -38508 31657 -38272
rect 31893 -38508 31935 -38272
rect 31615 -38592 31935 -38508
rect 31615 -38828 31657 -38592
rect 31893 -38828 31935 -38592
rect 31615 -38890 31935 -38828
rect 32615 -38272 32935 -38210
rect 32615 -38508 32657 -38272
rect 32893 -38508 32935 -38272
rect 32615 -38592 32935 -38508
rect 32615 -38828 32657 -38592
rect 32893 -38828 32935 -38592
rect 32615 -38890 32935 -38828
rect 33615 -38272 33935 -38210
rect 33615 -38508 33657 -38272
rect 33893 -38508 33935 -38272
rect 33615 -38592 33935 -38508
rect 33615 -38828 33657 -38592
rect 33893 -38828 33935 -38592
rect 33615 -38890 33935 -38828
rect 8275 -38932 34275 -38890
rect 8275 -39168 8317 -38932
rect 8553 -39168 8657 -38932
rect 8893 -39168 8997 -38932
rect 9233 -39168 9317 -38932
rect 9553 -39168 9657 -38932
rect 9893 -39168 9997 -38932
rect 10233 -39168 10317 -38932
rect 10553 -39168 10657 -38932
rect 10893 -39168 10997 -38932
rect 11233 -39168 11317 -38932
rect 11553 -39168 11657 -38932
rect 11893 -39168 11997 -38932
rect 12233 -39168 12317 -38932
rect 12553 -39168 12657 -38932
rect 12893 -39168 12997 -38932
rect 13233 -39168 13317 -38932
rect 13553 -39168 13657 -38932
rect 13893 -39168 13997 -38932
rect 14233 -39168 14317 -38932
rect 14553 -39168 14657 -38932
rect 14893 -39168 14997 -38932
rect 15233 -39168 15317 -38932
rect 15553 -39168 15657 -38932
rect 15893 -39168 15997 -38932
rect 16233 -39168 16317 -38932
rect 16553 -39168 16657 -38932
rect 16893 -39168 16997 -38932
rect 17233 -39168 17317 -38932
rect 17553 -39168 17657 -38932
rect 17893 -39168 17997 -38932
rect 18233 -39168 18317 -38932
rect 18553 -39168 18657 -38932
rect 18893 -39168 18997 -38932
rect 19233 -39168 19317 -38932
rect 19553 -39168 19657 -38932
rect 19893 -39168 19997 -38932
rect 20233 -39168 20317 -38932
rect 20553 -39168 20657 -38932
rect 20893 -39168 20997 -38932
rect 21233 -39168 21317 -38932
rect 21553 -39168 21657 -38932
rect 21893 -39168 21997 -38932
rect 22233 -39168 22317 -38932
rect 22553 -39168 22657 -38932
rect 22893 -39168 22997 -38932
rect 23233 -39168 23317 -38932
rect 23553 -39168 23657 -38932
rect 23893 -39168 23997 -38932
rect 24233 -39168 24317 -38932
rect 24553 -39168 24657 -38932
rect 24893 -39168 24997 -38932
rect 25233 -39168 25317 -38932
rect 25553 -39168 25657 -38932
rect 25893 -39168 25997 -38932
rect 26233 -39168 26317 -38932
rect 26553 -39168 26657 -38932
rect 26893 -39168 26997 -38932
rect 27233 -39168 27317 -38932
rect 27553 -39168 27657 -38932
rect 27893 -39168 27997 -38932
rect 28233 -39168 28317 -38932
rect 28553 -39168 28657 -38932
rect 28893 -39168 28997 -38932
rect 29233 -39168 29317 -38932
rect 29553 -39168 29657 -38932
rect 29893 -39168 29997 -38932
rect 30233 -39168 30317 -38932
rect 30553 -39168 30657 -38932
rect 30893 -39168 30997 -38932
rect 31233 -39168 31317 -38932
rect 31553 -39168 31657 -38932
rect 31893 -39168 31997 -38932
rect 32233 -39168 32317 -38932
rect 32553 -39168 32657 -38932
rect 32893 -39168 32997 -38932
rect 33233 -39168 33317 -38932
rect 33553 -39168 33657 -38932
rect 33893 -39168 33997 -38932
rect 34233 -39168 34275 -38932
rect 8275 -39210 34275 -39168
rect 8615 -39272 8935 -39210
rect 8615 -39508 8657 -39272
rect 8893 -39508 8935 -39272
rect 8615 -39592 8935 -39508
rect 8615 -39828 8657 -39592
rect 8893 -39828 8935 -39592
rect 8615 -39890 8935 -39828
rect 9615 -39272 9935 -39210
rect 9615 -39508 9657 -39272
rect 9893 -39508 9935 -39272
rect 9615 -39592 9935 -39508
rect 9615 -39828 9657 -39592
rect 9893 -39828 9935 -39592
rect 9615 -39890 9935 -39828
rect 10615 -39272 10935 -39210
rect 10615 -39508 10657 -39272
rect 10893 -39508 10935 -39272
rect 10615 -39592 10935 -39508
rect 10615 -39828 10657 -39592
rect 10893 -39828 10935 -39592
rect 10615 -39890 10935 -39828
rect 11615 -39272 11935 -39210
rect 11615 -39508 11657 -39272
rect 11893 -39508 11935 -39272
rect 11615 -39592 11935 -39508
rect 11615 -39828 11657 -39592
rect 11893 -39828 11935 -39592
rect 11615 -39890 11935 -39828
rect 12615 -39272 12935 -39210
rect 12615 -39508 12657 -39272
rect 12893 -39508 12935 -39272
rect 12615 -39592 12935 -39508
rect 12615 -39828 12657 -39592
rect 12893 -39828 12935 -39592
rect 12615 -39890 12935 -39828
rect 13615 -39272 13935 -39210
rect 13615 -39508 13657 -39272
rect 13893 -39508 13935 -39272
rect 13615 -39592 13935 -39508
rect 13615 -39828 13657 -39592
rect 13893 -39828 13935 -39592
rect 13615 -39890 13935 -39828
rect 14615 -39272 14935 -39210
rect 14615 -39508 14657 -39272
rect 14893 -39508 14935 -39272
rect 14615 -39592 14935 -39508
rect 14615 -39828 14657 -39592
rect 14893 -39828 14935 -39592
rect 14615 -39890 14935 -39828
rect 15615 -39272 15935 -39210
rect 15615 -39508 15657 -39272
rect 15893 -39508 15935 -39272
rect 15615 -39592 15935 -39508
rect 15615 -39828 15657 -39592
rect 15893 -39828 15935 -39592
rect 15615 -39890 15935 -39828
rect 16615 -39272 16935 -39210
rect 16615 -39508 16657 -39272
rect 16893 -39508 16935 -39272
rect 16615 -39592 16935 -39508
rect 16615 -39828 16657 -39592
rect 16893 -39828 16935 -39592
rect 16615 -39890 16935 -39828
rect 17615 -39272 17935 -39210
rect 17615 -39508 17657 -39272
rect 17893 -39508 17935 -39272
rect 17615 -39592 17935 -39508
rect 17615 -39828 17657 -39592
rect 17893 -39828 17935 -39592
rect 17615 -39890 17935 -39828
rect 18615 -39272 18935 -39210
rect 18615 -39508 18657 -39272
rect 18893 -39508 18935 -39272
rect 18615 -39592 18935 -39508
rect 18615 -39828 18657 -39592
rect 18893 -39828 18935 -39592
rect 18615 -39890 18935 -39828
rect 19615 -39272 19935 -39210
rect 19615 -39508 19657 -39272
rect 19893 -39508 19935 -39272
rect 19615 -39592 19935 -39508
rect 19615 -39828 19657 -39592
rect 19893 -39828 19935 -39592
rect 19615 -39890 19935 -39828
rect 20615 -39272 20935 -39210
rect 20615 -39508 20657 -39272
rect 20893 -39508 20935 -39272
rect 20615 -39592 20935 -39508
rect 20615 -39828 20657 -39592
rect 20893 -39828 20935 -39592
rect 20615 -39890 20935 -39828
rect 21615 -39272 21935 -39210
rect 21615 -39508 21657 -39272
rect 21893 -39508 21935 -39272
rect 21615 -39592 21935 -39508
rect 21615 -39828 21657 -39592
rect 21893 -39828 21935 -39592
rect 21615 -39890 21935 -39828
rect 22615 -39272 22935 -39210
rect 22615 -39508 22657 -39272
rect 22893 -39508 22935 -39272
rect 22615 -39592 22935 -39508
rect 22615 -39828 22657 -39592
rect 22893 -39828 22935 -39592
rect 22615 -39890 22935 -39828
rect 23615 -39272 23935 -39210
rect 23615 -39508 23657 -39272
rect 23893 -39508 23935 -39272
rect 23615 -39592 23935 -39508
rect 23615 -39828 23657 -39592
rect 23893 -39828 23935 -39592
rect 23615 -39890 23935 -39828
rect 24615 -39272 24935 -39210
rect 24615 -39508 24657 -39272
rect 24893 -39508 24935 -39272
rect 24615 -39592 24935 -39508
rect 24615 -39828 24657 -39592
rect 24893 -39828 24935 -39592
rect 24615 -39890 24935 -39828
rect 25615 -39272 25935 -39210
rect 25615 -39508 25657 -39272
rect 25893 -39508 25935 -39272
rect 25615 -39592 25935 -39508
rect 25615 -39828 25657 -39592
rect 25893 -39828 25935 -39592
rect 25615 -39890 25935 -39828
rect 26615 -39272 26935 -39210
rect 26615 -39508 26657 -39272
rect 26893 -39508 26935 -39272
rect 26615 -39592 26935 -39508
rect 26615 -39828 26657 -39592
rect 26893 -39828 26935 -39592
rect 26615 -39890 26935 -39828
rect 27615 -39272 27935 -39210
rect 27615 -39508 27657 -39272
rect 27893 -39508 27935 -39272
rect 27615 -39592 27935 -39508
rect 27615 -39828 27657 -39592
rect 27893 -39828 27935 -39592
rect 27615 -39890 27935 -39828
rect 28615 -39272 28935 -39210
rect 28615 -39508 28657 -39272
rect 28893 -39508 28935 -39272
rect 28615 -39592 28935 -39508
rect 28615 -39828 28657 -39592
rect 28893 -39828 28935 -39592
rect 28615 -39890 28935 -39828
rect 29615 -39272 29935 -39210
rect 29615 -39508 29657 -39272
rect 29893 -39508 29935 -39272
rect 29615 -39592 29935 -39508
rect 29615 -39828 29657 -39592
rect 29893 -39828 29935 -39592
rect 29615 -39890 29935 -39828
rect 30615 -39272 30935 -39210
rect 30615 -39508 30657 -39272
rect 30893 -39508 30935 -39272
rect 30615 -39592 30935 -39508
rect 30615 -39828 30657 -39592
rect 30893 -39828 30935 -39592
rect 30615 -39890 30935 -39828
rect 31615 -39272 31935 -39210
rect 31615 -39508 31657 -39272
rect 31893 -39508 31935 -39272
rect 31615 -39592 31935 -39508
rect 31615 -39828 31657 -39592
rect 31893 -39828 31935 -39592
rect 31615 -39890 31935 -39828
rect 32615 -39272 32935 -39210
rect 32615 -39508 32657 -39272
rect 32893 -39508 32935 -39272
rect 32615 -39592 32935 -39508
rect 32615 -39828 32657 -39592
rect 32893 -39828 32935 -39592
rect 32615 -39890 32935 -39828
rect 33615 -39272 33935 -39210
rect 33615 -39508 33657 -39272
rect 33893 -39508 33935 -39272
rect 33615 -39592 33935 -39508
rect 33615 -39828 33657 -39592
rect 33893 -39828 33935 -39592
rect 33615 -39890 33935 -39828
rect 8275 -39932 34275 -39890
rect 8275 -40168 8317 -39932
rect 8553 -40168 8657 -39932
rect 8893 -40168 8997 -39932
rect 9233 -40168 9317 -39932
rect 9553 -40168 9657 -39932
rect 9893 -40168 9997 -39932
rect 10233 -40168 10317 -39932
rect 10553 -40168 10657 -39932
rect 10893 -40168 10997 -39932
rect 11233 -40168 11317 -39932
rect 11553 -40168 11657 -39932
rect 11893 -40168 11997 -39932
rect 12233 -40168 12317 -39932
rect 12553 -40168 12657 -39932
rect 12893 -40168 12997 -39932
rect 13233 -40168 13317 -39932
rect 13553 -40168 13657 -39932
rect 13893 -40168 13997 -39932
rect 14233 -40168 14317 -39932
rect 14553 -40168 14657 -39932
rect 14893 -40168 14997 -39932
rect 15233 -40168 15317 -39932
rect 15553 -40168 15657 -39932
rect 15893 -40168 15997 -39932
rect 16233 -40168 16317 -39932
rect 16553 -40168 16657 -39932
rect 16893 -40168 16997 -39932
rect 17233 -40168 17317 -39932
rect 17553 -40168 17657 -39932
rect 17893 -40168 17997 -39932
rect 18233 -40168 18317 -39932
rect 18553 -40168 18657 -39932
rect 18893 -40168 18997 -39932
rect 19233 -40168 19317 -39932
rect 19553 -40168 19657 -39932
rect 19893 -40168 19997 -39932
rect 20233 -40168 20317 -39932
rect 20553 -40168 20657 -39932
rect 20893 -40168 20997 -39932
rect 21233 -40168 21317 -39932
rect 21553 -40168 21657 -39932
rect 21893 -40168 21997 -39932
rect 22233 -40168 22317 -39932
rect 22553 -40168 22657 -39932
rect 22893 -40168 22997 -39932
rect 23233 -40168 23317 -39932
rect 23553 -40168 23657 -39932
rect 23893 -40168 23997 -39932
rect 24233 -40168 24317 -39932
rect 24553 -40168 24657 -39932
rect 24893 -40168 24997 -39932
rect 25233 -40168 25317 -39932
rect 25553 -40168 25657 -39932
rect 25893 -40168 25997 -39932
rect 26233 -40168 26317 -39932
rect 26553 -40168 26657 -39932
rect 26893 -40168 26997 -39932
rect 27233 -40168 27317 -39932
rect 27553 -40168 27657 -39932
rect 27893 -40168 27997 -39932
rect 28233 -40168 28317 -39932
rect 28553 -40168 28657 -39932
rect 28893 -40168 28997 -39932
rect 29233 -40168 29317 -39932
rect 29553 -40168 29657 -39932
rect 29893 -40168 29997 -39932
rect 30233 -40168 30317 -39932
rect 30553 -40168 30657 -39932
rect 30893 -40168 30997 -39932
rect 31233 -40168 31317 -39932
rect 31553 -40168 31657 -39932
rect 31893 -40168 31997 -39932
rect 32233 -40168 32317 -39932
rect 32553 -40168 32657 -39932
rect 32893 -40168 32997 -39932
rect 33233 -40168 33317 -39932
rect 33553 -40168 33657 -39932
rect 33893 -40168 33997 -39932
rect 34233 -40168 34275 -39932
rect 8275 -40210 34275 -40168
rect 8615 -40272 8935 -40210
rect 8615 -40508 8657 -40272
rect 8893 -40508 8935 -40272
rect 8615 -40592 8935 -40508
rect 8615 -40828 8657 -40592
rect 8893 -40828 8935 -40592
rect 8615 -40890 8935 -40828
rect 9615 -40272 9935 -40210
rect 9615 -40508 9657 -40272
rect 9893 -40508 9935 -40272
rect 9615 -40592 9935 -40508
rect 9615 -40828 9657 -40592
rect 9893 -40828 9935 -40592
rect 9615 -40890 9935 -40828
rect 10615 -40272 10935 -40210
rect 10615 -40508 10657 -40272
rect 10893 -40508 10935 -40272
rect 10615 -40592 10935 -40508
rect 10615 -40828 10657 -40592
rect 10893 -40828 10935 -40592
rect 10615 -40890 10935 -40828
rect 11615 -40272 11935 -40210
rect 11615 -40508 11657 -40272
rect 11893 -40508 11935 -40272
rect 11615 -40592 11935 -40508
rect 11615 -40828 11657 -40592
rect 11893 -40828 11935 -40592
rect 11615 -40890 11935 -40828
rect 12615 -40272 12935 -40210
rect 12615 -40508 12657 -40272
rect 12893 -40508 12935 -40272
rect 12615 -40592 12935 -40508
rect 12615 -40828 12657 -40592
rect 12893 -40828 12935 -40592
rect 12615 -40890 12935 -40828
rect 13615 -40272 13935 -40210
rect 13615 -40508 13657 -40272
rect 13893 -40508 13935 -40272
rect 13615 -40592 13935 -40508
rect 13615 -40828 13657 -40592
rect 13893 -40828 13935 -40592
rect 13615 -40890 13935 -40828
rect 14615 -40272 14935 -40210
rect 14615 -40508 14657 -40272
rect 14893 -40508 14935 -40272
rect 14615 -40592 14935 -40508
rect 14615 -40828 14657 -40592
rect 14893 -40828 14935 -40592
rect 14615 -40890 14935 -40828
rect 15615 -40272 15935 -40210
rect 15615 -40508 15657 -40272
rect 15893 -40508 15935 -40272
rect 15615 -40592 15935 -40508
rect 15615 -40828 15657 -40592
rect 15893 -40828 15935 -40592
rect 15615 -40890 15935 -40828
rect 16615 -40272 16935 -40210
rect 16615 -40508 16657 -40272
rect 16893 -40508 16935 -40272
rect 16615 -40592 16935 -40508
rect 16615 -40828 16657 -40592
rect 16893 -40828 16935 -40592
rect 16615 -40890 16935 -40828
rect 17615 -40272 17935 -40210
rect 17615 -40508 17657 -40272
rect 17893 -40508 17935 -40272
rect 17615 -40592 17935 -40508
rect 17615 -40828 17657 -40592
rect 17893 -40828 17935 -40592
rect 17615 -40890 17935 -40828
rect 18615 -40272 18935 -40210
rect 18615 -40508 18657 -40272
rect 18893 -40508 18935 -40272
rect 18615 -40592 18935 -40508
rect 18615 -40828 18657 -40592
rect 18893 -40828 18935 -40592
rect 18615 -40890 18935 -40828
rect 19615 -40272 19935 -40210
rect 19615 -40508 19657 -40272
rect 19893 -40508 19935 -40272
rect 19615 -40592 19935 -40508
rect 19615 -40828 19657 -40592
rect 19893 -40828 19935 -40592
rect 19615 -40890 19935 -40828
rect 20615 -40272 20935 -40210
rect 20615 -40508 20657 -40272
rect 20893 -40508 20935 -40272
rect 20615 -40592 20935 -40508
rect 20615 -40828 20657 -40592
rect 20893 -40828 20935 -40592
rect 20615 -40890 20935 -40828
rect 21615 -40272 21935 -40210
rect 21615 -40508 21657 -40272
rect 21893 -40508 21935 -40272
rect 21615 -40592 21935 -40508
rect 21615 -40828 21657 -40592
rect 21893 -40828 21935 -40592
rect 21615 -40890 21935 -40828
rect 22615 -40272 22935 -40210
rect 22615 -40508 22657 -40272
rect 22893 -40508 22935 -40272
rect 22615 -40592 22935 -40508
rect 22615 -40828 22657 -40592
rect 22893 -40828 22935 -40592
rect 22615 -40890 22935 -40828
rect 23615 -40272 23935 -40210
rect 23615 -40508 23657 -40272
rect 23893 -40508 23935 -40272
rect 23615 -40592 23935 -40508
rect 23615 -40828 23657 -40592
rect 23893 -40828 23935 -40592
rect 23615 -40890 23935 -40828
rect 24615 -40272 24935 -40210
rect 24615 -40508 24657 -40272
rect 24893 -40508 24935 -40272
rect 24615 -40592 24935 -40508
rect 24615 -40828 24657 -40592
rect 24893 -40828 24935 -40592
rect 24615 -40890 24935 -40828
rect 25615 -40272 25935 -40210
rect 25615 -40508 25657 -40272
rect 25893 -40508 25935 -40272
rect 25615 -40592 25935 -40508
rect 25615 -40828 25657 -40592
rect 25893 -40828 25935 -40592
rect 25615 -40890 25935 -40828
rect 26615 -40272 26935 -40210
rect 26615 -40508 26657 -40272
rect 26893 -40508 26935 -40272
rect 26615 -40592 26935 -40508
rect 26615 -40828 26657 -40592
rect 26893 -40828 26935 -40592
rect 26615 -40890 26935 -40828
rect 27615 -40272 27935 -40210
rect 27615 -40508 27657 -40272
rect 27893 -40508 27935 -40272
rect 27615 -40592 27935 -40508
rect 27615 -40828 27657 -40592
rect 27893 -40828 27935 -40592
rect 27615 -40890 27935 -40828
rect 28615 -40272 28935 -40210
rect 28615 -40508 28657 -40272
rect 28893 -40508 28935 -40272
rect 28615 -40592 28935 -40508
rect 28615 -40828 28657 -40592
rect 28893 -40828 28935 -40592
rect 28615 -40890 28935 -40828
rect 29615 -40272 29935 -40210
rect 29615 -40508 29657 -40272
rect 29893 -40508 29935 -40272
rect 29615 -40592 29935 -40508
rect 29615 -40828 29657 -40592
rect 29893 -40828 29935 -40592
rect 29615 -40890 29935 -40828
rect 30615 -40272 30935 -40210
rect 30615 -40508 30657 -40272
rect 30893 -40508 30935 -40272
rect 30615 -40592 30935 -40508
rect 30615 -40828 30657 -40592
rect 30893 -40828 30935 -40592
rect 30615 -40890 30935 -40828
rect 31615 -40272 31935 -40210
rect 31615 -40508 31657 -40272
rect 31893 -40508 31935 -40272
rect 31615 -40592 31935 -40508
rect 31615 -40828 31657 -40592
rect 31893 -40828 31935 -40592
rect 31615 -40890 31935 -40828
rect 32615 -40272 32935 -40210
rect 32615 -40508 32657 -40272
rect 32893 -40508 32935 -40272
rect 32615 -40592 32935 -40508
rect 32615 -40828 32657 -40592
rect 32893 -40828 32935 -40592
rect 32615 -40890 32935 -40828
rect 33615 -40272 33935 -40210
rect 33615 -40508 33657 -40272
rect 33893 -40508 33935 -40272
rect 33615 -40592 33935 -40508
rect 33615 -40828 33657 -40592
rect 33893 -40828 33935 -40592
rect 33615 -40890 33935 -40828
rect 8275 -40932 34275 -40890
rect 8275 -41168 8317 -40932
rect 8553 -41168 8657 -40932
rect 8893 -41168 8997 -40932
rect 9233 -41168 9317 -40932
rect 9553 -41168 9657 -40932
rect 9893 -41168 9997 -40932
rect 10233 -41168 10317 -40932
rect 10553 -41168 10657 -40932
rect 10893 -41168 10997 -40932
rect 11233 -41168 11317 -40932
rect 11553 -41168 11657 -40932
rect 11893 -41168 11997 -40932
rect 12233 -41168 12317 -40932
rect 12553 -41168 12657 -40932
rect 12893 -41168 12997 -40932
rect 13233 -41168 13317 -40932
rect 13553 -41168 13657 -40932
rect 13893 -41168 13997 -40932
rect 14233 -41168 14317 -40932
rect 14553 -41168 14657 -40932
rect 14893 -41168 14997 -40932
rect 15233 -41168 15317 -40932
rect 15553 -41168 15657 -40932
rect 15893 -41168 15997 -40932
rect 16233 -41168 16317 -40932
rect 16553 -41168 16657 -40932
rect 16893 -41168 16997 -40932
rect 17233 -41168 17317 -40932
rect 17553 -41168 17657 -40932
rect 17893 -41168 17997 -40932
rect 18233 -41168 18317 -40932
rect 18553 -41168 18657 -40932
rect 18893 -41168 18997 -40932
rect 19233 -41168 19317 -40932
rect 19553 -41168 19657 -40932
rect 19893 -41168 19997 -40932
rect 20233 -41168 20317 -40932
rect 20553 -41168 20657 -40932
rect 20893 -41168 20997 -40932
rect 21233 -41168 21317 -40932
rect 21553 -41168 21657 -40932
rect 21893 -41168 21997 -40932
rect 22233 -41168 22317 -40932
rect 22553 -41168 22657 -40932
rect 22893 -41168 22997 -40932
rect 23233 -41168 23317 -40932
rect 23553 -41168 23657 -40932
rect 23893 -41168 23997 -40932
rect 24233 -41168 24317 -40932
rect 24553 -41168 24657 -40932
rect 24893 -41168 24997 -40932
rect 25233 -41168 25317 -40932
rect 25553 -41168 25657 -40932
rect 25893 -41168 25997 -40932
rect 26233 -41168 26317 -40932
rect 26553 -41168 26657 -40932
rect 26893 -41168 26997 -40932
rect 27233 -41168 27317 -40932
rect 27553 -41168 27657 -40932
rect 27893 -41168 27997 -40932
rect 28233 -41168 28317 -40932
rect 28553 -41168 28657 -40932
rect 28893 -41168 28997 -40932
rect 29233 -41168 29317 -40932
rect 29553 -41168 29657 -40932
rect 29893 -41168 29997 -40932
rect 30233 -41168 30317 -40932
rect 30553 -41168 30657 -40932
rect 30893 -41168 30997 -40932
rect 31233 -41168 31317 -40932
rect 31553 -41168 31657 -40932
rect 31893 -41168 31997 -40932
rect 32233 -41168 32317 -40932
rect 32553 -41168 32657 -40932
rect 32893 -41168 32997 -40932
rect 33233 -41168 33317 -40932
rect 33553 -41168 33657 -40932
rect 33893 -41168 33997 -40932
rect 34233 -41168 34275 -40932
rect 8275 -41210 34275 -41168
rect 8615 -41272 8935 -41210
rect 8615 -41508 8657 -41272
rect 8893 -41508 8935 -41272
rect 8615 -41592 8935 -41508
rect 8615 -41828 8657 -41592
rect 8893 -41828 8935 -41592
rect 8615 -41890 8935 -41828
rect 9615 -41272 9935 -41210
rect 9615 -41508 9657 -41272
rect 9893 -41508 9935 -41272
rect 9615 -41592 9935 -41508
rect 9615 -41828 9657 -41592
rect 9893 -41828 9935 -41592
rect 9615 -41890 9935 -41828
rect 10615 -41272 10935 -41210
rect 10615 -41508 10657 -41272
rect 10893 -41508 10935 -41272
rect 10615 -41592 10935 -41508
rect 10615 -41828 10657 -41592
rect 10893 -41828 10935 -41592
rect 10615 -41890 10935 -41828
rect 11615 -41272 11935 -41210
rect 11615 -41508 11657 -41272
rect 11893 -41508 11935 -41272
rect 11615 -41592 11935 -41508
rect 11615 -41828 11657 -41592
rect 11893 -41828 11935 -41592
rect 11615 -41890 11935 -41828
rect 12615 -41272 12935 -41210
rect 12615 -41508 12657 -41272
rect 12893 -41508 12935 -41272
rect 12615 -41592 12935 -41508
rect 12615 -41828 12657 -41592
rect 12893 -41828 12935 -41592
rect 12615 -41890 12935 -41828
rect 13615 -41272 13935 -41210
rect 13615 -41508 13657 -41272
rect 13893 -41508 13935 -41272
rect 13615 -41592 13935 -41508
rect 13615 -41828 13657 -41592
rect 13893 -41828 13935 -41592
rect 13615 -41890 13935 -41828
rect 14615 -41272 14935 -41210
rect 14615 -41508 14657 -41272
rect 14893 -41508 14935 -41272
rect 14615 -41592 14935 -41508
rect 14615 -41828 14657 -41592
rect 14893 -41828 14935 -41592
rect 14615 -41890 14935 -41828
rect 15615 -41272 15935 -41210
rect 15615 -41508 15657 -41272
rect 15893 -41508 15935 -41272
rect 15615 -41592 15935 -41508
rect 15615 -41828 15657 -41592
rect 15893 -41828 15935 -41592
rect 15615 -41890 15935 -41828
rect 16615 -41272 16935 -41210
rect 16615 -41508 16657 -41272
rect 16893 -41508 16935 -41272
rect 16615 -41592 16935 -41508
rect 16615 -41828 16657 -41592
rect 16893 -41828 16935 -41592
rect 16615 -41890 16935 -41828
rect 17615 -41272 17935 -41210
rect 17615 -41508 17657 -41272
rect 17893 -41508 17935 -41272
rect 17615 -41592 17935 -41508
rect 17615 -41828 17657 -41592
rect 17893 -41828 17935 -41592
rect 17615 -41890 17935 -41828
rect 18615 -41272 18935 -41210
rect 18615 -41508 18657 -41272
rect 18893 -41508 18935 -41272
rect 18615 -41592 18935 -41508
rect 18615 -41828 18657 -41592
rect 18893 -41828 18935 -41592
rect 18615 -41890 18935 -41828
rect 19615 -41272 19935 -41210
rect 19615 -41508 19657 -41272
rect 19893 -41508 19935 -41272
rect 19615 -41592 19935 -41508
rect 19615 -41828 19657 -41592
rect 19893 -41828 19935 -41592
rect 19615 -41890 19935 -41828
rect 20615 -41272 20935 -41210
rect 20615 -41508 20657 -41272
rect 20893 -41508 20935 -41272
rect 20615 -41592 20935 -41508
rect 20615 -41828 20657 -41592
rect 20893 -41828 20935 -41592
rect 20615 -41890 20935 -41828
rect 21615 -41272 21935 -41210
rect 21615 -41508 21657 -41272
rect 21893 -41508 21935 -41272
rect 21615 -41592 21935 -41508
rect 21615 -41828 21657 -41592
rect 21893 -41828 21935 -41592
rect 21615 -41890 21935 -41828
rect 22615 -41272 22935 -41210
rect 22615 -41508 22657 -41272
rect 22893 -41508 22935 -41272
rect 22615 -41592 22935 -41508
rect 22615 -41828 22657 -41592
rect 22893 -41828 22935 -41592
rect 22615 -41890 22935 -41828
rect 23615 -41272 23935 -41210
rect 23615 -41508 23657 -41272
rect 23893 -41508 23935 -41272
rect 23615 -41592 23935 -41508
rect 23615 -41828 23657 -41592
rect 23893 -41828 23935 -41592
rect 23615 -41890 23935 -41828
rect 24615 -41272 24935 -41210
rect 24615 -41508 24657 -41272
rect 24893 -41508 24935 -41272
rect 24615 -41592 24935 -41508
rect 24615 -41828 24657 -41592
rect 24893 -41828 24935 -41592
rect 24615 -41890 24935 -41828
rect 25615 -41272 25935 -41210
rect 25615 -41508 25657 -41272
rect 25893 -41508 25935 -41272
rect 25615 -41592 25935 -41508
rect 25615 -41828 25657 -41592
rect 25893 -41828 25935 -41592
rect 25615 -41890 25935 -41828
rect 26615 -41272 26935 -41210
rect 26615 -41508 26657 -41272
rect 26893 -41508 26935 -41272
rect 26615 -41592 26935 -41508
rect 26615 -41828 26657 -41592
rect 26893 -41828 26935 -41592
rect 26615 -41890 26935 -41828
rect 27615 -41272 27935 -41210
rect 27615 -41508 27657 -41272
rect 27893 -41508 27935 -41272
rect 27615 -41592 27935 -41508
rect 27615 -41828 27657 -41592
rect 27893 -41828 27935 -41592
rect 27615 -41890 27935 -41828
rect 28615 -41272 28935 -41210
rect 28615 -41508 28657 -41272
rect 28893 -41508 28935 -41272
rect 28615 -41592 28935 -41508
rect 28615 -41828 28657 -41592
rect 28893 -41828 28935 -41592
rect 28615 -41890 28935 -41828
rect 29615 -41272 29935 -41210
rect 29615 -41508 29657 -41272
rect 29893 -41508 29935 -41272
rect 29615 -41592 29935 -41508
rect 29615 -41828 29657 -41592
rect 29893 -41828 29935 -41592
rect 29615 -41890 29935 -41828
rect 30615 -41272 30935 -41210
rect 30615 -41508 30657 -41272
rect 30893 -41508 30935 -41272
rect 30615 -41592 30935 -41508
rect 30615 -41828 30657 -41592
rect 30893 -41828 30935 -41592
rect 30615 -41890 30935 -41828
rect 31615 -41272 31935 -41210
rect 31615 -41508 31657 -41272
rect 31893 -41508 31935 -41272
rect 31615 -41592 31935 -41508
rect 31615 -41828 31657 -41592
rect 31893 -41828 31935 -41592
rect 31615 -41890 31935 -41828
rect 32615 -41272 32935 -41210
rect 32615 -41508 32657 -41272
rect 32893 -41508 32935 -41272
rect 32615 -41592 32935 -41508
rect 32615 -41828 32657 -41592
rect 32893 -41828 32935 -41592
rect 32615 -41890 32935 -41828
rect 33615 -41272 33935 -41210
rect 33615 -41508 33657 -41272
rect 33893 -41508 33935 -41272
rect 33615 -41592 33935 -41508
rect 33615 -41828 33657 -41592
rect 33893 -41828 33935 -41592
rect 33615 -41890 33935 -41828
rect 8275 -41932 34275 -41890
rect 8275 -42168 8317 -41932
rect 8553 -42168 8657 -41932
rect 8893 -42168 8997 -41932
rect 9233 -42168 9317 -41932
rect 9553 -42168 9657 -41932
rect 9893 -42168 9997 -41932
rect 10233 -42168 10317 -41932
rect 10553 -42168 10657 -41932
rect 10893 -42168 10997 -41932
rect 11233 -42168 11317 -41932
rect 11553 -42168 11657 -41932
rect 11893 -42168 11997 -41932
rect 12233 -42168 12317 -41932
rect 12553 -42168 12657 -41932
rect 12893 -42168 12997 -41932
rect 13233 -42168 13317 -41932
rect 13553 -42168 13657 -41932
rect 13893 -42168 13997 -41932
rect 14233 -42168 14317 -41932
rect 14553 -42168 14657 -41932
rect 14893 -42168 14997 -41932
rect 15233 -42168 15317 -41932
rect 15553 -42168 15657 -41932
rect 15893 -42168 15997 -41932
rect 16233 -42168 16317 -41932
rect 16553 -42168 16657 -41932
rect 16893 -42168 16997 -41932
rect 17233 -42168 17317 -41932
rect 17553 -42168 17657 -41932
rect 17893 -42168 17997 -41932
rect 18233 -42168 18317 -41932
rect 18553 -42168 18657 -41932
rect 18893 -42168 18997 -41932
rect 19233 -42168 19317 -41932
rect 19553 -42168 19657 -41932
rect 19893 -42168 19997 -41932
rect 20233 -42168 20317 -41932
rect 20553 -42168 20657 -41932
rect 20893 -42168 20997 -41932
rect 21233 -42168 21317 -41932
rect 21553 -42168 21657 -41932
rect 21893 -42168 21997 -41932
rect 22233 -42168 22317 -41932
rect 22553 -42168 22657 -41932
rect 22893 -42168 22997 -41932
rect 23233 -42168 23317 -41932
rect 23553 -42168 23657 -41932
rect 23893 -42168 23997 -41932
rect 24233 -42168 24317 -41932
rect 24553 -42168 24657 -41932
rect 24893 -42168 24997 -41932
rect 25233 -42168 25317 -41932
rect 25553 -42168 25657 -41932
rect 25893 -42168 25997 -41932
rect 26233 -42168 26317 -41932
rect 26553 -42168 26657 -41932
rect 26893 -42168 26997 -41932
rect 27233 -42168 27317 -41932
rect 27553 -42168 27657 -41932
rect 27893 -42168 27997 -41932
rect 28233 -42168 28317 -41932
rect 28553 -42168 28657 -41932
rect 28893 -42168 28997 -41932
rect 29233 -42168 29317 -41932
rect 29553 -42168 29657 -41932
rect 29893 -42168 29997 -41932
rect 30233 -42168 30317 -41932
rect 30553 -42168 30657 -41932
rect 30893 -42168 30997 -41932
rect 31233 -42168 31317 -41932
rect 31553 -42168 31657 -41932
rect 31893 -42168 31997 -41932
rect 32233 -42168 32317 -41932
rect 32553 -42168 32657 -41932
rect 32893 -42168 32997 -41932
rect 33233 -42168 33317 -41932
rect 33553 -42168 33657 -41932
rect 33893 -42168 33997 -41932
rect 34233 -42168 34275 -41932
rect 8275 -42210 34275 -42168
rect 8615 -42272 8935 -42210
rect 8615 -42508 8657 -42272
rect 8893 -42508 8935 -42272
rect 8615 -42592 8935 -42508
rect 8615 -42828 8657 -42592
rect 8893 -42828 8935 -42592
rect 8615 -42890 8935 -42828
rect 9615 -42272 9935 -42210
rect 9615 -42508 9657 -42272
rect 9893 -42508 9935 -42272
rect 9615 -42592 9935 -42508
rect 9615 -42828 9657 -42592
rect 9893 -42828 9935 -42592
rect 9615 -42890 9935 -42828
rect 10615 -42272 10935 -42210
rect 10615 -42508 10657 -42272
rect 10893 -42508 10935 -42272
rect 10615 -42592 10935 -42508
rect 10615 -42828 10657 -42592
rect 10893 -42828 10935 -42592
rect 10615 -42890 10935 -42828
rect 11615 -42272 11935 -42210
rect 11615 -42508 11657 -42272
rect 11893 -42508 11935 -42272
rect 11615 -42592 11935 -42508
rect 11615 -42828 11657 -42592
rect 11893 -42828 11935 -42592
rect 11615 -42890 11935 -42828
rect 12615 -42272 12935 -42210
rect 12615 -42508 12657 -42272
rect 12893 -42508 12935 -42272
rect 12615 -42592 12935 -42508
rect 12615 -42828 12657 -42592
rect 12893 -42828 12935 -42592
rect 12615 -42890 12935 -42828
rect 13615 -42272 13935 -42210
rect 13615 -42508 13657 -42272
rect 13893 -42508 13935 -42272
rect 13615 -42592 13935 -42508
rect 13615 -42828 13657 -42592
rect 13893 -42828 13935 -42592
rect 13615 -42890 13935 -42828
rect 14615 -42272 14935 -42210
rect 14615 -42508 14657 -42272
rect 14893 -42508 14935 -42272
rect 14615 -42592 14935 -42508
rect 14615 -42828 14657 -42592
rect 14893 -42828 14935 -42592
rect 14615 -42890 14935 -42828
rect 15615 -42272 15935 -42210
rect 15615 -42508 15657 -42272
rect 15893 -42508 15935 -42272
rect 15615 -42592 15935 -42508
rect 15615 -42828 15657 -42592
rect 15893 -42828 15935 -42592
rect 15615 -42890 15935 -42828
rect 16615 -42272 16935 -42210
rect 16615 -42508 16657 -42272
rect 16893 -42508 16935 -42272
rect 16615 -42592 16935 -42508
rect 16615 -42828 16657 -42592
rect 16893 -42828 16935 -42592
rect 16615 -42890 16935 -42828
rect 17615 -42272 17935 -42210
rect 17615 -42508 17657 -42272
rect 17893 -42508 17935 -42272
rect 17615 -42592 17935 -42508
rect 17615 -42828 17657 -42592
rect 17893 -42828 17935 -42592
rect 17615 -42890 17935 -42828
rect 18615 -42272 18935 -42210
rect 18615 -42508 18657 -42272
rect 18893 -42508 18935 -42272
rect 18615 -42592 18935 -42508
rect 18615 -42828 18657 -42592
rect 18893 -42828 18935 -42592
rect 18615 -42890 18935 -42828
rect 19615 -42272 19935 -42210
rect 19615 -42508 19657 -42272
rect 19893 -42508 19935 -42272
rect 19615 -42592 19935 -42508
rect 19615 -42828 19657 -42592
rect 19893 -42828 19935 -42592
rect 19615 -42890 19935 -42828
rect 20615 -42272 20935 -42210
rect 20615 -42508 20657 -42272
rect 20893 -42508 20935 -42272
rect 20615 -42592 20935 -42508
rect 20615 -42828 20657 -42592
rect 20893 -42828 20935 -42592
rect 20615 -42890 20935 -42828
rect 21615 -42272 21935 -42210
rect 21615 -42508 21657 -42272
rect 21893 -42508 21935 -42272
rect 21615 -42592 21935 -42508
rect 21615 -42828 21657 -42592
rect 21893 -42828 21935 -42592
rect 21615 -42890 21935 -42828
rect 22615 -42272 22935 -42210
rect 22615 -42508 22657 -42272
rect 22893 -42508 22935 -42272
rect 22615 -42592 22935 -42508
rect 22615 -42828 22657 -42592
rect 22893 -42828 22935 -42592
rect 22615 -42890 22935 -42828
rect 23615 -42272 23935 -42210
rect 23615 -42508 23657 -42272
rect 23893 -42508 23935 -42272
rect 23615 -42592 23935 -42508
rect 23615 -42828 23657 -42592
rect 23893 -42828 23935 -42592
rect 23615 -42890 23935 -42828
rect 24615 -42272 24935 -42210
rect 24615 -42508 24657 -42272
rect 24893 -42508 24935 -42272
rect 24615 -42592 24935 -42508
rect 24615 -42828 24657 -42592
rect 24893 -42828 24935 -42592
rect 24615 -42890 24935 -42828
rect 25615 -42272 25935 -42210
rect 25615 -42508 25657 -42272
rect 25893 -42508 25935 -42272
rect 25615 -42592 25935 -42508
rect 25615 -42828 25657 -42592
rect 25893 -42828 25935 -42592
rect 25615 -42890 25935 -42828
rect 26615 -42272 26935 -42210
rect 26615 -42508 26657 -42272
rect 26893 -42508 26935 -42272
rect 26615 -42592 26935 -42508
rect 26615 -42828 26657 -42592
rect 26893 -42828 26935 -42592
rect 26615 -42890 26935 -42828
rect 27615 -42272 27935 -42210
rect 27615 -42508 27657 -42272
rect 27893 -42508 27935 -42272
rect 27615 -42592 27935 -42508
rect 27615 -42828 27657 -42592
rect 27893 -42828 27935 -42592
rect 27615 -42890 27935 -42828
rect 28615 -42272 28935 -42210
rect 28615 -42508 28657 -42272
rect 28893 -42508 28935 -42272
rect 28615 -42592 28935 -42508
rect 28615 -42828 28657 -42592
rect 28893 -42828 28935 -42592
rect 28615 -42890 28935 -42828
rect 29615 -42272 29935 -42210
rect 29615 -42508 29657 -42272
rect 29893 -42508 29935 -42272
rect 29615 -42592 29935 -42508
rect 29615 -42828 29657 -42592
rect 29893 -42828 29935 -42592
rect 29615 -42890 29935 -42828
rect 30615 -42272 30935 -42210
rect 30615 -42508 30657 -42272
rect 30893 -42508 30935 -42272
rect 30615 -42592 30935 -42508
rect 30615 -42828 30657 -42592
rect 30893 -42828 30935 -42592
rect 30615 -42890 30935 -42828
rect 31615 -42272 31935 -42210
rect 31615 -42508 31657 -42272
rect 31893 -42508 31935 -42272
rect 31615 -42592 31935 -42508
rect 31615 -42828 31657 -42592
rect 31893 -42828 31935 -42592
rect 31615 -42890 31935 -42828
rect 32615 -42272 32935 -42210
rect 32615 -42508 32657 -42272
rect 32893 -42508 32935 -42272
rect 32615 -42592 32935 -42508
rect 32615 -42828 32657 -42592
rect 32893 -42828 32935 -42592
rect 32615 -42890 32935 -42828
rect 33615 -42272 33935 -42210
rect 33615 -42508 33657 -42272
rect 33893 -42508 33935 -42272
rect 33615 -42592 33935 -42508
rect 33615 -42828 33657 -42592
rect 33893 -42828 33935 -42592
rect 33615 -42890 33935 -42828
rect 8275 -42932 34275 -42890
rect 8275 -43168 8317 -42932
rect 8553 -43168 8657 -42932
rect 8893 -43168 8997 -42932
rect 9233 -43168 9317 -42932
rect 9553 -43168 9657 -42932
rect 9893 -43168 9997 -42932
rect 10233 -43168 10317 -42932
rect 10553 -43168 10657 -42932
rect 10893 -43168 10997 -42932
rect 11233 -43168 11317 -42932
rect 11553 -43168 11657 -42932
rect 11893 -43168 11997 -42932
rect 12233 -43168 12317 -42932
rect 12553 -43168 12657 -42932
rect 12893 -43168 12997 -42932
rect 13233 -43168 13317 -42932
rect 13553 -43168 13657 -42932
rect 13893 -43168 13997 -42932
rect 14233 -43168 14317 -42932
rect 14553 -43168 14657 -42932
rect 14893 -43168 14997 -42932
rect 15233 -43168 15317 -42932
rect 15553 -43168 15657 -42932
rect 15893 -43168 15997 -42932
rect 16233 -43168 16317 -42932
rect 16553 -43168 16657 -42932
rect 16893 -43168 16997 -42932
rect 17233 -43168 17317 -42932
rect 17553 -43168 17657 -42932
rect 17893 -43168 17997 -42932
rect 18233 -43168 18317 -42932
rect 18553 -43168 18657 -42932
rect 18893 -43168 18997 -42932
rect 19233 -43168 19317 -42932
rect 19553 -43168 19657 -42932
rect 19893 -43168 19997 -42932
rect 20233 -43168 20317 -42932
rect 20553 -43168 20657 -42932
rect 20893 -43168 20997 -42932
rect 21233 -43168 21317 -42932
rect 21553 -43168 21657 -42932
rect 21893 -43168 21997 -42932
rect 22233 -43168 22317 -42932
rect 22553 -43168 22657 -42932
rect 22893 -43168 22997 -42932
rect 23233 -43168 23317 -42932
rect 23553 -43168 23657 -42932
rect 23893 -43168 23997 -42932
rect 24233 -43168 24317 -42932
rect 24553 -43168 24657 -42932
rect 24893 -43168 24997 -42932
rect 25233 -43168 25317 -42932
rect 25553 -43168 25657 -42932
rect 25893 -43168 25997 -42932
rect 26233 -43168 26317 -42932
rect 26553 -43168 26657 -42932
rect 26893 -43168 26997 -42932
rect 27233 -43168 27317 -42932
rect 27553 -43168 27657 -42932
rect 27893 -43168 27997 -42932
rect 28233 -43168 28317 -42932
rect 28553 -43168 28657 -42932
rect 28893 -43168 28997 -42932
rect 29233 -43168 29317 -42932
rect 29553 -43168 29657 -42932
rect 29893 -43168 29997 -42932
rect 30233 -43168 30317 -42932
rect 30553 -43168 30657 -42932
rect 30893 -43168 30997 -42932
rect 31233 -43168 31317 -42932
rect 31553 -43168 31657 -42932
rect 31893 -43168 31997 -42932
rect 32233 -43168 32317 -42932
rect 32553 -43168 32657 -42932
rect 32893 -43168 32997 -42932
rect 33233 -43168 33317 -42932
rect 33553 -43168 33657 -42932
rect 33893 -43168 33997 -42932
rect 34233 -43168 34275 -42932
rect 8275 -43210 34275 -43168
rect 8615 -43272 8935 -43210
rect 8615 -43508 8657 -43272
rect 8893 -43508 8935 -43272
rect 8615 -43592 8935 -43508
rect 8615 -43828 8657 -43592
rect 8893 -43828 8935 -43592
rect 8615 -43890 8935 -43828
rect 9615 -43272 9935 -43210
rect 9615 -43508 9657 -43272
rect 9893 -43508 9935 -43272
rect 9615 -43592 9935 -43508
rect 9615 -43828 9657 -43592
rect 9893 -43828 9935 -43592
rect 9615 -43890 9935 -43828
rect 10615 -43272 10935 -43210
rect 10615 -43508 10657 -43272
rect 10893 -43508 10935 -43272
rect 10615 -43592 10935 -43508
rect 10615 -43828 10657 -43592
rect 10893 -43828 10935 -43592
rect 10615 -43890 10935 -43828
rect 11615 -43272 11935 -43210
rect 11615 -43508 11657 -43272
rect 11893 -43508 11935 -43272
rect 11615 -43592 11935 -43508
rect 11615 -43828 11657 -43592
rect 11893 -43828 11935 -43592
rect 11615 -43890 11935 -43828
rect 12615 -43272 12935 -43210
rect 12615 -43508 12657 -43272
rect 12893 -43508 12935 -43272
rect 12615 -43592 12935 -43508
rect 12615 -43828 12657 -43592
rect 12893 -43828 12935 -43592
rect 12615 -43890 12935 -43828
rect 13615 -43272 13935 -43210
rect 13615 -43508 13657 -43272
rect 13893 -43508 13935 -43272
rect 13615 -43592 13935 -43508
rect 13615 -43828 13657 -43592
rect 13893 -43828 13935 -43592
rect 13615 -43890 13935 -43828
rect 14615 -43272 14935 -43210
rect 14615 -43508 14657 -43272
rect 14893 -43508 14935 -43272
rect 14615 -43592 14935 -43508
rect 14615 -43828 14657 -43592
rect 14893 -43828 14935 -43592
rect 14615 -43890 14935 -43828
rect 15615 -43272 15935 -43210
rect 15615 -43508 15657 -43272
rect 15893 -43508 15935 -43272
rect 15615 -43592 15935 -43508
rect 15615 -43828 15657 -43592
rect 15893 -43828 15935 -43592
rect 15615 -43890 15935 -43828
rect 16615 -43272 16935 -43210
rect 16615 -43508 16657 -43272
rect 16893 -43508 16935 -43272
rect 16615 -43592 16935 -43508
rect 16615 -43828 16657 -43592
rect 16893 -43828 16935 -43592
rect 16615 -43890 16935 -43828
rect 17615 -43272 17935 -43210
rect 17615 -43508 17657 -43272
rect 17893 -43508 17935 -43272
rect 17615 -43592 17935 -43508
rect 17615 -43828 17657 -43592
rect 17893 -43828 17935 -43592
rect 17615 -43890 17935 -43828
rect 18615 -43272 18935 -43210
rect 18615 -43508 18657 -43272
rect 18893 -43508 18935 -43272
rect 18615 -43592 18935 -43508
rect 18615 -43828 18657 -43592
rect 18893 -43828 18935 -43592
rect 18615 -43890 18935 -43828
rect 19615 -43272 19935 -43210
rect 19615 -43508 19657 -43272
rect 19893 -43508 19935 -43272
rect 19615 -43592 19935 -43508
rect 19615 -43828 19657 -43592
rect 19893 -43828 19935 -43592
rect 19615 -43890 19935 -43828
rect 20615 -43272 20935 -43210
rect 20615 -43508 20657 -43272
rect 20893 -43508 20935 -43272
rect 20615 -43592 20935 -43508
rect 20615 -43828 20657 -43592
rect 20893 -43828 20935 -43592
rect 20615 -43890 20935 -43828
rect 21615 -43272 21935 -43210
rect 21615 -43508 21657 -43272
rect 21893 -43508 21935 -43272
rect 21615 -43592 21935 -43508
rect 21615 -43828 21657 -43592
rect 21893 -43828 21935 -43592
rect 21615 -43890 21935 -43828
rect 22615 -43272 22935 -43210
rect 22615 -43508 22657 -43272
rect 22893 -43508 22935 -43272
rect 22615 -43592 22935 -43508
rect 22615 -43828 22657 -43592
rect 22893 -43828 22935 -43592
rect 22615 -43890 22935 -43828
rect 23615 -43272 23935 -43210
rect 23615 -43508 23657 -43272
rect 23893 -43508 23935 -43272
rect 23615 -43592 23935 -43508
rect 23615 -43828 23657 -43592
rect 23893 -43828 23935 -43592
rect 23615 -43890 23935 -43828
rect 24615 -43272 24935 -43210
rect 24615 -43508 24657 -43272
rect 24893 -43508 24935 -43272
rect 24615 -43592 24935 -43508
rect 24615 -43828 24657 -43592
rect 24893 -43828 24935 -43592
rect 24615 -43890 24935 -43828
rect 25615 -43272 25935 -43210
rect 25615 -43508 25657 -43272
rect 25893 -43508 25935 -43272
rect 25615 -43592 25935 -43508
rect 25615 -43828 25657 -43592
rect 25893 -43828 25935 -43592
rect 25615 -43890 25935 -43828
rect 26615 -43272 26935 -43210
rect 26615 -43508 26657 -43272
rect 26893 -43508 26935 -43272
rect 26615 -43592 26935 -43508
rect 26615 -43828 26657 -43592
rect 26893 -43828 26935 -43592
rect 26615 -43890 26935 -43828
rect 27615 -43272 27935 -43210
rect 27615 -43508 27657 -43272
rect 27893 -43508 27935 -43272
rect 27615 -43592 27935 -43508
rect 27615 -43828 27657 -43592
rect 27893 -43828 27935 -43592
rect 27615 -43890 27935 -43828
rect 28615 -43272 28935 -43210
rect 28615 -43508 28657 -43272
rect 28893 -43508 28935 -43272
rect 28615 -43592 28935 -43508
rect 28615 -43828 28657 -43592
rect 28893 -43828 28935 -43592
rect 28615 -43890 28935 -43828
rect 29615 -43272 29935 -43210
rect 29615 -43508 29657 -43272
rect 29893 -43508 29935 -43272
rect 29615 -43592 29935 -43508
rect 29615 -43828 29657 -43592
rect 29893 -43828 29935 -43592
rect 29615 -43890 29935 -43828
rect 30615 -43272 30935 -43210
rect 30615 -43508 30657 -43272
rect 30893 -43508 30935 -43272
rect 30615 -43592 30935 -43508
rect 30615 -43828 30657 -43592
rect 30893 -43828 30935 -43592
rect 30615 -43890 30935 -43828
rect 31615 -43272 31935 -43210
rect 31615 -43508 31657 -43272
rect 31893 -43508 31935 -43272
rect 31615 -43592 31935 -43508
rect 31615 -43828 31657 -43592
rect 31893 -43828 31935 -43592
rect 31615 -43890 31935 -43828
rect 32615 -43272 32935 -43210
rect 32615 -43508 32657 -43272
rect 32893 -43508 32935 -43272
rect 32615 -43592 32935 -43508
rect 32615 -43828 32657 -43592
rect 32893 -43828 32935 -43592
rect 32615 -43890 32935 -43828
rect 33615 -43272 33935 -43210
rect 33615 -43508 33657 -43272
rect 33893 -43508 33935 -43272
rect 33615 -43592 33935 -43508
rect 33615 -43828 33657 -43592
rect 33893 -43828 33935 -43592
rect 33615 -43890 33935 -43828
rect 8275 -43932 34275 -43890
rect 8275 -44168 8317 -43932
rect 8553 -44168 8657 -43932
rect 8893 -44168 8997 -43932
rect 9233 -44168 9317 -43932
rect 9553 -44168 9657 -43932
rect 9893 -44168 9997 -43932
rect 10233 -44168 10317 -43932
rect 10553 -44168 10657 -43932
rect 10893 -44168 10997 -43932
rect 11233 -44168 11317 -43932
rect 11553 -44168 11657 -43932
rect 11893 -44168 11997 -43932
rect 12233 -44168 12317 -43932
rect 12553 -44168 12657 -43932
rect 12893 -44168 12997 -43932
rect 13233 -44168 13317 -43932
rect 13553 -44168 13657 -43932
rect 13893 -44168 13997 -43932
rect 14233 -44168 14317 -43932
rect 14553 -44168 14657 -43932
rect 14893 -44168 14997 -43932
rect 15233 -44168 15317 -43932
rect 15553 -44168 15657 -43932
rect 15893 -44168 15997 -43932
rect 16233 -44168 16317 -43932
rect 16553 -44168 16657 -43932
rect 16893 -44168 16997 -43932
rect 17233 -44168 17317 -43932
rect 17553 -44168 17657 -43932
rect 17893 -44168 17997 -43932
rect 18233 -44168 18317 -43932
rect 18553 -44168 18657 -43932
rect 18893 -44168 18997 -43932
rect 19233 -44168 19317 -43932
rect 19553 -44168 19657 -43932
rect 19893 -44168 19997 -43932
rect 20233 -44168 20317 -43932
rect 20553 -44168 20657 -43932
rect 20893 -44168 20997 -43932
rect 21233 -44168 21317 -43932
rect 21553 -44168 21657 -43932
rect 21893 -44168 21997 -43932
rect 22233 -44168 22317 -43932
rect 22553 -44168 22657 -43932
rect 22893 -44168 22997 -43932
rect 23233 -44168 23317 -43932
rect 23553 -44168 23657 -43932
rect 23893 -44168 23997 -43932
rect 24233 -44168 24317 -43932
rect 24553 -44168 24657 -43932
rect 24893 -44168 24997 -43932
rect 25233 -44168 25317 -43932
rect 25553 -44168 25657 -43932
rect 25893 -44168 25997 -43932
rect 26233 -44168 26317 -43932
rect 26553 -44168 26657 -43932
rect 26893 -44168 26997 -43932
rect 27233 -44168 27317 -43932
rect 27553 -44168 27657 -43932
rect 27893 -44168 27997 -43932
rect 28233 -44168 28317 -43932
rect 28553 -44168 28657 -43932
rect 28893 -44168 28997 -43932
rect 29233 -44168 29317 -43932
rect 29553 -44168 29657 -43932
rect 29893 -44168 29997 -43932
rect 30233 -44168 30317 -43932
rect 30553 -44168 30657 -43932
rect 30893 -44168 30997 -43932
rect 31233 -44168 31317 -43932
rect 31553 -44168 31657 -43932
rect 31893 -44168 31997 -43932
rect 32233 -44168 32317 -43932
rect 32553 -44168 32657 -43932
rect 32893 -44168 32997 -43932
rect 33233 -44168 33317 -43932
rect 33553 -44168 33657 -43932
rect 33893 -44168 33997 -43932
rect 34233 -44168 34275 -43932
rect 8275 -44210 34275 -44168
tri -22905 -44550 -22875 -44520 ne
rect -22875 -44550 -17675 -44520
tri -17675 -44550 -17645 -44520 nw
rect -4275 -44550 5725 -44428
rect 8615 -44272 8935 -44210
rect 8615 -44508 8657 -44272
rect 8893 -44508 8935 -44272
rect -49485 -44828 -49443 -44592
rect -49207 -44828 -49165 -44592
rect -49485 -44890 -49165 -44828
rect 8615 -44592 8935 -44508
rect 8615 -44828 8657 -44592
rect 8893 -44828 8935 -44592
rect 8615 -44890 8935 -44828
rect 9615 -44272 9935 -44210
rect 9615 -44508 9657 -44272
rect 9893 -44508 9935 -44272
rect 9615 -44592 9935 -44508
rect 9615 -44828 9657 -44592
rect 9893 -44828 9935 -44592
rect 9615 -44890 9935 -44828
rect 10615 -44272 10935 -44210
rect 10615 -44508 10657 -44272
rect 10893 -44508 10935 -44272
rect 10615 -44592 10935 -44508
rect 10615 -44828 10657 -44592
rect 10893 -44828 10935 -44592
rect 10615 -44890 10935 -44828
rect 11615 -44272 11935 -44210
rect 11615 -44508 11657 -44272
rect 11893 -44508 11935 -44272
rect 11615 -44592 11935 -44508
rect 11615 -44828 11657 -44592
rect 11893 -44828 11935 -44592
rect 11615 -44890 11935 -44828
rect 12615 -44272 12935 -44210
rect 12615 -44508 12657 -44272
rect 12893 -44508 12935 -44272
rect 12615 -44592 12935 -44508
rect 12615 -44828 12657 -44592
rect 12893 -44828 12935 -44592
rect 12615 -44890 12935 -44828
rect 13615 -44272 13935 -44210
rect 13615 -44508 13657 -44272
rect 13893 -44508 13935 -44272
rect 13615 -44592 13935 -44508
rect 13615 -44828 13657 -44592
rect 13893 -44828 13935 -44592
rect 13615 -44890 13935 -44828
rect 14615 -44272 14935 -44210
rect 14615 -44508 14657 -44272
rect 14893 -44508 14935 -44272
rect 14615 -44592 14935 -44508
rect 14615 -44828 14657 -44592
rect 14893 -44828 14935 -44592
rect 14615 -44890 14935 -44828
rect 15615 -44272 15935 -44210
rect 15615 -44508 15657 -44272
rect 15893 -44508 15935 -44272
rect 15615 -44592 15935 -44508
rect 15615 -44828 15657 -44592
rect 15893 -44828 15935 -44592
rect 15615 -44890 15935 -44828
rect 16615 -44272 16935 -44210
rect 16615 -44508 16657 -44272
rect 16893 -44508 16935 -44272
rect 16615 -44592 16935 -44508
rect 16615 -44828 16657 -44592
rect 16893 -44828 16935 -44592
rect 16615 -44890 16935 -44828
rect 17615 -44272 17935 -44210
rect 17615 -44508 17657 -44272
rect 17893 -44508 17935 -44272
rect 17615 -44592 17935 -44508
rect 17615 -44828 17657 -44592
rect 17893 -44828 17935 -44592
rect 17615 -44890 17935 -44828
rect 18615 -44272 18935 -44210
rect 18615 -44508 18657 -44272
rect 18893 -44508 18935 -44272
rect 18615 -44592 18935 -44508
rect 18615 -44828 18657 -44592
rect 18893 -44828 18935 -44592
rect 18615 -44890 18935 -44828
rect 19615 -44272 19935 -44210
rect 19615 -44508 19657 -44272
rect 19893 -44508 19935 -44272
rect 19615 -44592 19935 -44508
rect 19615 -44828 19657 -44592
rect 19893 -44828 19935 -44592
rect 19615 -44890 19935 -44828
rect 20615 -44272 20935 -44210
rect 20615 -44508 20657 -44272
rect 20893 -44508 20935 -44272
rect 20615 -44592 20935 -44508
rect 20615 -44828 20657 -44592
rect 20893 -44828 20935 -44592
rect 20615 -44890 20935 -44828
rect 21615 -44272 21935 -44210
rect 21615 -44508 21657 -44272
rect 21893 -44508 21935 -44272
rect 21615 -44592 21935 -44508
rect 21615 -44828 21657 -44592
rect 21893 -44828 21935 -44592
rect 21615 -44890 21935 -44828
rect 22615 -44272 22935 -44210
rect 22615 -44508 22657 -44272
rect 22893 -44508 22935 -44272
rect 22615 -44592 22935 -44508
rect 22615 -44828 22657 -44592
rect 22893 -44828 22935 -44592
rect 22615 -44890 22935 -44828
rect 23615 -44272 23935 -44210
rect 23615 -44508 23657 -44272
rect 23893 -44508 23935 -44272
rect 23615 -44592 23935 -44508
rect 23615 -44828 23657 -44592
rect 23893 -44828 23935 -44592
rect 23615 -44890 23935 -44828
rect 24615 -44272 24935 -44210
rect 24615 -44508 24657 -44272
rect 24893 -44508 24935 -44272
rect 24615 -44592 24935 -44508
rect 24615 -44828 24657 -44592
rect 24893 -44828 24935 -44592
rect 24615 -44890 24935 -44828
rect 25615 -44272 25935 -44210
rect 25615 -44508 25657 -44272
rect 25893 -44508 25935 -44272
rect 25615 -44592 25935 -44508
rect 25615 -44828 25657 -44592
rect 25893 -44828 25935 -44592
rect 25615 -44890 25935 -44828
rect 26615 -44272 26935 -44210
rect 26615 -44508 26657 -44272
rect 26893 -44508 26935 -44272
rect 26615 -44592 26935 -44508
rect 26615 -44828 26657 -44592
rect 26893 -44828 26935 -44592
rect 26615 -44890 26935 -44828
rect 27615 -44272 27935 -44210
rect 27615 -44508 27657 -44272
rect 27893 -44508 27935 -44272
rect 27615 -44592 27935 -44508
rect 27615 -44828 27657 -44592
rect 27893 -44828 27935 -44592
rect 27615 -44890 27935 -44828
rect 28615 -44272 28935 -44210
rect 28615 -44508 28657 -44272
rect 28893 -44508 28935 -44272
rect 28615 -44592 28935 -44508
rect 28615 -44828 28657 -44592
rect 28893 -44828 28935 -44592
rect 28615 -44890 28935 -44828
rect 29615 -44272 29935 -44210
rect 29615 -44508 29657 -44272
rect 29893 -44508 29935 -44272
rect 29615 -44592 29935 -44508
rect 29615 -44828 29657 -44592
rect 29893 -44828 29935 -44592
rect 29615 -44890 29935 -44828
rect 30615 -44272 30935 -44210
rect 30615 -44508 30657 -44272
rect 30893 -44508 30935 -44272
rect 30615 -44592 30935 -44508
rect 30615 -44828 30657 -44592
rect 30893 -44828 30935 -44592
rect 30615 -44890 30935 -44828
rect 31615 -44272 31935 -44210
rect 31615 -44508 31657 -44272
rect 31893 -44508 31935 -44272
rect 31615 -44592 31935 -44508
rect 31615 -44828 31657 -44592
rect 31893 -44828 31935 -44592
rect 31615 -44890 31935 -44828
rect 32615 -44272 32935 -44210
rect 32615 -44508 32657 -44272
rect 32893 -44508 32935 -44272
rect 32615 -44592 32935 -44508
rect 32615 -44828 32657 -44592
rect 32893 -44828 32935 -44592
rect 32615 -44890 32935 -44828
rect 33615 -44272 33935 -44210
rect 33615 -44508 33657 -44272
rect 33893 -44508 33935 -44272
rect 33615 -44592 33935 -44508
rect 33615 -44828 33657 -44592
rect 33893 -44828 33935 -44592
rect 33615 -44890 33935 -44828
rect -74825 -44932 -48825 -44890
rect -74825 -45168 -74783 -44932
rect -74547 -45168 -74443 -44932
rect -74207 -45168 -74103 -44932
rect -73867 -45168 -73783 -44932
rect -73547 -45168 -73443 -44932
rect -73207 -45168 -73103 -44932
rect -72867 -45168 -72783 -44932
rect -72547 -45168 -72443 -44932
rect -72207 -45168 -72103 -44932
rect -71867 -45168 -71783 -44932
rect -71547 -45168 -71443 -44932
rect -71207 -45168 -71103 -44932
rect -70867 -45168 -70783 -44932
rect -70547 -45168 -70443 -44932
rect -70207 -45168 -70103 -44932
rect -69867 -45168 -69783 -44932
rect -69547 -45168 -69443 -44932
rect -69207 -45168 -69103 -44932
rect -68867 -45168 -68783 -44932
rect -68547 -45168 -68443 -44932
rect -68207 -45168 -68103 -44932
rect -67867 -45168 -67783 -44932
rect -67547 -45168 -67443 -44932
rect -67207 -45168 -67103 -44932
rect -66867 -45168 -66783 -44932
rect -66547 -45168 -66443 -44932
rect -66207 -45168 -66103 -44932
rect -65867 -45168 -65783 -44932
rect -65547 -45168 -65443 -44932
rect -65207 -45168 -65103 -44932
rect -64867 -45168 -64783 -44932
rect -64547 -45168 -64443 -44932
rect -64207 -45168 -64103 -44932
rect -63867 -45168 -63783 -44932
rect -63547 -45168 -63443 -44932
rect -63207 -45168 -63103 -44932
rect -62867 -45168 -62783 -44932
rect -62547 -45168 -62443 -44932
rect -62207 -45168 -62103 -44932
rect -61867 -45168 -61783 -44932
rect -61547 -45168 -61443 -44932
rect -61207 -45168 -61103 -44932
rect -60867 -45168 -60783 -44932
rect -60547 -45168 -60443 -44932
rect -60207 -45168 -60103 -44932
rect -59867 -45168 -59783 -44932
rect -59547 -45168 -59443 -44932
rect -59207 -45168 -59103 -44932
rect -58867 -45168 -58783 -44932
rect -58547 -45168 -58443 -44932
rect -58207 -45168 -58103 -44932
rect -57867 -45168 -57783 -44932
rect -57547 -45168 -57443 -44932
rect -57207 -45168 -57103 -44932
rect -56867 -45168 -56783 -44932
rect -56547 -45168 -56443 -44932
rect -56207 -45168 -56103 -44932
rect -55867 -45168 -55783 -44932
rect -55547 -45168 -55443 -44932
rect -55207 -45168 -55103 -44932
rect -54867 -45168 -54783 -44932
rect -54547 -45168 -54443 -44932
rect -54207 -45168 -54103 -44932
rect -53867 -45168 -53783 -44932
rect -53547 -45168 -53443 -44932
rect -53207 -45168 -53103 -44932
rect -52867 -45168 -52783 -44932
rect -52547 -45168 -52443 -44932
rect -52207 -45168 -52103 -44932
rect -51867 -45168 -51783 -44932
rect -51547 -45168 -51443 -44932
rect -51207 -45168 -51103 -44932
rect -50867 -45168 -50783 -44932
rect -50547 -45168 -50443 -44932
rect -50207 -45168 -50103 -44932
rect -49867 -45168 -49783 -44932
rect -49547 -45168 -49443 -44932
rect -49207 -45168 -49103 -44932
rect -48867 -45168 -48825 -44932
rect -74825 -45210 -48825 -45168
rect 8275 -44932 34275 -44890
rect 8275 -45168 8317 -44932
rect 8553 -45168 8657 -44932
rect 8893 -45168 8997 -44932
rect 9233 -45168 9317 -44932
rect 9553 -45168 9657 -44932
rect 9893 -45168 9997 -44932
rect 10233 -45168 10317 -44932
rect 10553 -45168 10657 -44932
rect 10893 -45168 10997 -44932
rect 11233 -45168 11317 -44932
rect 11553 -45168 11657 -44932
rect 11893 -45168 11997 -44932
rect 12233 -45168 12317 -44932
rect 12553 -45168 12657 -44932
rect 12893 -45168 12997 -44932
rect 13233 -45168 13317 -44932
rect 13553 -45168 13657 -44932
rect 13893 -45168 13997 -44932
rect 14233 -45168 14317 -44932
rect 14553 -45168 14657 -44932
rect 14893 -45168 14997 -44932
rect 15233 -45168 15317 -44932
rect 15553 -45168 15657 -44932
rect 15893 -45168 15997 -44932
rect 16233 -45168 16317 -44932
rect 16553 -45168 16657 -44932
rect 16893 -45168 16997 -44932
rect 17233 -45168 17317 -44932
rect 17553 -45168 17657 -44932
rect 17893 -45168 17997 -44932
rect 18233 -45168 18317 -44932
rect 18553 -45168 18657 -44932
rect 18893 -45168 18997 -44932
rect 19233 -45168 19317 -44932
rect 19553 -45168 19657 -44932
rect 19893 -45168 19997 -44932
rect 20233 -45168 20317 -44932
rect 20553 -45168 20657 -44932
rect 20893 -45168 20997 -44932
rect 21233 -45168 21317 -44932
rect 21553 -45168 21657 -44932
rect 21893 -45168 21997 -44932
rect 22233 -45168 22317 -44932
rect 22553 -45168 22657 -44932
rect 22893 -45168 22997 -44932
rect 23233 -45168 23317 -44932
rect 23553 -45168 23657 -44932
rect 23893 -45168 23997 -44932
rect 24233 -45168 24317 -44932
rect 24553 -45168 24657 -44932
rect 24893 -45168 24997 -44932
rect 25233 -45168 25317 -44932
rect 25553 -45168 25657 -44932
rect 25893 -45168 25997 -44932
rect 26233 -45168 26317 -44932
rect 26553 -45168 26657 -44932
rect 26893 -45168 26997 -44932
rect 27233 -45168 27317 -44932
rect 27553 -45168 27657 -44932
rect 27893 -45168 27997 -44932
rect 28233 -45168 28317 -44932
rect 28553 -45168 28657 -44932
rect 28893 -45168 28997 -44932
rect 29233 -45168 29317 -44932
rect 29553 -45168 29657 -44932
rect 29893 -45168 29997 -44932
rect 30233 -45168 30317 -44932
rect 30553 -45168 30657 -44932
rect 30893 -45168 30997 -44932
rect 31233 -45168 31317 -44932
rect 31553 -45168 31657 -44932
rect 31893 -45168 31997 -44932
rect 32233 -45168 32317 -44932
rect 32553 -45168 32657 -44932
rect 32893 -45168 32997 -44932
rect 33233 -45168 33317 -44932
rect 33553 -45168 33657 -44932
rect 33893 -45168 33997 -44932
rect 34233 -45168 34275 -44932
rect 8275 -45210 34275 -45168
rect -74485 -45272 -74165 -45210
rect -74485 -45508 -74443 -45272
rect -74207 -45508 -74165 -45272
rect -74485 -45592 -74165 -45508
rect -74485 -45828 -74443 -45592
rect -74207 -45828 -74165 -45592
rect -74485 -45890 -74165 -45828
rect -73485 -45272 -73165 -45210
rect -73485 -45508 -73443 -45272
rect -73207 -45508 -73165 -45272
rect -73485 -45592 -73165 -45508
rect -73485 -45828 -73443 -45592
rect -73207 -45828 -73165 -45592
rect -73485 -45890 -73165 -45828
rect -72485 -45272 -72165 -45210
rect -72485 -45508 -72443 -45272
rect -72207 -45508 -72165 -45272
rect -72485 -45592 -72165 -45508
rect -72485 -45828 -72443 -45592
rect -72207 -45828 -72165 -45592
rect -72485 -45890 -72165 -45828
rect -71485 -45272 -71165 -45210
rect -71485 -45508 -71443 -45272
rect -71207 -45508 -71165 -45272
rect -71485 -45592 -71165 -45508
rect -71485 -45828 -71443 -45592
rect -71207 -45828 -71165 -45592
rect -71485 -45890 -71165 -45828
rect -70485 -45272 -70165 -45210
rect -70485 -45508 -70443 -45272
rect -70207 -45508 -70165 -45272
rect -70485 -45592 -70165 -45508
rect -70485 -45828 -70443 -45592
rect -70207 -45828 -70165 -45592
rect -70485 -45890 -70165 -45828
rect -69485 -45272 -69165 -45210
rect -69485 -45508 -69443 -45272
rect -69207 -45508 -69165 -45272
rect -69485 -45592 -69165 -45508
rect -69485 -45828 -69443 -45592
rect -69207 -45828 -69165 -45592
rect -69485 -45890 -69165 -45828
rect -68485 -45272 -68165 -45210
rect -68485 -45508 -68443 -45272
rect -68207 -45508 -68165 -45272
rect -68485 -45592 -68165 -45508
rect -68485 -45828 -68443 -45592
rect -68207 -45828 -68165 -45592
rect -68485 -45890 -68165 -45828
rect -67485 -45272 -67165 -45210
rect -67485 -45508 -67443 -45272
rect -67207 -45508 -67165 -45272
rect -67485 -45592 -67165 -45508
rect -67485 -45828 -67443 -45592
rect -67207 -45828 -67165 -45592
rect -67485 -45890 -67165 -45828
rect -66485 -45272 -66165 -45210
rect -66485 -45508 -66443 -45272
rect -66207 -45508 -66165 -45272
rect -66485 -45592 -66165 -45508
rect -66485 -45828 -66443 -45592
rect -66207 -45828 -66165 -45592
rect -66485 -45890 -66165 -45828
rect -65485 -45272 -65165 -45210
rect -65485 -45508 -65443 -45272
rect -65207 -45508 -65165 -45272
rect -65485 -45592 -65165 -45508
rect -65485 -45828 -65443 -45592
rect -65207 -45828 -65165 -45592
rect -65485 -45890 -65165 -45828
rect -64485 -45272 -64165 -45210
rect -64485 -45508 -64443 -45272
rect -64207 -45508 -64165 -45272
rect -64485 -45592 -64165 -45508
rect -64485 -45828 -64443 -45592
rect -64207 -45828 -64165 -45592
rect -64485 -45890 -64165 -45828
rect -63485 -45272 -63165 -45210
rect -63485 -45508 -63443 -45272
rect -63207 -45508 -63165 -45272
rect -63485 -45592 -63165 -45508
rect -63485 -45828 -63443 -45592
rect -63207 -45828 -63165 -45592
rect -63485 -45890 -63165 -45828
rect -62485 -45272 -62165 -45210
rect -62485 -45508 -62443 -45272
rect -62207 -45508 -62165 -45272
rect -62485 -45592 -62165 -45508
rect -62485 -45828 -62443 -45592
rect -62207 -45828 -62165 -45592
rect -62485 -45890 -62165 -45828
rect -61485 -45272 -61165 -45210
rect -61485 -45508 -61443 -45272
rect -61207 -45508 -61165 -45272
rect -61485 -45592 -61165 -45508
rect -61485 -45828 -61443 -45592
rect -61207 -45828 -61165 -45592
rect -61485 -45890 -61165 -45828
rect -60485 -45272 -60165 -45210
rect -60485 -45508 -60443 -45272
rect -60207 -45508 -60165 -45272
rect -60485 -45592 -60165 -45508
rect -60485 -45828 -60443 -45592
rect -60207 -45828 -60165 -45592
rect -60485 -45890 -60165 -45828
rect -59485 -45272 -59165 -45210
rect -59485 -45508 -59443 -45272
rect -59207 -45508 -59165 -45272
rect -59485 -45592 -59165 -45508
rect -59485 -45828 -59443 -45592
rect -59207 -45828 -59165 -45592
rect -59485 -45890 -59165 -45828
rect -58485 -45272 -58165 -45210
rect -58485 -45508 -58443 -45272
rect -58207 -45508 -58165 -45272
rect -58485 -45592 -58165 -45508
rect -58485 -45828 -58443 -45592
rect -58207 -45828 -58165 -45592
rect -58485 -45890 -58165 -45828
rect -57485 -45272 -57165 -45210
rect -57485 -45508 -57443 -45272
rect -57207 -45508 -57165 -45272
rect -57485 -45592 -57165 -45508
rect -57485 -45828 -57443 -45592
rect -57207 -45828 -57165 -45592
rect -57485 -45890 -57165 -45828
rect -56485 -45272 -56165 -45210
rect -56485 -45508 -56443 -45272
rect -56207 -45508 -56165 -45272
rect -56485 -45592 -56165 -45508
rect -56485 -45828 -56443 -45592
rect -56207 -45828 -56165 -45592
rect -56485 -45890 -56165 -45828
rect -55485 -45272 -55165 -45210
rect -55485 -45508 -55443 -45272
rect -55207 -45508 -55165 -45272
rect -55485 -45592 -55165 -45508
rect -55485 -45828 -55443 -45592
rect -55207 -45828 -55165 -45592
rect -55485 -45890 -55165 -45828
rect -54485 -45272 -54165 -45210
rect -54485 -45508 -54443 -45272
rect -54207 -45508 -54165 -45272
rect -54485 -45592 -54165 -45508
rect -54485 -45828 -54443 -45592
rect -54207 -45828 -54165 -45592
rect -54485 -45890 -54165 -45828
rect -53485 -45272 -53165 -45210
rect -53485 -45508 -53443 -45272
rect -53207 -45508 -53165 -45272
rect -53485 -45592 -53165 -45508
rect -53485 -45828 -53443 -45592
rect -53207 -45828 -53165 -45592
rect -53485 -45890 -53165 -45828
rect -52485 -45272 -52165 -45210
rect -52485 -45508 -52443 -45272
rect -52207 -45508 -52165 -45272
rect -52485 -45592 -52165 -45508
rect -52485 -45828 -52443 -45592
rect -52207 -45828 -52165 -45592
rect -52485 -45890 -52165 -45828
rect -51485 -45272 -51165 -45210
rect -51485 -45508 -51443 -45272
rect -51207 -45508 -51165 -45272
rect -51485 -45592 -51165 -45508
rect -51485 -45828 -51443 -45592
rect -51207 -45828 -51165 -45592
rect -51485 -45890 -51165 -45828
rect -50485 -45272 -50165 -45210
rect -50485 -45508 -50443 -45272
rect -50207 -45508 -50165 -45272
rect -50485 -45592 -50165 -45508
rect -50485 -45828 -50443 -45592
rect -50207 -45828 -50165 -45592
rect -50485 -45890 -50165 -45828
rect -49485 -45272 -49165 -45210
rect -49485 -45508 -49443 -45272
rect -49207 -45508 -49165 -45272
rect -49485 -45592 -49165 -45508
rect -49485 -45828 -49443 -45592
rect -49207 -45828 -49165 -45592
rect -49485 -45890 -49165 -45828
rect 8615 -45272 8935 -45210
rect 8615 -45508 8657 -45272
rect 8893 -45508 8935 -45272
rect 8615 -45592 8935 -45508
rect 8615 -45828 8657 -45592
rect 8893 -45828 8935 -45592
rect 8615 -45890 8935 -45828
rect 9615 -45272 9935 -45210
rect 9615 -45508 9657 -45272
rect 9893 -45508 9935 -45272
rect 9615 -45592 9935 -45508
rect 9615 -45828 9657 -45592
rect 9893 -45828 9935 -45592
rect 9615 -45890 9935 -45828
rect 10615 -45272 10935 -45210
rect 10615 -45508 10657 -45272
rect 10893 -45508 10935 -45272
rect 10615 -45592 10935 -45508
rect 10615 -45828 10657 -45592
rect 10893 -45828 10935 -45592
rect 10615 -45890 10935 -45828
rect 11615 -45272 11935 -45210
rect 11615 -45508 11657 -45272
rect 11893 -45508 11935 -45272
rect 11615 -45592 11935 -45508
rect 11615 -45828 11657 -45592
rect 11893 -45828 11935 -45592
rect 11615 -45890 11935 -45828
rect 12615 -45272 12935 -45210
rect 12615 -45508 12657 -45272
rect 12893 -45508 12935 -45272
rect 12615 -45592 12935 -45508
rect 12615 -45828 12657 -45592
rect 12893 -45828 12935 -45592
rect 12615 -45890 12935 -45828
rect 13615 -45272 13935 -45210
rect 13615 -45508 13657 -45272
rect 13893 -45508 13935 -45272
rect 13615 -45592 13935 -45508
rect 13615 -45828 13657 -45592
rect 13893 -45828 13935 -45592
rect 13615 -45890 13935 -45828
rect 14615 -45272 14935 -45210
rect 14615 -45508 14657 -45272
rect 14893 -45508 14935 -45272
rect 14615 -45592 14935 -45508
rect 14615 -45828 14657 -45592
rect 14893 -45828 14935 -45592
rect 14615 -45890 14935 -45828
rect 15615 -45272 15935 -45210
rect 15615 -45508 15657 -45272
rect 15893 -45508 15935 -45272
rect 15615 -45592 15935 -45508
rect 15615 -45828 15657 -45592
rect 15893 -45828 15935 -45592
rect 15615 -45890 15935 -45828
rect 16615 -45272 16935 -45210
rect 16615 -45508 16657 -45272
rect 16893 -45508 16935 -45272
rect 16615 -45592 16935 -45508
rect 16615 -45828 16657 -45592
rect 16893 -45828 16935 -45592
rect 16615 -45890 16935 -45828
rect 17615 -45272 17935 -45210
rect 17615 -45508 17657 -45272
rect 17893 -45508 17935 -45272
rect 17615 -45592 17935 -45508
rect 17615 -45828 17657 -45592
rect 17893 -45828 17935 -45592
rect 17615 -45890 17935 -45828
rect 18615 -45272 18935 -45210
rect 18615 -45508 18657 -45272
rect 18893 -45508 18935 -45272
rect 18615 -45592 18935 -45508
rect 18615 -45828 18657 -45592
rect 18893 -45828 18935 -45592
rect 18615 -45890 18935 -45828
rect 19615 -45272 19935 -45210
rect 19615 -45508 19657 -45272
rect 19893 -45508 19935 -45272
rect 19615 -45592 19935 -45508
rect 19615 -45828 19657 -45592
rect 19893 -45828 19935 -45592
rect 19615 -45890 19935 -45828
rect 20615 -45272 20935 -45210
rect 20615 -45508 20657 -45272
rect 20893 -45508 20935 -45272
rect 20615 -45592 20935 -45508
rect 20615 -45828 20657 -45592
rect 20893 -45828 20935 -45592
rect 20615 -45890 20935 -45828
rect 21615 -45272 21935 -45210
rect 21615 -45508 21657 -45272
rect 21893 -45508 21935 -45272
rect 21615 -45592 21935 -45508
rect 21615 -45828 21657 -45592
rect 21893 -45828 21935 -45592
rect 21615 -45890 21935 -45828
rect 22615 -45272 22935 -45210
rect 22615 -45508 22657 -45272
rect 22893 -45508 22935 -45272
rect 22615 -45592 22935 -45508
rect 22615 -45828 22657 -45592
rect 22893 -45828 22935 -45592
rect 22615 -45890 22935 -45828
rect 23615 -45272 23935 -45210
rect 23615 -45508 23657 -45272
rect 23893 -45508 23935 -45272
rect 23615 -45592 23935 -45508
rect 23615 -45828 23657 -45592
rect 23893 -45828 23935 -45592
rect 23615 -45890 23935 -45828
rect 24615 -45272 24935 -45210
rect 24615 -45508 24657 -45272
rect 24893 -45508 24935 -45272
rect 24615 -45592 24935 -45508
rect 24615 -45828 24657 -45592
rect 24893 -45828 24935 -45592
rect 24615 -45890 24935 -45828
rect 25615 -45272 25935 -45210
rect 25615 -45508 25657 -45272
rect 25893 -45508 25935 -45272
rect 25615 -45592 25935 -45508
rect 25615 -45828 25657 -45592
rect 25893 -45828 25935 -45592
rect 25615 -45890 25935 -45828
rect 26615 -45272 26935 -45210
rect 26615 -45508 26657 -45272
rect 26893 -45508 26935 -45272
rect 26615 -45592 26935 -45508
rect 26615 -45828 26657 -45592
rect 26893 -45828 26935 -45592
rect 26615 -45890 26935 -45828
rect 27615 -45272 27935 -45210
rect 27615 -45508 27657 -45272
rect 27893 -45508 27935 -45272
rect 27615 -45592 27935 -45508
rect 27615 -45828 27657 -45592
rect 27893 -45828 27935 -45592
rect 27615 -45890 27935 -45828
rect 28615 -45272 28935 -45210
rect 28615 -45508 28657 -45272
rect 28893 -45508 28935 -45272
rect 28615 -45592 28935 -45508
rect 28615 -45828 28657 -45592
rect 28893 -45828 28935 -45592
rect 28615 -45890 28935 -45828
rect 29615 -45272 29935 -45210
rect 29615 -45508 29657 -45272
rect 29893 -45508 29935 -45272
rect 29615 -45592 29935 -45508
rect 29615 -45828 29657 -45592
rect 29893 -45828 29935 -45592
rect 29615 -45890 29935 -45828
rect 30615 -45272 30935 -45210
rect 30615 -45508 30657 -45272
rect 30893 -45508 30935 -45272
rect 30615 -45592 30935 -45508
rect 30615 -45828 30657 -45592
rect 30893 -45828 30935 -45592
rect 30615 -45890 30935 -45828
rect 31615 -45272 31935 -45210
rect 31615 -45508 31657 -45272
rect 31893 -45508 31935 -45272
rect 31615 -45592 31935 -45508
rect 31615 -45828 31657 -45592
rect 31893 -45828 31935 -45592
rect 31615 -45890 31935 -45828
rect 32615 -45272 32935 -45210
rect 32615 -45508 32657 -45272
rect 32893 -45508 32935 -45272
rect 32615 -45592 32935 -45508
rect 32615 -45828 32657 -45592
rect 32893 -45828 32935 -45592
rect 32615 -45890 32935 -45828
rect 33615 -45272 33935 -45210
rect 33615 -45508 33657 -45272
rect 33893 -45508 33935 -45272
rect 33615 -45592 33935 -45508
rect 33615 -45828 33657 -45592
rect 33893 -45828 33935 -45592
rect 33615 -45890 33935 -45828
rect -74825 -45932 -48825 -45890
rect -74825 -46168 -74783 -45932
rect -74547 -46168 -74443 -45932
rect -74207 -46168 -74103 -45932
rect -73867 -46168 -73783 -45932
rect -73547 -46168 -73443 -45932
rect -73207 -46168 -73103 -45932
rect -72867 -46168 -72783 -45932
rect -72547 -46168 -72443 -45932
rect -72207 -46168 -72103 -45932
rect -71867 -46168 -71783 -45932
rect -71547 -46168 -71443 -45932
rect -71207 -46168 -71103 -45932
rect -70867 -46168 -70783 -45932
rect -70547 -46168 -70443 -45932
rect -70207 -46168 -70103 -45932
rect -69867 -46168 -69783 -45932
rect -69547 -46168 -69443 -45932
rect -69207 -46168 -69103 -45932
rect -68867 -46168 -68783 -45932
rect -68547 -46168 -68443 -45932
rect -68207 -46168 -68103 -45932
rect -67867 -46168 -67783 -45932
rect -67547 -46168 -67443 -45932
rect -67207 -46168 -67103 -45932
rect -66867 -46168 -66783 -45932
rect -66547 -46168 -66443 -45932
rect -66207 -46168 -66103 -45932
rect -65867 -46168 -65783 -45932
rect -65547 -46168 -65443 -45932
rect -65207 -46168 -65103 -45932
rect -64867 -46168 -64783 -45932
rect -64547 -46168 -64443 -45932
rect -64207 -46168 -64103 -45932
rect -63867 -46168 -63783 -45932
rect -63547 -46168 -63443 -45932
rect -63207 -46168 -63103 -45932
rect -62867 -46168 -62783 -45932
rect -62547 -46168 -62443 -45932
rect -62207 -46168 -62103 -45932
rect -61867 -46168 -61783 -45932
rect -61547 -46168 -61443 -45932
rect -61207 -46168 -61103 -45932
rect -60867 -46168 -60783 -45932
rect -60547 -46168 -60443 -45932
rect -60207 -46168 -60103 -45932
rect -59867 -46168 -59783 -45932
rect -59547 -46168 -59443 -45932
rect -59207 -46168 -59103 -45932
rect -58867 -46168 -58783 -45932
rect -58547 -46168 -58443 -45932
rect -58207 -46168 -58103 -45932
rect -57867 -46168 -57783 -45932
rect -57547 -46168 -57443 -45932
rect -57207 -46168 -57103 -45932
rect -56867 -46168 -56783 -45932
rect -56547 -46168 -56443 -45932
rect -56207 -46168 -56103 -45932
rect -55867 -46168 -55783 -45932
rect -55547 -46168 -55443 -45932
rect -55207 -46168 -55103 -45932
rect -54867 -46168 -54783 -45932
rect -54547 -46168 -54443 -45932
rect -54207 -46168 -54103 -45932
rect -53867 -46168 -53783 -45932
rect -53547 -46168 -53443 -45932
rect -53207 -46168 -53103 -45932
rect -52867 -46168 -52783 -45932
rect -52547 -46168 -52443 -45932
rect -52207 -46168 -52103 -45932
rect -51867 -46168 -51783 -45932
rect -51547 -46168 -51443 -45932
rect -51207 -46168 -51103 -45932
rect -50867 -46168 -50783 -45932
rect -50547 -46168 -50443 -45932
rect -50207 -46168 -50103 -45932
rect -49867 -46168 -49783 -45932
rect -49547 -46168 -49443 -45932
rect -49207 -46168 -49103 -45932
rect -48867 -46168 -48825 -45932
rect -74825 -46210 -48825 -46168
rect 8275 -45932 34275 -45890
rect 8275 -46168 8317 -45932
rect 8553 -46168 8657 -45932
rect 8893 -46168 8997 -45932
rect 9233 -46168 9317 -45932
rect 9553 -46168 9657 -45932
rect 9893 -46168 9997 -45932
rect 10233 -46168 10317 -45932
rect 10553 -46168 10657 -45932
rect 10893 -46168 10997 -45932
rect 11233 -46168 11317 -45932
rect 11553 -46168 11657 -45932
rect 11893 -46168 11997 -45932
rect 12233 -46168 12317 -45932
rect 12553 -46168 12657 -45932
rect 12893 -46168 12997 -45932
rect 13233 -46168 13317 -45932
rect 13553 -46168 13657 -45932
rect 13893 -46168 13997 -45932
rect 14233 -46168 14317 -45932
rect 14553 -46168 14657 -45932
rect 14893 -46168 14997 -45932
rect 15233 -46168 15317 -45932
rect 15553 -46168 15657 -45932
rect 15893 -46168 15997 -45932
rect 16233 -46168 16317 -45932
rect 16553 -46168 16657 -45932
rect 16893 -46168 16997 -45932
rect 17233 -46168 17317 -45932
rect 17553 -46168 17657 -45932
rect 17893 -46168 17997 -45932
rect 18233 -46168 18317 -45932
rect 18553 -46168 18657 -45932
rect 18893 -46168 18997 -45932
rect 19233 -46168 19317 -45932
rect 19553 -46168 19657 -45932
rect 19893 -46168 19997 -45932
rect 20233 -46168 20317 -45932
rect 20553 -46168 20657 -45932
rect 20893 -46168 20997 -45932
rect 21233 -46168 21317 -45932
rect 21553 -46168 21657 -45932
rect 21893 -46168 21997 -45932
rect 22233 -46168 22317 -45932
rect 22553 -46168 22657 -45932
rect 22893 -46168 22997 -45932
rect 23233 -46168 23317 -45932
rect 23553 -46168 23657 -45932
rect 23893 -46168 23997 -45932
rect 24233 -46168 24317 -45932
rect 24553 -46168 24657 -45932
rect 24893 -46168 24997 -45932
rect 25233 -46168 25317 -45932
rect 25553 -46168 25657 -45932
rect 25893 -46168 25997 -45932
rect 26233 -46168 26317 -45932
rect 26553 -46168 26657 -45932
rect 26893 -46168 26997 -45932
rect 27233 -46168 27317 -45932
rect 27553 -46168 27657 -45932
rect 27893 -46168 27997 -45932
rect 28233 -46168 28317 -45932
rect 28553 -46168 28657 -45932
rect 28893 -46168 28997 -45932
rect 29233 -46168 29317 -45932
rect 29553 -46168 29657 -45932
rect 29893 -46168 29997 -45932
rect 30233 -46168 30317 -45932
rect 30553 -46168 30657 -45932
rect 30893 -46168 30997 -45932
rect 31233 -46168 31317 -45932
rect 31553 -46168 31657 -45932
rect 31893 -46168 31997 -45932
rect 32233 -46168 32317 -45932
rect 32553 -46168 32657 -45932
rect 32893 -46168 32997 -45932
rect 33233 -46168 33317 -45932
rect 33553 -46168 33657 -45932
rect 33893 -46168 33997 -45932
rect 34233 -46168 34275 -45932
rect 8275 -46210 34275 -46168
rect -74485 -46272 -74165 -46210
rect -74485 -46508 -74443 -46272
rect -74207 -46508 -74165 -46272
rect -74485 -46550 -74165 -46508
rect -73485 -46272 -73165 -46210
rect -73485 -46508 -73443 -46272
rect -73207 -46508 -73165 -46272
rect -73485 -46550 -73165 -46508
rect -72485 -46272 -72165 -46210
rect -72485 -46508 -72443 -46272
rect -72207 -46508 -72165 -46272
rect -72485 -46550 -72165 -46508
rect -71485 -46272 -71165 -46210
rect -71485 -46508 -71443 -46272
rect -71207 -46508 -71165 -46272
rect -71485 -46550 -71165 -46508
rect -70485 -46272 -70165 -46210
rect -70485 -46508 -70443 -46272
rect -70207 -46508 -70165 -46272
rect -70485 -46550 -70165 -46508
rect -69485 -46272 -69165 -46210
rect -69485 -46508 -69443 -46272
rect -69207 -46508 -69165 -46272
rect -69485 -46550 -69165 -46508
rect -68485 -46272 -68165 -46210
rect -68485 -46508 -68443 -46272
rect -68207 -46508 -68165 -46272
rect -68485 -46550 -68165 -46508
rect -67485 -46272 -67165 -46210
rect -67485 -46508 -67443 -46272
rect -67207 -46508 -67165 -46272
rect -67485 -46550 -67165 -46508
rect -66485 -46272 -66165 -46210
rect -66485 -46508 -66443 -46272
rect -66207 -46508 -66165 -46272
rect -66485 -46550 -66165 -46508
rect -65485 -46272 -65165 -46210
rect -65485 -46508 -65443 -46272
rect -65207 -46508 -65165 -46272
rect -65485 -46550 -65165 -46508
rect -64485 -46272 -64165 -46210
rect -64485 -46508 -64443 -46272
rect -64207 -46508 -64165 -46272
rect -64485 -46550 -64165 -46508
rect -63485 -46272 -63165 -46210
rect -63485 -46508 -63443 -46272
rect -63207 -46508 -63165 -46272
rect -63485 -46550 -63165 -46508
rect -62485 -46272 -62165 -46210
rect -62485 -46508 -62443 -46272
rect -62207 -46508 -62165 -46272
rect -62485 -46550 -62165 -46508
rect -61485 -46272 -61165 -46210
rect -61485 -46508 -61443 -46272
rect -61207 -46508 -61165 -46272
rect -61485 -46550 -61165 -46508
rect -60485 -46272 -60165 -46210
rect -60485 -46508 -60443 -46272
rect -60207 -46508 -60165 -46272
rect -60485 -46550 -60165 -46508
rect -59485 -46272 -59165 -46210
rect -59485 -46508 -59443 -46272
rect -59207 -46508 -59165 -46272
rect -59485 -46550 -59165 -46508
rect -58485 -46272 -58165 -46210
rect -58485 -46508 -58443 -46272
rect -58207 -46508 -58165 -46272
rect -58485 -46550 -58165 -46508
rect -57485 -46272 -57165 -46210
rect -57485 -46508 -57443 -46272
rect -57207 -46508 -57165 -46272
rect -57485 -46550 -57165 -46508
rect -56485 -46272 -56165 -46210
rect -56485 -46508 -56443 -46272
rect -56207 -46508 -56165 -46272
rect -56485 -46550 -56165 -46508
rect -55485 -46272 -55165 -46210
rect -55485 -46508 -55443 -46272
rect -55207 -46508 -55165 -46272
rect -55485 -46550 -55165 -46508
rect -54485 -46272 -54165 -46210
rect -54485 -46508 -54443 -46272
rect -54207 -46508 -54165 -46272
rect -54485 -46550 -54165 -46508
rect -53485 -46272 -53165 -46210
rect -53485 -46508 -53443 -46272
rect -53207 -46508 -53165 -46272
rect -53485 -46550 -53165 -46508
rect -52485 -46272 -52165 -46210
rect -52485 -46508 -52443 -46272
rect -52207 -46508 -52165 -46272
rect -52485 -46550 -52165 -46508
rect -51485 -46272 -51165 -46210
rect -51485 -46508 -51443 -46272
rect -51207 -46508 -51165 -46272
rect -51485 -46550 -51165 -46508
rect -50485 -46272 -50165 -46210
rect -50485 -46508 -50443 -46272
rect -50207 -46508 -50165 -46272
rect -50485 -46550 -50165 -46508
rect -49485 -46272 -49165 -46210
rect -49485 -46508 -49443 -46272
rect -49207 -46508 -49165 -46272
rect -49485 -46550 -49165 -46508
rect 8615 -46272 8935 -46210
rect 8615 -46508 8657 -46272
rect 8893 -46508 8935 -46272
rect 8615 -46550 8935 -46508
rect 9615 -46272 9935 -46210
rect 9615 -46508 9657 -46272
rect 9893 -46508 9935 -46272
rect 9615 -46550 9935 -46508
rect 10615 -46272 10935 -46210
rect 10615 -46508 10657 -46272
rect 10893 -46508 10935 -46272
rect 10615 -46550 10935 -46508
rect 11615 -46272 11935 -46210
rect 11615 -46508 11657 -46272
rect 11893 -46508 11935 -46272
rect 11615 -46550 11935 -46508
rect 12615 -46272 12935 -46210
rect 12615 -46508 12657 -46272
rect 12893 -46508 12935 -46272
rect 12615 -46550 12935 -46508
rect 13615 -46272 13935 -46210
rect 13615 -46508 13657 -46272
rect 13893 -46508 13935 -46272
rect 13615 -46550 13935 -46508
rect 14615 -46272 14935 -46210
rect 14615 -46508 14657 -46272
rect 14893 -46508 14935 -46272
rect 14615 -46550 14935 -46508
rect 15615 -46272 15935 -46210
rect 15615 -46508 15657 -46272
rect 15893 -46508 15935 -46272
rect 15615 -46550 15935 -46508
rect 16615 -46272 16935 -46210
rect 16615 -46508 16657 -46272
rect 16893 -46508 16935 -46272
rect 16615 -46550 16935 -46508
rect 17615 -46272 17935 -46210
rect 17615 -46508 17657 -46272
rect 17893 -46508 17935 -46272
rect 17615 -46550 17935 -46508
rect 18615 -46272 18935 -46210
rect 18615 -46508 18657 -46272
rect 18893 -46508 18935 -46272
rect 18615 -46550 18935 -46508
rect 19615 -46272 19935 -46210
rect 19615 -46508 19657 -46272
rect 19893 -46508 19935 -46272
rect 19615 -46550 19935 -46508
rect 20615 -46272 20935 -46210
rect 20615 -46508 20657 -46272
rect 20893 -46508 20935 -46272
rect 20615 -46550 20935 -46508
rect 21615 -46272 21935 -46210
rect 21615 -46508 21657 -46272
rect 21893 -46508 21935 -46272
rect 21615 -46550 21935 -46508
rect 22615 -46272 22935 -46210
rect 22615 -46508 22657 -46272
rect 22893 -46508 22935 -46272
rect 22615 -46550 22935 -46508
rect 23615 -46272 23935 -46210
rect 23615 -46508 23657 -46272
rect 23893 -46508 23935 -46272
rect 23615 -46550 23935 -46508
rect 24615 -46272 24935 -46210
rect 24615 -46508 24657 -46272
rect 24893 -46508 24935 -46272
rect 24615 -46550 24935 -46508
rect 25615 -46272 25935 -46210
rect 25615 -46508 25657 -46272
rect 25893 -46508 25935 -46272
rect 25615 -46550 25935 -46508
rect 26615 -46272 26935 -46210
rect 26615 -46508 26657 -46272
rect 26893 -46508 26935 -46272
rect 26615 -46550 26935 -46508
rect 27615 -46272 27935 -46210
rect 27615 -46508 27657 -46272
rect 27893 -46508 27935 -46272
rect 27615 -46550 27935 -46508
rect 28615 -46272 28935 -46210
rect 28615 -46508 28657 -46272
rect 28893 -46508 28935 -46272
rect 28615 -46550 28935 -46508
rect 29615 -46272 29935 -46210
rect 29615 -46508 29657 -46272
rect 29893 -46508 29935 -46272
rect 29615 -46550 29935 -46508
rect 30615 -46272 30935 -46210
rect 30615 -46508 30657 -46272
rect 30893 -46508 30935 -46272
rect 30615 -46550 30935 -46508
rect 31615 -46272 31935 -46210
rect 31615 -46508 31657 -46272
rect 31893 -46508 31935 -46272
rect 31615 -46550 31935 -46508
rect 32615 -46272 32935 -46210
rect 32615 -46508 32657 -46272
rect 32893 -46508 32935 -46272
rect 32615 -46550 32935 -46508
rect 33615 -46272 33935 -46210
rect 33615 -46508 33657 -46272
rect 33893 -46508 33935 -46272
rect 33615 -46550 33935 -46508
<< rm5 >>
rect -32665 7478 -30434 8172
rect -10115 7478 -7884 8172
<< fillblock >>
rect -74825 -28000 34654 28000
rect -48275 -46550 7725 -28000
<< labels >>
flabel metal3 s -57246 46206 -56845 46655 2 FreeSans 2000 0 0 0 Toggle
port 1 nsew
flabel metal3 s -21476 44243 -19660 46234 2 FreeSans 2000 0 0 0 Vdd
port 2 nsew
flabel metal3 s 22307 43278 25064 45617 2 FreeSans 2000 0 0 0 Gnd
port 3 nsew
flabel metal5 s -21182 -39506 -19396 -37434 2 FreeSans 2000 0 0 0 Port3
port 4 nsew
flabel metal5 s -68123 -893 -66309 806 2 FreeSans 2000 0 0 0 Port1
port 5 nsew
flabel metal5 s 25508 -735 27083 1120 2 FreeSans 2000 0 0 0 Port2
port 6 nsew
<< properties >>
string FIXED_BBOX -84822 -56100 44278 39000
string path -1426.300 1206.050 -1426.300 819.400 -1264.250 819.400 
<< end >>
